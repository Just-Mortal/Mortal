`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Dh8jYaDEjUNIISk6T5qegPKxinMKzapW2xSzbNSXvzIwV5MTAPgGIZ8+0S4bW/f
ZdkTEtfKwX0hMZLkHQYft4N4O5UOSk64VZxa2aG9taPgbXEJRopgOJ3zeeDx8Eaw
f5BWs8n7oWu5Jk8ldeMmiDV+8uXR5TYiphGxL+oQyXtbB5nS4myqxMif8CgODUyp
zWGAtU0rugunBPNUMCkWzgHCA8eHc29J4QfqZ+UZlZhTxCjGKp7tTsTtPS+E++6H
KAia9yRrRJvK9OSHhDKa4loAditmHYuoTqaYigEQkqcqUvDaNAntX3wilmpTZM/e
uyK3Wyus1OBa1ICdA1B1nlK1g2gDqVJUKYpk4zRu8MVoM/5lgrfmMea6vswV3fE1
12G6ay8ibKq27SetPgE0SuhDI7vminP2Tjr8lwP4Udd3zPyYdIR+GSv1ySTWlTEg
FzndGQ+G7yzG6remue9AhA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4ymXuwoYm2JmJlpCvrUsm1tn7DrV5iECy7L0hiS6yTKZVFHIBwJtKPRAWeLZ5e2
dS2sBBhpsOa0yBa+2RZvdexp0L8BBSeoFwNPSGi3TKFMR6nlB34KkKETw9UzEM91
k+OvywlTldur6UYSCNjgC0Npqjuec+kwpOWCp06JWJW7bAkOP2TqmXT3reEjBMPG
sbD71MY6zo3Vf2hZYTG6BmXZ8CIMg8ag8npfI6p6gMGr0OcPAnUDkKTuQ8lW/GEb
Lu2aaFF8lfXS4XkPKtTDliKI50yjhzgz6bLoTkaMkFS1vWrHvgbtk49/TDrmQhaZ
QGp78/O51mdHY5ZmVj+c6AMTnla8JcHL3/NNAcMA5v1twFDARxABrsrvjlso3z/o
p9gjqsS85iY/TPvy1uosfFW4OryE4AbnAgrkF96e7ke2XxunpIkEYZvfJCgOWsvE
U4G+NW+kyX0cpWJG4XlqRdoSX+qOrSzGboOrM0KuEjJ40s6lAY/p7v6uy9zZph1k
Db+RP7jlFeW7buEOwRkITdPJ9Z6FqCm0nbkZLUx3DmhJLhtrej0h0kVbHSI3+sQZ
sGkRvLZ+uUAqXGsitoMSKiO/6Hg1O4wAnaxFLNpEXH3iXfuiSkcqvLQGZMpd2dnG
bt8mRlkEgNjPYWWUoCxWrqOU7b/OoTSx09i3Gsfr64+j9t2ffDbtiSIV00HX0MaU
iHrXfWzqusQW9BunHwF5G1wOcCfXIOrVjtbCxC9t5i1dq/qTJxHxytdU636ZbpID
mGHbDs7KzmJRXlHIRG0bnGVvEeK2w2Xu6y33ft05vNeinaGUdc8UAOCS/0ywQlTt
ItCjbSi82fDHKpMZAnR+foni0zPnzVQ7B5QaLcUiU/pRgVm1PbXXjMBtDujTfAe+
q5JqNsfZQ8cGj3JA9vjuQbRpFyR3BjW1EbuKo6rUFyHKlXD26t8KewoRKareFsxh
rnFlHcOypHgoxjcQzD7bhYxp5c4cJJDN4mxTBEWDo/K1kFja9R6hGvWx+10V04D9
vM3fsydDxDrdDe0Uu5EJKJi13Tbp6GSaAxhs3Qtstj7WhI4b7prpiTkPpx8/FWeB
SDqCCBXpWWHoQLqv/B7QaezGyanu7FoEHilY1xSyojjm/2w0bI+pVXJf6LpwzkRv
U6JlmsI9Xv/hexeJCbD8VAWjQ8ehqKAxjUwZOIw0t+4IagKs7q/TvGW8kCxEowE6
hev1Kho1FaidXGZ6KLDuJy8TtyQsuDki+2jQkRJAYYH4CIFnOC733XF3cHP5qLin
TgPVOFZy1PmHXvjWxS423XuuFS7aLLnCLvvZneKOywVRW6byHJcCzsRUMilkVwqt
YyS4OI+eGmvu25+7XjbxkA3GGQxhpEcZgz3FUcRyIscEelkGQpN2VRIiZcGq85Fy
AY6m2wN3df94U9QWVpLPA1t1s1WWd6ANtfeKLjtPPnZ+RUU+N5zMxEe+cq8DRApk
yyQG9LEGb2EVaK2rt9eugFV9VEEmPxDxEgvFPk9/uvePcD3yvypCAmbOSCRHS3q/
joT0JTnREKmQpLfLh/28IQOy3LOxpBFPksfNjhdU9X/XJInfLzJIrGrPuZYi3EZd
AQr5W0g1BYiyjrvtSblH61D0tW+kCd2DXT6zgry9Q7UTObFOQf9RyECgDWKodqHo
f2qqUD6C8d8dJJooauZ081l9NvpcXbfRFb9dr3iZtsgrh2JJXQ28pDsMO1sCQrSv
yI74oIQvGxICjkZAtUIIpzI7EcTqHGD6YKxQAZJO70v9M2LnR2ocMLgYjFdrNlv4
iQKz05bf9tnjXV2l+UHNETcyFuuMVlydIvG4ZN7ZwQtHj6S+T0VIWPZlnFAGZcTl
TtKiaF9BPbBYy2Kg5nTu7c0GIkwt6LFCPKRj6CUJPTLlQwC67mF8Z1XYXooHTHVF
JUb5rfqJI4hW+jJMRbDAdDU6lWU7qnTCrQP4Ztq0I7/LqencUwC0ZLFY6cXiGZHB
rgVn/UzGS02QJ+3Y/QMeOTAyEAzb8jGAOBpcE7plSJ3tlv1s3wKkNfWuIHiv53qh
W9DB7w6SUabtHylPU64f9IKOhacknLzlOr50TJF7m722lCM58oyrByYSQsGgD38g
+YjLXl3JDcnWVkLgFAFsMTu1OhkVHy17fZ4cMLYMsKIy3Nrnx0GY4oF8Tnb8n2GN
Jcwl5glHaDXQVpIdru/SjO2W3HgwVnsCyehofl4oyv7+g30ayRRKLTzyQsplsXpm
OyltDvwBYNAJO7d60JBandnvaGOhmCmcD0DklcPGVaxqLG7squ5B98oB7TaQz+Ds
VYuPiFjcabpY+Wv5OpkwevdGFm94JWeapJCB/chQLiwRnntQFnjz78mU5Y9Z0DLT
hUjM11KuQVjpDO6Zepd6wH0RDgneMAE9AgaHsNrxnL4Xz1jCmWmPXcAl2dO9tuCW
z2NacehbaxDR9T9dAJmab0sfnh8PYwb+HbKVt7LEXKIdMfMuGrTp95gx8ZbO8QgU
PrIeY/Sr1LTiPljArHk+ERu64oSMuGuJkl6EFwdqziuMIkXnOZ+Njq6vhpfV9fkz
beDCKNYCyPVQ9tQyYyKmaMjCIuYb5vYjOle/htVXR7+sQNUqeAu8z4zMuGNrYCTD
G8594jbl7fQYS6gjWC2yMP1GeQi/HQc/1yXggB7pLYCywgEaWWvwmvnN3lLHmtLH
qhaYLyn5sPD0EfmU9NJSugKaA17qOW1/kXOEcZgAlEmvySgu897YqvpfDtuTBr7h
ceO6NJTuCpTJB+Wl0h/zVQLax6eCGUcNF6w9fAbzQ4HpmnQF6iNyaKOM2ciQySMf
MMzeK0d1/F8hIErpjJsqs0Zi4BDNZeJJw5wb8u7YLx8z6vRroXqs2kwAuUaKSsyl
RbvVURwJrSxouR4qQeX+sfphkeGpAcJXOqMPZcd1bsBv+K8A8kF2sY+NfonZgjG6
lqbDkC79hDK8CsBTW6EKbx8JNUVdu3MBg/xdyEn21BLraZkjHYrkXy35JxCxkQIO
xtDLb2TdsZ3Br0HpoGkvAlKmd+vFNZyRGG2R1Uy2HZ8Ssa4cgnor9lU1DX0TuZIb
SBr9+E4Yu3mM72APfs76dsJf3q581PG4sYlvfEeOwj0AdKNQYUZwnTybA5IULGyG
h3vhlwUjMgEjwrMgR+I9v5ST0v/OSZYB+Z++jrefVeqRSxQd57TqQiGLUWImfvGs
ncgdmM8Od8EnHZC32eMU+2vGj+eO7Y43GM1wHDTK30VrGKOeP6eyZjC+mPuH4G1/
Hs/sv85fqCxg2y28rrvoDXMqT6N6sbhCpBqiRaq37BiA28nL2+4+ZR1DbZovtGID
W96TIuV1PQp/SseWMZ0EWPVkaksG4j2XTt42QpZZ1C5zms88sK4O/H5QDYMOUssR
4ye3ZbmpTR0TnKUkAmTaQSzbrKni00vKjkzk+EsmIjPB1XUAiiQICs1eZvqZhUq0
n+10hGQcsmLtBP8Dt6TVNt63u8DWJCIqgUllN0W/yGU4RnPK5F7cXPGKI0gwdl3j
TCPLvOy3F1ktAHiGHaU7qYx6QOftSLSAHe5hIv5LGpkq9KKJu5gQug034jbWbTZF
Z2fRTMnl6G2j7hzCEy+Y5vL6SJifZXKQB5o58UTc+l6/znR11K56elw3HMRdnPg/
sgO+rKt4yABVva6Sj1VAWYXqiYbEXaEurXtTz+x/3VyvfdGhCOTgfbsK/Ojjp63B
uU3a/7+/aAzvh4E7lHw2VNrDogxw6v2geqjUQln6tgicClmtN1lLMzhvAj1UWWbw
Zv8WIb0kVujtDE4oxNmVMCxWuLAOKQAuLUBRxYz3/SLL0gN2MNmeNttkOIMHLuT2
QagA3yUH7rnWJJyZJLe0q+QwN+7irsrjBp9QHLAT5iWJdtktpaMkB8sjXIK55NOR
9O8+I6jymbkeFruo0zem8iG5cHSIT67M3v37js0iqq6l6FGgIbxVPFVOGPDzOJkF
z+6DQyt210Vj1dk7ebxgeqvrf5KcPVO/HrliqTLqjPes8MANUmnx57/oFSeA+34a
cm3U4H/H+hOIFQl5JxJOMXDktMalQx4EQvcEGKxDvr/FinM+BBcWrQkjqa+NKgE7
NS1zvRd+qo96yTt2v2M6XbLrz3mL2UIWXd0y+ohWON7ceN0qPBG9lqbLBTKnuOxY
KWtel/jYLjk0Hl1CdbOJhYGYGpJ4qj61BjG0UQxITfqAS3xQN769vj9dFeceiv0l
b9C043GapGDymjyz6pmetbUucaC8yulSxW0kPB9hZ5wT0wvvjxBtYnabUYIWSa7m
6F4CPM7JOpCeI/U5/5k1nqlDaQpVLUyHaggYxTf70gcXvXHYE3AUMfmIJh7qjl1Q
v0gU1fniAe6j5gxPKJFQcvTUwbPPWbqKJ1YqjUgVU+xirgRPHLW3xqqBcVNR3OoO
62Ysriv3UXifNWpB2XGwhntoa2jQ+FT+MhLDcj7l9Uk4hhrgiY4uZnEmu/oOaZEv
dHN5pK9n7a6rwFibVskZDMiE1VxZF05vyDdTTXV3O4aA2nFVek2DPxLkpYPRtjVv
55ZdJMt7dpqYujfZUgJb0nwvy5BHqWfiJ/2BtyViQHNr3CFqRxIJBse4/SNGAgH0
Ly0JE+3JQ1ADKn8QFYKTRJ6rBMBCH65h9voMmxZ6S2c0lDgYQWZp011Adb8Av/yS
Fe9mcYbusUUrbiLjQKTJRGlXjV9X4X7TP2i9ehRB+SzD4Pffe/wP5c7Bu4/Im3MV
BJzz2UfM3YY+yr/2+bjlZExgtxdLHIQXd3kNWs9Mk7BrJ5gzmGHxFcYi85yKCiXy
a00nZedlU1VbHPtZslLsxNJQ78iv1mYdE7dxagsU4tpvr6VWd8y7tGnayWfX4/+H
GyxmA9onXWWpNH1sD7gDsJi/DM75iPHj+boGVvSOa6at9hJS+q9L+6+lscLrpdcl
+CkQM+jS37W5YqN5euCCS+ztz2XZtblh+YVnr2TjxDAozLFtHHHs2le2BqSTu4Ia
QKw8zy8kLoUQ0gVc2ETg5B06UKGiS5jYa9whsZjEoOOS36f8rLq1yhxmvozT83Ec
O8f4C55/MCH/WmEWKRvrmWbMxvUIDejdoL08aUsknEdkz5MTlbiYSmJAoUWUkLRy
pTACD64AhbpV/TsHDESsUPBnLTUg5gyMTVOAMexbx/7eSJ8o75SzEuHZ0eiLyq04
OD9lKVOGR0F3eq9rvF7z8SJ3PsQYb37EmMbZVbWw5RRK4SNobHpBXHlXlwqoO5x2
JOvIZyeCnUpOjc/P3mV2IKyI7BUqDzE/i8Js1TASINYZIGSAT1KuN8WlB9DQuCRB
fiMBKSHUKkZQ5sInz4HCeKRYFcpu9ReW52VJoLVLtMULwdH1YvQ2BQqZ67pxbpO0
oIrvk8Oh+nc7f8I7nBtmXCczX+FBMYgN43R1HxjgSAucDvybiwGetRgn1J8wPwLq
OJ+lQs+ojANKASD0JeK0k2jlBSgLdOFnl1ptsW9DUc2TBbVK4RVGzakFHwgrFRSz
WD1QO7X3fx2hnchsAdXCnTgx7970XJrMAWBh4kmolKRLL4jGOy3qzSO/IjUwfDMA
4VyecYQ/n8l4wZ0/KPtbd6YDyXYG85LdL9Gto0DwBnv19Uo+3csVE6HJr4RZRfPM
LFslVQX86lSZstIgcRPypiVnTfJulev7wBDD//3nnXhzdIBEmXQ3/RLrUdarplVU
oJUashA8wS7NPhWH3vakxevqK8bUr7KbQ03pZ5phmBog70H2UIA6vTjwlV6xAzbk
I2ApFHg2bfpSCA3HtlVdgJ0khJGw8IzQdo9D/8aAgjT9qj4PVB+YXXg7XOR9hB8u
6hPEJ2SqL/K8NRgR60EP3176KXHdu1mnPgRV/pouTMmf3BPKDhGwjDnhO1z3FFGV
B7B26sL5flWwypFtL9MoLTR/HZUFcHJGlOXzNzFgl4fQ3UNEs/uBYVCFLqNQBBOK
xh+0YvRZiPcYiEHbILYTnVYFSIK7o+rX4uVgQ+laSIqLqJIR0bzcNJrbrsPSQmGH
i+7bWNf1u8Ghrdj7C1Sdvma7y5KDcl8sHPxF9YlkifQSCx/FJ+k/kq2P2GCx8lDs
y3aGiI7M4ipt7di8X8ilK//FB0Zg0WQuGh6ZrhXvpG4u9hOO4QODlb+JBWt7DJPu
7fEjJORCEWIFTnZ5SukRFnWsl5UuZT6kUp0BtbzrMpfBNtV8a4Kv4zeJEVHrBYy0
zmI7tpziXa1kK7+oa96lnqkVQg+n8zhgy7t+KIIDgEgAQcscE0qL7p63vXpCT7Ls
pn35Ly1C9aCnDF6Uo3g+N1Nemv7nyRYGwc2pDktoQMSrgqTI+Zx9uBYSpDXcZsXH
VW4GrPVUxneB4O0MUrQNiUfHrvemvqUswAQITm9Eezy6bIPQZ1+sMT4JYXwFkiW/
tXMIr/nJwMufT2U/g+no4SkZH9kYyCxMZMiXJTHgNtAxQ0STFS6vUYvT/Nq4NIVe
wnkx1LjX1t0EdaZtLhiAAU1/K9/dwr8zoFdiBVsshQqOWOEreNkFvHBaq9D7Trnf
KoV+MQheiDJsz45tlup3uwtM38ZFdI8Qd150ZC5oFVbwaVVepI8vWbs6LzbUNzMY
6892UVgEc30i9pSxsfqw2ufZkDRz3cfx3JrPSkfFWnbpReekn+3OJcb/SvuCEjAm
AA+ob2N5nQsPcDE5OpvrQdp+0mIdz4HGhdrEzGidkrx6xcxoB1k0iCmENIUmvCSD
R0p5qzbOOnOGFKdsl0D/B2f2AsRargexwhD7qhgBWjbKC1dCDgekJkvkIXGSoMcX
uhba+6As6yG3pwTSWK157BWvsv+156BixY/HZLaQdWSskQZkOuKgS/jgRuZA46x4
Pvkf0VUYr6ShG2JNBkczp874NmpnpstRStb7EMMFz3byM+kAdSj8UN0o65R+/7vp
ebtOjj2IfkoRCvxHssEHpCAydkrHLrIGjX1Z+5DkMEQ0rTt7cZql9dPFGWsZIZwF
tPnaYM27tCgUTr4EyHbvo5q0rpB7U4Om8NckD23WJK8Y/rWk3IwcI5OBbbj3sI5J
guXfQ+iqqR8yrn1o166phDbj+R5CMkYyDMgpNfn9Wh3U5jBXXqj0jP3Bt3xZIUtN
FtG4uoO6etnaMQvKhxdySGqKG+9fDy8Bd9SBxRRjKxCivfUXciKqWGUNybp+cjXs
GI5SRZ93sfAGNZMqXZSCdKdW9amgvd8+BHGDJm855+Ar8G4bA61H91F0UmsV60ev
Rds92/Af5Ipe5Kx7MdAHPy2lsbH4lm0YPeyRpxjv62NG1NITLTZ4qGlr5UwQJceK
4MpWr+XFyzAGSgGrinxycnbs3mf9Wh13zhADMyoYyy1vmrV9U5Xj4pOO9XCtZJkO
lycBNgGhvlKpI/XHhrfw8aoEIt1rujDbwCDAT8cDQcIXAGqhunNCvBn52IAeXExg
tKacIWFjWMwcZRliFsP8Zi5Anx2qwQSssBuzvvISBDf3KnXtW0zkWyF85oeIwzA0
owbV4/DAjEmjRDvvtLcLuczVsZeQNgYu9Rvy/xHNC/Q0thaOnr+t9GtW2saoyI1I
ZCSiNMORveH5d7SYFJD5hOgUHr5bZdQFaqTcOlaVJ7poVJ4lORrJ6l6tCycsd/Vu
2ulppwR4i+fI+kKKHiMOEOJW/xrZ9G93vOAaaV/qCC/Y1XmphhCD5/6PFDskuABo
89sknyV4oXl/I7hE/fOqBeMmqwN3YWFaOnGijc0XHS5399/XxEJQjr3ruqhZSiXy
8ojLtsiWICK4w266PK6UPB8odTRlLS1aDhxAc/rPenTYXdAMAWlr9rNcp9w5Ei2O
Wzqr0vhI4zXxJz+2C9B0A5/+vvpsxgmmZJ5SIF2X24aEuYerbdzsX227/9jfgy/M
QOpWcmnRGMMSVNwI0R7sl/Ie4nLMnBu5rd8pUAA5y9rtd3LqfRMQDDCPLh+IVnC0
T4iCeYzoxDgzYE262op2RV/JhLDjLkQohuVf9Ot8AIfkNcvJ7d5N/Tl1dnZ/Ee41
Nma+Uq9FhQnaCp7PFDSBixFxwSStMJerXN0GP1fWIY4Z4bIC82jV2sgZnjNkoVVx
guNJo306+f0/jYkZCWlAcpXaCL2yxBi85WTzeZZxgA6nAnR3JzQ5m7VKFLp/dLMM
khz0vnNRR1rP0s8S2dyOt1VAiaqXlUpvTYZukee5qZl2W85EGHMcPdc7xfQZx34b
2d+elE9cb3WgE20koJ2q2cNQih4mQ5Q+ZE7+yddHuTyBZosoc8CQ0hAmlVbk+1kZ
gzBmayhSzYUBwf62+cAsfmuzdMCDHCUGnuXsaziiUWHY+Ak1JmrF+aEFocl7qumL
WFBZKDteGccmyeSU0b7zi6FvHawlMdrmBcsMVL0bIcrjx+DJu8tJSjJ3AsMLCLEr
pYSGVH5YknyE9mlOaf0gCLhqzsHXOs9ceYbNJyay5XIKpXv+75ayUGkaurhMSLDm
tMnIFeoMzhFNV4YQOUnjX7cn4bXKchtM6ELwBBXmQk6eEoDj5l6RL/i50I5hfYKL
X0S+lwLhAaUKM85MvApVK3YTYfViIOoRSAi5n3rOk7FrOh+rLecCKH3ESaSmwY2N
1t7zhx2TzIGyF7zMJUttfx1OH5V4d5d7RlIq5QD6WzZtUX0u4VcAPNFCnpmFhTC5
hzxkkAshuWGeEuMjyec1QEyioNl4J93yYACZKvOPjTMQ9lHpERp9PoFDJH3TMNJZ
96cJhLeTvaiVDolJQLCHltlIOff6CGCMXi6zb4CI39xZJqi23ggqdlzZSg7db4+H
/F3zOJISyX2yWQUI+E9IQk3e+DT66P6KjmyWLdZuu+FxfCxW6fjOrb9HTxT6/3Jg
3wi5/G9FraT+DfuwNq9EbTqm2aumgIpoOGKtx5DscSHWr2H5boifxHm7J3Waoa08
5u0Nm2lxFNRXYB9b6EFPPs85KzKtvueVXSKGMECs9HzUqv5ckRl9asHeFbD/wePn
95fTb9nT7eWQxoxQpy80IzJ2ugP5yeIE2LdE99EdsRDa3Hff4D2vBfLH6/orJnza
c22WEP/3HictrPcVDwvbDJ0aJibi9GZwPRlmUqiGAnshDm1zeh1sRi59jJ9ZFiSW
oHIvtpxORFO3Ugsnhj7f6N0/3Cx5ZPSca8VE3LlzH1xIkSw1Ylo+B5ejil8/zFOt
LCs92Z6kBdsqywJu3D3UZwJcZHykOkNw1YsKF67F0V73K89MxQaDGxF6cP6nQ629
Ww252aGD9zhQtdr3vCmLguKnRKtIBE3+y3mILaW9PVOe7gSTH4ksrCc9UFtecO0L
X1tA0stqozm7R19DfyqbKOcZYYBtLzoks01sqnN3oDHdxORNvYmaxCDgCVUrBUu8
8nxOkJQQZuBonv6DmkQs8sagd/666J5IG9NeVpptCRWu4OxfTxy6EbaywpNLp5DO
TYYpsecbSkp9zZbjyXQ1rwhFLFNnkkPq9n6/VQjijzDtUjFhZBnG+6fFpASulDLT
D7wfeRQRBbfekNXU7FRid/vHkexTHSW+zg8t2AQtngrYMaA8fzJPWTURxJkmBVjs
Mdszm+2aNnu4eWhXsKzP8S0BPHzBsxDNrQYURHA6MxjvdpNznGPpIt8v6BaLnPbL
BS7e7IzTAlS9x2My0Pt5os7sGdJARD2GvhBWCeOaMAitl/d267byFJ73C/tYTnHD
LjIHKlJF/g3JZApuvp5qETeX3AX28icN8wkTtAmuR1cl3vPf0t2N8CwF8yOtMbo9
J3wvWhRJfHPoB1nXLabKlkIlidKueScUE+F2a0s7aZ0cwyumWWPJ+gYGcjyySyXk
uOQUMDSsQHdm2MMKfH2X+HWI60iSyBmqJdFweK4y81C7q3cuICWxajda79qK87i3
O1954kgp9ksDVdUfW8jlLdE8LjbXKXcp0Yd+XXsiy3H6zyiKzUiKDhDnHylKQx6p
sPS2X32c94No3xPC/AqLLB1ItmoAhsc2cqbX1tWYPYAETLSEKwKahMsZ+5Yva4IG
qO6PTHtIThKwloqjC3riUOglJNq+O71k9c2pl//mGC7janoH5AButxkUJyuvAWay
YhIW26oPtl24brwev/NSNcoanjVnn3iceFlezDdmEs6WUBJGnbGynHgvDQOUw0zA
0bT4xBjDJ582Cg0Gn04mNIomLLo9dScHxNJCUPEZgfEOMoGHIyyAW51iT1OaIw1Z
PenMvXle6CgiDcP+hhbAqzER+B7MtLr15ZsgparEuQ/Fm7XErkipDuwIa5+VCvuC
K7s2ZqOsyVCpJJpsZUC2XMTv0SpWRqDGzV1n91B4I8TQAwiRXxljJy4NjdvcIbCh
Ym96RwWQv+lyGRjBa/cU1J0EUX8rf92O98nV2UbZpQx0FbwWPSONyE3AW6BbR+lV
fdm50bvirvHgaJA49XC84S/ZmsdEptwoR9oZoup059FBmaQyN+4EOjTBy31MJfM1
2VWgVYSgZCvdt4Kf5Yy7dLoKepY26j3H8+mq2kTjlWli0dRWMhMQY1YCMSXau2Um
HNyLSuSXQcJHCYs0sfptKA==
`protect END_PROTECTED

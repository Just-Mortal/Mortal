`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yF1snTSuulS2m79VEE0k+RqMGQ1FgzrbBpkrt8gyfYaWvOGJIbrtvA5EDpGPuAuu
Frl4OyXSx3NDlVswF/NUjpDt7lOjadzsh4kifzgw99VXgJptzYyda9RG7vv+17Q6
4qxSRbMDBPntbQ8SU3hFh16BzkZ1ThjNIFiHJtvPsHrrDpdGwRcxMTOoP8sLLMr1
EoOxXVL5h/B+1rVmrHfXJJwq6GuJkALi4orSLuMsrsB0xbwpWVxJfUSUe+01vzet
amsuomsC7h1zUiNBSnYSnGyTboPb5VOHJekGJrqz5jmxs9tP9tRnRYy0pRZ4Ty34
BQY9tNN82LjdtwSduAreCmfikDzpcHwAPLkIJJZ1MvnQ94kyXcc8b7njW9hiJ1/6
gv703swmHdydirMzdV2CzOXOQgufOv3yLVjq1pEWyJoOTwgaAOyZCuVaarfi/OG3
9bLBODqC7ZIlXhPcc8vb6mXPYmN3m9RFUOS/4B7go7FTlUmcLXDqHDpyc+/u7Wos
DZz6xa/UVrluP9YVmLWCW02gXVfWeKCgwMgw4wlHvDpWTd5V/L0+cmEkMnuYQOxp
X98l5+pkTKNNOSOA5m5u4RYbb2dEdIdpCF6PDN7R1wjYMCtfWTq0sy4X6nATFPrg
fbJeH0PHhE7LksKWC0qb309cRczzjz0e3j3ifJQ1wl+l6I1rx/UU4rlfTCbDW6PC
/ivNGt4u/5GK3gHFfAKqQMKwcrZy6kJ5TCnwdiesjj5r2OWz5tnHpk4Micdz+7OQ
P3eqVQkVTPMBw6lfhgGW5EJf7WJ8wKyANOXP+wibcd/7nZ1IwIRuHX4XcR49qHnM
8KyliJZyh7gBZf2x9nyEaHPTYq2RxSLEqAwGslHkoJnlxlG8rrH2RD9nmDdRf+zv
Na5ch/E84hfemjFNV56PZcuQpDxn9s3IvXjNspEjgOOqlEfOwLDK/o1vDkO5bl0l
ccI2M5hkixT7SMnNVlrv+QTehxqEId9Ss3enlrHKDwHZX0JtCOxS+DAUJX8sFrDt
RCorWMcq248yRXomvg0kDP+UcQA87Y1FRGWb0iKl4QYcpJ/xtkkGS4UcoSDPLIOg
R7zP0u5/DvWBmpr46s0b3J1IIYdLXH1s8OwCdXzfHF4cz4qk2UEdXU0Tc/CPoAHs
0vDggPiOXNVSj5GTu8GcO+AjfS/CkQ3i+G5zrEOhVA8hIAjW+pLoV7uS+Ip+s2r5
rlAi3c4VLZasYmFokOi0dynr9w+d4Ugoy1NJ+fy8V0nWFnzpu49A+kuPzPRJ/Yl2
Y1Rny/m+sCirtGpo5TCJ/R1Mh/LOzbq/pwaIVteks/bIXHD86rdgKhoAmkfvG8UM
/w1FGl+qaULB4Z+/5FBFogxghaSShpLBtMXgG/1Dbvba+HCKqfD0QWkYJ9OCw6Qb
sQvBfyY+boDTgUu6UtUqHtbloKsT61WJ85HXtrJuKPGrvY9we3M7yaTYVIajltFD
mfO7Yvwd50h4NgkdP/rUj0tLXwVrMBmQSc8KEOSF99ibL4EdRBLjbAms2P6FdZhq
/Pj+oqKNGvvzkxOBQskug0bvoDR5LhX0pIeakGdrP4BBqebKlAjuAtMAXImapbbq
91Q32fxwJ3xd/q9YyDM1OtZzsMJOAG+92AGanGbYrkH90c31isv295JWB0L8eMQ9
vRcNDdtdBD9AEnJYgAKIfqWXYUqhqVmErp3145Sq730HAhFVo7zyPHUvAbtN5R7s
Rg3x5w5jesGh2DLoU5nRsnomWgiZSN22Tcy1Y608TSnwfNiSVBvVSZCwjtr1cqY6
0+kujdg7jPm5AWoYPuPsfa4bCQ2C51dT12NVJoGXGXNO1bi0KJB6xMFSMSmaJu1J
D1brWAnZBEuV1DIWi9KAvg3AlRUANr/Th/gKNCUuOuwHjb28YMSZ/bkObINV9JX7
1+wDsekfK/YrPkYAz39Z18z9fxSGMRYbP+KNEQpgAZ+/li3AoSQM/KDBdHpoaC+c
hxqJBf5ymc/at2uu456CbAZf8Fxem/ajXcLX5Hoz0u6JggBWA/C8iQzCXhur/cDX
8+PH9mwDiRoIuDuNPCWTCw+lRuR3loPBavU7PVaxl1z5uewa335KNk/vSq7rv2WB
pAfKF1V7ezajKb7QGPnOVVSj3/wKTCu3FnpEIlP84op8VTTN0skMBfXD6MuyTpBA
GzITC3Irh4gOpjlJRLnc1LeEZxtTXzsPQBUd5Ozz3s8SieSbYu0PHOF/4HOk4yOo
+AQK+cccME+N6fTrjCPFyx0CI9ISkqfc7qBDp3ohFP5dEfP0gHk9O047XKrnqUYG
IbAqVrsyecprvkNYyPC5OtTZxBXqxePZJ9N1d3QrXjKXl4+it4+G3U7bHzknjkLO
gz+SdKSpgfVhm0Ln8l3PeXHquv6M1nmMFLAIayoXuSn0QkmERX1QW7dJYpu7njni
qzLf8rqjux2a4kH3m8swOnC4gzLYe95CbZXQDgcKEtUYqyQK0x+/+inmsb6hWtVI
nHbAKMAHwLnJOSPysBP0hX/8DkteSrEdvJNtx4Kx5MkCCJOz6FhBymwYVLKl7JxH
borRRG0nRc2DuZLjjl+k997erWPMjeJub1h+vmxsyGk+mHmwNNMOg0WS7sX9vLZe
E4J/vRElWqLYe6AvhSiv8Fx+D039EGMkpMETRgE5tm0yVdvQ6VP1VUyNykz1FAMC
B5wvafYv2foiqxBxZgJZH8xS3bilwJ8oeDtKwBX3MZtjaJg/3OI4vOvRp1d5Grdt
J0PjdI+FPE/Vz3OIqNb3rs5i3cxyxBj7fGc8Ia8mNi8ctLbMUukW05lzEsEd8eQR
DTVLlPNGAhyll0euciSAn/8+khCnwDy8M78bLIMSFKmU7YqBXtN314ASUEFOEVW6
wpQzbFBbxLT8mc5bUw4CvXK+jO2wPjmxdAjsy1tZ/9Xs4xoT0Fgemq+5LiKGAw0m
UOUFhvbfzGWumArJyn8XdOrbc2JNcIc+aEE0wHSxi7NvZ97c8e8FbM1apbmyzxvZ
qkUSNvaeG+tHtMw8hgfPmKUem9etF0t/Ek4ix1MTK4azqqMiHvvrPYvenkGr7EqD
gS2CgQ/PlXqJkRQT/LYrwKJH2mA5KwVyKUKx/VOM4xWahqrsUBCoM24n31pWWo//
42giJEmQaec5evDQ1gCShhBT+2QWTPNYlAn8dghlkaoHIqVJsj7XHUiIhwWmSJnz
w2lUSxom66XLkim/G2DroY4gENQH/fiMVehhwFqChY6n7pdCUz4eXTcjJ2x5yTPu
WOVOusrqU95CEnffUt7TDL5y2y5mIt1ApBraTUdF+VVp3PoTH4bSMwXskwt4xTvR
EJ4io8ulnzk06EI7DS8n+3k3Omaj9NZ4NgWEEqJHo7aDCaxwHFQn125SzmJzxiyw
pENLspNsfNWVNbpcpDL2o8gr7mbsFRWRawbe7JpFa/DXSoNpF8oWmJQq7XiD9RhQ
tabm6tcibt7iaXw5iVVTCvHCeDKozxmhQBtWPNTH9c/KPq7mLeTDcVZRhDdxRVdi
wRHaa2vpVssZ8E7f0IYZDSmquOAQBOMAUFu6t8miNAT8jD++BXg0yLjrrgVw0zg7
nNNfHfoDRdwUPtp7MtxImHsIq5IzOOYl2zr9YaychUkf3uFr9bF+OEj/JzK4pTLz
PrS+/qe/X0YGGrknanreNZeaC9JHYgpWrwb1uttewJwhpsovx3AlfTHup+NhkPLI
l5OJb5tJgCqDxsDt5W6G+UiQy4wAi2mPQNbBOVuIkxwc/vXuIaITL5hA8Bdjx8bm
SnXmRrqU8Zc8eN1DAiaJOA==
`protect END_PROTECTED

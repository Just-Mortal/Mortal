`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjXmllRSN8jROfkeSs+QrywOGBNNTA+3jXYAL2R+WsrY+BVXBYKC09GVJyfcbfUr
FG3SMtA8PfEXOELct+64KTIvF9rbrV9IYVgu1Uwvx2xGLSjG5DvAOH4uJPXoXR23
r28OSiPtS2tj63aXVs9STlJxBhvjmXqzWCjD2MjeeWdfVujRA853hhwbUS7FlfX8
VLsxTx3l657HCzsf845rnrYE7z3RFyQhWcPTJU+OfIfn3JFpzvnHFvWn8v1WXLo+
yyLvwrYzw4hDiVU7OBgZe+gG7oJX8gUxuLQsycabY5sbZw9KlUuwyeaNszufH7N0
VbiQfG34cqzHCROXAf+4LJ2RfJfvM8EFaUQmA7FsKQ2YxfBmqvd750S49nk2jG0k
L2Im8MY9tt45YQtInfatUxAn6qNtsaYtpVh690jmtG4rytX68D5mG/M5ZNi1hPwZ
nd3YC0sKRy4vv2dNhpE/NB0ek5yd88EzuzC4MrhSBvGMrdOZgkZn2D4qeuGCys+H
9WvJPjTDGm3+LQQmVaMc3y1s9wPVfSvHpxeS7vRmYSgWWWXMMY5V+X/jkDilynKh
PUnLG0eJvPkIrvWjBeSghNT1imJSyx6cGiO+1T02LDPph0LMdhmSw0sOW3pN4Bdj
667YnxdQz6DrwQKC40xIPnjX9VoJV8kMsaIJCpYqvvcXzyPpyiKCBtDuJm+/U+UN
sPt6A3RGzuJjyy+46BNUtTJZGSXuR5UxNjrPG/UindXV2JXtHrmkkESIJxJUgLVZ
SE/Qbl31+1X+mU1Zm00btrgkasPnJihNuqM3e1ZxkBt4GNmWm3mOgOVZmL++xPcp
qFZIYPaKfJLIyrNpd72NHUJ+28sputE7m8jcPCK4HQBn9MisRLOmlbQlReq6i5oB
yhAPor5YR0izQ914dptwUfWbr9pHBlDMHFlHZIjGkHSNmgDNxitgRnlIrpEmGgTF
AIKeIXdAq8ukqRS2/4cQEJSwnyhPfCf0crKUcL/sM3JO+eWWGajmrQKM4etM1aqj
eFLJi/K3S2c7hsIVE2UZn8XldrZKU1quflGuECiReTy3k5pxWmaWkOYnYjKChw4k
LI4kjhWX2oLw8iYeovsoKPUyj0Wvzs72yuyzKVrULOmDntCMHFE4dcBTTBYxXab+
BTHB2+bWXJ5JpKFo5yQNQ7PQpl771ym/XKAOmNezaYUSDPcfyLXfacQLPHTyzWzu
karimA75FTYOFI1poE6TMUJAfTTcorwYSs11ehubPhbNBr5BvsegFz1qZIdEvaNd
nEY9vxjmy89sIUg1UgTTUgxvNWT3bID4yy7GzCvHRoXVWjjlFrfjf6gCyWo2wF+4
CzC0DUeWPJYMy31+PptvlykUtfhsjJaEeOcrqCW/697wnwGI3HS0dKh3YprDN0cB
gD5dtDJvLMb81lip6aJvH9LWZzEz1TsB+20tUaRy2df+oDQ+q5yt6W8p02Ebo11T
cizSJUjdkkHlwzVLBzN6s6BVYfcWu8sra7x0m6feWiPLQtjG4Riq3cVNHtJcRO2y
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RH3H6PC40+7cl+p5p81ANLXLYYB7QjA81Z5DlWehTVVuDD70hNMEOHKAxl8bTFmp
ORV+kry3WlqVdd4mjkxI9eEpJcOMKN1tynjkNUGXkKGD3jNMpTPPIws2dYpQRWRs
9GMZEKO+54gEuzl6mYDyuIVqgGXj1UJyCWZrFOsDI2KMf02UglyFUgwFgiFSO8ps
czJas2osw65PVSeQZe7EJCSuM7kQj3tfh+qgQ5IOHKn29MTDQNTXCYz6qHvJuxLp
7Im0k8x4Nfi+lSn8fbgO2zlyKx+1gkd2j6xGhp/TqLTyhkuxJYtgses6X6XCjYRY
nUauBxhi/4rO5pyKTzf6P8SFFSabz8mwdnQahgj9otvoEi59LxL0nuNrqNwk7ULH
q1FnCTjeCQCNlgEvWyejGd6WnsBGU+3nOdesn2SOwVwLDn2KhA3ZAjtp7/BziMVx
uNLMaCMFg+3gYR149iY+3XVvgUHgy4lbuqyqzg8+VUiSRW+9Egv7gD8olXso7HfJ
7kaePqUAr6e7UCXmlBm6oTAxopIUSchGUqcr9ESuqGjZNdNailOYH4/Vjj0FZIuI
lTi/Q4FymfECH3nJM8QrFLmlExNfda01LTGwypiAslXnv6/k8vgScEtkz1mrEkwg
QaPJdJOxvFuC6bY/jpPsgHstEICGAsw/cpkl1mEaCVaEICQaiQp27AjIfHFpD7X4
nFWU/rFtTu/Pv5e9olJABQXBDzmSrJQ8NSXTZ64jDJwavO8agZUvNN33zfDKrDQH
mz2Ph3yqhcWjReLxRwqSsBecUlx63U1upOUsLWc466rJgYRx65ypZoagO9EmDTEG
6C5XcX03Dz949sRzrQ7G2cIk1JirRi7kEjzF4pezckVVDkUMHoIACvacWHKVt9zc
Fmct13RM4FNvK3zbbkDDbeU4cv9H5ixZUJW0udA9jlIBhGW55n62lEW+RyRBxFcM
YInLnHqBbOfmarMN8zVNjmATpyaSgrRroDwxGVQTTlZzxovdlP3kLhitYW8tJfnO
NieoZMdsWTf/IxkxXEKe2bxTyFEyQkt0iN62dMkJRmSpLNdh1yrRpVlCs1XyiIcY
SSZKVkN+kHO/Rgd7sU+b8AyYGs2azzSrUL9orPMf3gXIKAJXXAfaGIBUU0iE2bsV
XwxI/p+fV74DXdd1/ho50QqPhF6ArM3a7b/P0sujrCedEbvWK74/bs7Azy9O+9Su
SgvXaD0dlCBqTS7hrId6eiWVVhW2raWwXsqVABzg6CkVZngslaWZo+PyHT2iYsq9
dqwUSD3fSyV+x+xzsy1F4x4XNrnru5orojY9KAbbGIeuQqAsIO2M/XWNPeFnetqw
CojJEn31wNgcGoKJsLsimwpBonVUVu8sIDfssuTyMGrmj2xhb3x9rtDTCOTK7oIR
rDCRy9ePX1WYS49f5SmVybr0Q7OaQ2ur8dn0jiVW0AjYPqS4Nj3DhYr/8WcalNuD
WNtTue0orILeGA3bPNVT9WLaXIvhgT7GwEoD08c4HgMTXrX9vfq4FnTTg1dQmNHW
PFXx1QHXSZRt6E6cWhkCtvHTMA0Y30nE69fA3+O/LuiT4MRR3zrBSGSd1TB2T40J
oMRQcvi9KL5aTSEh0ksn0eeblxGO54KtlnEBkeQ8VY+3vnsvnbSYmXcZC5PoNupk
CAQG14VboMO2ExQ1+k6AWVB9E/6iAHACUqg/tSIB1ByLhOGywobXTL5ss55XSYfB
ExXBbqwTijjiT3Vt1Ab2m0ZDP/j8Ocg/pVXiF0EIwPwgjeVCoakgSJHXqYmzt+/W
ho+E+iJM6hwxppiGT2c4+vxBN+BiE8rup69o+pKrDJDj7uNtXsOv1RBLDmySSJB5
sc5bXFspi0sjdmAhibSyjdzdFx3aUcqaI0Wx8BEkmu/Vaqi3xMQpQ3n9mykCo66n
a0tom/hwNm17DhL+jE0YaGZE2bXz7eOTnBrkoOskSb+QlzZFT7UjKbnTDgu4VzEn
qwLzyJ4ONwfKd+NuEN3aRc/1+fwY/xZmBukJK0M/uejefIlOY6cD0ELPA/74eXgD
uQVJ+cysGD8wT5fTsuyoW+Nh61oghUzXFdT7V1u4+FmV08fgXZgcE+StLz1b2d4g
wROPYf6WjzhdMiFEuIBfhWXjyNzNjkqUfcu6l9K06Hbu+eo/NogggSN1EE96zhVX
aysm8JtPOcu3bzjm9n3HL5Dq4JnbuKiaM7JXahjsamdPrsyWqLmUcHGwNdrN9kt2
AYPkYeC3etsqWgBfyvUrJPXDYn7DEE5OvO22uVrLIq8v+NHe7Y2R8Iv4fntsIqtv
HPTRbchPEh1ZZWHd3vUHEzFBdJoiLz685ymZQJp8IMmQFVJELAQTmKyYHRtL07q4
dhp16wiGKVlVCcTQoueLTG3+iRDx7eqq7tL7FVedIDowi0Wbz1K88PwIXlqnN9dT
Jj2QCgL/KH1JJti4Ft1WNwtR5Q83GXQYaOiDruG5Hg3NyhMbA+LTWjLW1mTv9vNC
LzNiwMzZHLaXNk/V7igCryzkSemRa4N7YwKyYXO3rQjWPhudkUcx+Vaeud/VyG1M
Rnba+xJbOIyXqc2D7O3d2TR3Bdj7ObJMwGRGZ/crR8MtuL0mKm1J0VxD3ztpS9OV
b3FsL0Gc2vRtwLzZtPMwuWuL1xBN3bPmhgrxNHm3dn/3lHN596YDoaO9YNb0DXVd
bn7VqD8krv/FePwHQyS6HXllQUTMKSE2ecNOnd+xx767GKU9fZQtb2ifJpWQz2me
kSi31zqb0ipjK00o33p4SWDE9mQWJCDnV/iCtePHhCeMxllWhG8/SWvye+KJNDmM
ndAFo5gQ2y9MVPkWkL9/f3EjHzBg9xyLdeYp3CFM457Ku0h5htfEyJJplcUEomvP
fHvPbxVyuOIkYTMEAt7e8kjALS2YmQ1iHGZ6iKmBW6DjDpo5kY6ZDcewlAnlW1Ju
ShU6hsbz5MxPGM3OeC4Ugj3UgHXZvyIe26eOegMU3t8w+4Ylgi7nbdz0hcNpGM4Q
rIF0QFLF9td6Ovn/oajQN0s4rJ79Ds8V6G1UKS0YaI4Yx6sMcyZCxf29vLltOTZc
X/Umy3Im2tUaXHiFpQOdF5yXYPW+V6m+MKIcb+dWd1IbAzlEEIjuSElZqytmWGex
B2uVKQEKkGsywJ1VipK8PPBDpMVzY6UK3RNZJTWTAKE/8UZLD2piWX0b4KIH9Oam
sJTpGimxFv/i+zSpWW8QJHgDop8WK0sTyRzF/YVefotXljeeU2fQIITHXXUBlZAL
zNbeuXEk57kERQnRVvHZonekPAbqcw9ye6XE0jN+AuOfxRh6I5oGmfLN7MOA6S1y
IFnbrX0+pD/TKR8P0gn5rAj+lzkc+ZLH70UFLU9x+iAwSUOc4e3+2hUzTUky0TT9
ck1sC//7sc8pddVTk1hKZnlqph36zZSXIjTlp5cMHRPabzUsDkKfT/3av6FjFuVd
rbSankkMwqeRM5MIFmZidC4QOx04AFiDCo4hjLLmOMZZVFMUdCzhA1v5RJJ23ZhK
W9CeQFyKvOw5/ZR4AZmZ3BaU2Nl7yQ7mdJ7zew+63TfH5K4e2/rb5i6Doc8XcXIq
05jeu35eq8ESABBnk1xt3PJoTN0Kok4Gulx8XPqDyq9MRce84CPLLF7WpwKoQ6zQ
XTBF1qw0dGkw4Tv2OybzcJl/SoDYiDedYquSh5UQ4Ll0UFqpW5DxdaQZa7PoVpE0
FKjavktxtGuCNOlLj6uy0OrnXQBT0TbRhNeqgr4RqHVbJQIfJcOsdZtrkSGHtO/8
CacgijUMOBAKYLMXwG1In7iQgmidILhqgqZxPsCulBUdkpvhgAFTjbCoJpiJKkzc
Sl36XvbOr/x9kRM1OYA+3mU3AbE7THdeGP6zTknrtjYY0h2VNsKyWasUYZ/KNjSW
GZ2qZRYxnTpbvXH8z1Ly18boNOYSjOoCslqCkNZpPKQz4egpUtbCZ2mGwAZd66qT
Hn0oBKY0hHDYepuoN/g6r95RABIEB7gfa4wRIBzp/YsJ3iy+wljYcYxwAGlT5OCS
58l0zb7alTnaKEl+DdcX9baH1acwJ4MXFJyCZQrfwhXy/f8sKpj1oayfqCoaEFi1
1nNk3VNCc21qk9hJ/eU92StwzWMDP9cShLEoiIv6gIrCGQLYRV5BFwBRZfXhdQhI
JO+nnQY2kRNxI3fSq5Kj9ttcTobY9ft9a3wj41mnxQEjHPlurfyBmenuOIE12Uc6
JKsZ2qk+Y5fUIuE6ZukqBtwGAU24B3UJIraCge86wKTZvKujdZmnmyQV1JuW0kgK
RwyTE+igmmrBJRr+l/Q4e05zIhr4NJmzTOyijIn12H4ZiKmZrSwS6aQQpcMb4f5m
M7bCPl4Any3zhf9a4tXl/YwAjG557Gp7mVLcC+3EYsFAgy/AjmoNZI05PCWTf3VB
d5vpqo6OexxiHZyKEr+Mn89nb1+1G86/AoDEgDxyvFubJnrbPuPwjpsQAsQsr6Wk
/C+k4Jxaz6j/qAqV14slrvGkCzfiDQzbkW4KmCDbLXbMIBOZnZSf5Y/bW78e67gZ
zQDIQ0TbawmYDNRtbtPQWOp8Ep+OiQbeqO3vZBSj+VefmA4O2xJL3ucv1U2Z7x3M
+u9RFkeGsXxAkhP2lHxCAAqMrKUylsIJLzhvsSUQqOhAuFVFeXChGlnEHf+Ok7vV
Ut8phjOMWVzvRKMFiutLcwp8pfyjipjEVM84ggzI5kfQ3HOqpTez1CvUT7+4pJ/b
EjY5/Xns5qwDxtfpbK7+bULvUEZR2WXI2TZhf+3ySmjI7qnsWa4zTrYyNtcrX8Nr
HaCu0SFQK6CAqgyrecIcT57MqIA308thI+4i/BjSt3Wp8JHUzyP4Sb/U/TUSfUBI
dHLZMWnl2h2N/bsEJY6RY29z0hpP3/GQgGSv4a6MI2Q9PD3BnD6sX3sESsRRgjUT
08vAsl5n8E4dit5RdYAA9bLGS9AN3dKrAPo6FLwB7nvmqlVynvYiJBaqlYbEr3OE
0YMVNi5zAjZ6E30kp1/n+1MHgzS1AjKAlWRpHQPseK6uwe2+TsjEm/tLmj64WPF8
HVicYy2BrZUYiCvtCgviRuLY021NvhaTpV+bPaaKGCevXjhtDmH9RkdZ2iZByaNi
4XYApQ3+0FjDfevwZ513Q/12R7wB8yDuMoBkPXz8oHNi5J5FZcwiAfxg3oCjSiOG
glVdnx8LM93mew6tZs/VKx+lczv+t/+M0XkTZTSzWDF2hwkbzCJmJ/dsL4Jg3pwF
gMoPd1lkCOai/pJ8VcWa373dGw6lY+ZgHM6nBH+BxArzYOvmhn0Baj/ikur2O7EZ
1OMlV4E7CPp7CqIY6RGqRNmxnXk/DxOC5a3Kx8xd3V6nPLl1RDT7U9F7S1tpIIKn
GiGSbykBpQ34EIIobWCsArBdcxZulkF8zwQHbspwLs4yJMkaya9xLODscv77dSUK
d+/WzMcz2KRqgSf0wMpYf1dHqjtHbQAyYwYoyDPWcUwq7KPFRrjHfuva2g+bFiIV
j4d5J1j5QfbfJJVqh4YCXHd/UtIopbe6ccv00HH4wb8Vtp3fyzFRbcQfNfZ5bZvi
R3XZEX1yCB5kRhbJn6y+Frz/peBE2p314C2GN3hFdqEeiZGWTLWvFVSjm2fL3lMv
vndppwyiixGR0MMgbvFD4FmUW41gqIX7J0L2bBmNzLtWVdvM3UBe3YGIapiW0wGq
ewqMLAQSpYyV8/uZ28KCCVjVI2uBXcJJduRkgTFOa80Pq/ak57ILiSxYkNaWKses
8+qLjDGa9H8LimQPYYFUkTPhgtSEBuvBesindKbUBU78kY6Uuobs+YY/GDxG0Mdw
fbZ8997lW63jlbuotdRYBx81PECqviNJ6OsXhrvdzzgS+VV0rUMjJ+ih8tnitpCF
g7HpZ1g2up6ckqbTZCTpi+freopBAueIbCjP22jq1AwMcT8Rlt1vV6ygI0Z8n8hA
2unT108FtPk4kJq3UNFLX1OBbAf8Y9/rJpd+H7G5ey+FFNHWGYfxn6If6xb7G/3T
/jZWBFVv3h0xogi2lCvtvD2mUKn4pKPIBFn6Fq8067SuDQV8iP107/cJxxNVTJoi
LpaG3B70Y2iOj5drCOC+1Vobx53bLI68+FE+nFZhwC3b/k/aTS9CE83m83qSUu/n
KuucflbkEUFeWjgm5har2gqFHvpCe2xaw9NBv5VtjswCJIMumd2Z3p/MFmAmoh3/
ieeKixu3NxNFyjPrQAHN+AeYtRoBKO91l50hK23V73jrwN6oiTpCVO1jXPOV9VCW
sWUgC8V/DLWfseYDVKeNEbqO550EBlW6H+F6e5/30HXIPTl5tGsj5XAQtGEZhynO
/RXtgifmVXXkvG6fq0ykQSHA8lWVN2F0MBosX4dNHT8Wg6wWtTfWi/sMLPfQtNc2
eN0b7dpRtEPGhTlZRcbfBK+2Ud3RmDDVWzwZuambtXbJ2KQdu1AIqi3Q0yl20mci
IeTcmWSvomvU2S8TrTtK6iWxwZGNsx+xhfo4lECr64e1Er82IwhocOS5VlHYgDiV
gYrA6dwbLkD4dCQqFvI5k2UaIemaAMcnE6WaEAIgmJWS9u48Rtj6eV3BklYTyqlR
s1bTr6/pdSgsJe31lgSNKukH4YWtywMba3rC4ofMkrlLDT/I7/Yn1BDRF0MLNXLz
2UstzHQcEm1+65jSLSnlyqYTGbPWSVyjXj295bRiKEXC6yeyhAH1m0+yiT61CJnX
Z1WC0KZ9iMmt7tOA7sFl0vPU7OQRjuBMcxZDV6zXWwK64g5rjY2UmqXH148pZM+H
ka7Jq4s199dWO9aiaC5jkMBBdsfT0wIJs1eM58to3J5LgTwEa6sIDOo4wbKnikyf
MT378XuBnhd7rqS9P84qrFKJqirkdMFOweoVEt1EpkUVCHSHWjSpaBygdUARYNMc
4L83gHsoeYNvHnG8iz+tNE9/Mde7dJ1Hxr3Dxwi7hto2WtkN0LrR1WboyaTi+yIP
IfN24rIkTTHvpUBrPOP4iHr8xcIBU48Ns9La8K1ma5X8lo5fUYKur1IJ+IZXEtXn
GuAWH2LW+Z/G/d2RK8ab7fnxMLVBj/DwUctryc3Q5d5tIR6T4NqLmUduADj2JSem
sIqFOHvKv6myf8G25RQKKsZDqOnQez+LzFfmWsQCChkHKhYc1SM0cRqkuHY70KOV
Pvh30/WJ/SyLhYkDqbNndXWPlmCcev8xzfiaakNwz6lVY6gk3dYq97hDuVT4xKmZ
UE1BSslwQVHi5YTE43pqdYb6j85YijQ/TPL6xEGiYgYwYEj9xaA4kdASj3PrtnOO
wcL3fqwn1hsYz65Z6p0lj5SXOna+rryqJTMEgTMH/04es+vuAiXwCEYdjDFjDfUS
yJCpF2kF9EeVt71lwFm5XSZ9+Q8OzlzaEjgI9UC9X9lvN5YFmGD+7W88UggMOwDt
XrXK1nEzzq97k52FL047f/6eYd0rKQa78ln2Y01K/IgWKBwWhE5XI/8RT0jkYRtC
OQVy5R/AGxiBvCNqKXSINVlOZ0KRwCgNEMl+vQVie1bOJfTb4PWHkB0cU8BCZ9Ww
Lh7yrhMEEvAH87pLAZ5CgW4RgivW5rIjbxVoJ8cx8tGXwxYCjzfuFu6NksiAVqJD
rVRDw5NfYuF7Y9uhtrAzzQs55RK/8qvIOcFpp9AOunZ/84l4QbK9LITAoIVJmfxc
S5O2XMNf7J7nI6nptB5MjtGtnjqDXYwBW84tKZq6u7/1NIL9whSQgf42O8AKHy05
ILG5iYO8rIhmHXyenG23IIZ3M9bkgrcQMGE2hR3lsPfWbFotapl71COfbs01EUu2
S+vWj51Bd5wh5zpHO2uvI1JEvFMPVSbYcnkgeqOoqkAyAgAWs5tE0bxB2Cav97HC
3l33tJJG9SSNP4SfhIHK5BZ7TKrpGuGZFuGPKag9nLRvVALltLSxXSlxYPeILzP4
dZWo3YV35WB/l3f/7qBIT1XujhFY4MruMssct45hmzF4+tavaSEi/mjUxD5vGTkO
5O6/rCs59N1ca9aqJYATq3uTxQbIqgSZdWt9IyeDFXALk4Bxm17eURKlQSjU/YsC
xQ+XwEaMUzEX6VzT0Fo1GvVaamEBvpmwBlq6PSgGxjCa1HSHXmk4z/7EzDN/fguq
QdBvJG+81H6vcybzRGyyN/U5skpGP6bIBs+PoRTPZ9hiv9rid+nX4b2asuufq7As
ZPoVhkQC3kAHx9kiThf6NX4bv2gRA5BZt3d+YzCbL/z+ntGDqrkzhlJ9Ok7ww+em
7agkjE1yyfcflztdQNCc7ipjPfD5rCLywEC10Cw4P1WImdTlFrU14OejNuU/Ec1j
XsJDJIjJD5HHnL2ztD6XQFEInM0aQwP8zOS5WxQOEUlfMR/SnWDCZDbSzaA8+C3n
FelqMp0ZR0Uw9QM0s2nkBpFESJ7GsdjIGQXiOo5QhLRtT0dqU1N/wDoyJ2NXse3o
jfxeGoKArUq+AXVg2zT89SpPu1piqWFrRUEuc+mFUH+zB2ZSH0gZ4Uxj+OCx7SuX
Wf0G8ZJMizzREpdnhjgml61qKQ5vDcnxQ0j270dgu6HDdTjy00HWsXPCIErO7bT/
3LMxi/fLX5erm6Jy/AToCIu6ZlCA/PfAwJem3CdUMH8aVYoVu7ZAnCxFuFDXqkfu
mruJUUAPWLuAO82H9sldvR0gz6ZUIk3Oo2rQVDPv5EWDZtp2y4yVsdaNmxdx5Z/4
gEcSeRm1mm3PFLCBu92TRxii3tB1W/ZiwRkKGKUgFPg0LE6txKIy0mnuJ3jPPpQK
954QMCeeqb6zgwysdlPdM4wFipRWkadU4h/0gHbUqzYemcJTq1oBy0OpVQ7NcV1u
HYKF3/jUSiooXi1PvC3VDWT70INHtnEKoipp5N+shOe4XgrDGMy3nA3OSN9qpUzr
vSxAqQJ8pG9Q4Be1U5eIgmRJrv1iLgMFY1gR2ZCi7JBetMhPUl9/7GrvWfdC9AoU
5lQYWyAfABbDuiPTRryHnqELqnXfY9zkQoMSN1i+uoc+M5zynCwsqKWBrRTxXM5E
QMWLPdPrVbacXyBWssRoKMNPjgcNam7J6Z6ziDYnm1v7lhaDh3GvVdj3j3ldBOEY
6GQlmAA5T6kmyEvHMn/IKf/Qqro4klZO6WSCY709nqzIz2lQUWJdpHl1ou3M2DDT
uV3Kh4eOQ3yi2XP9H86O8RwqjhhtPvMaRaTzkrGCx1GJiAckbnMxTxCHpbLIy8CB
ilZ4s+ytnryZwex/Qf+tsolPrgMt/R0OTZy8k1rBYKnuVkHT6o5ogSyejeSIAiC2
Muk+FSCqDziu9QmplGdAnaqrMMjAHuPSbecgB+S7wrGxevL2agB64SLOOc/x+293
9f7XSX5wkEmPDfGisL95yqtT4HvTg5U+6MBmIQlZB9g1S9OfIN8s5fm7vHsilZPr
+XRiC+BWyDQv2c4EoNfr2prdFzzNLh2dfCxVpsG9zzV5Pe9pnE8qF2KKMmLXDi+p
o1jdSYYtoI/BosfqZJ6XG3q4RdPoy5CCuoYWPRz0ff1ZADEBAo9FPfDBdG96RYRt
7TuaRFvM/eTYSpNEj89ybHZswkzE9TPpaa2e/O2ZrMRP7RfHIsPFEEU+ACy3erXa
oQeTjJ5k97xAiO58Ov38YEde6mnDI3G7OZdrwcJrklzEPMjSY5Oq4+Thy9GBNpJO
k20zFSq15Qa5sOAr2c1Y0tOHTCuls+8o4xmkH+Nn14bLhd+qhAxHLaOvdITl/gLg
Kh4IZIWHbNj5uA7JQ0gSp7mv+sbymb6X6/hgSt5ZiJS8os6GaEkDXgnlOejyxKv2
MQRz7B51dKn2JG6TD14lN0lJAlPgDKPy35YXfSv1qKYAVMLNXITvtP8FplNMocLz
CN5o4JsMzjn0JAV3ARWJXdlzLb8hctIWQuWhSiIssw1IsxxgoaFjWFI5ZHpnmQDC
lOC2unDqsDAVRC9WVLxQAFejBIj0NgrR3GDKwN0myz77gnaifhd5oXUZ96sm6Ew1
IaY9SA5T/EH5Ws+SjJFfKLiDtWFeCXn29HuPvljq7XKn7XV7alOTNwYHjZgNDh+G
3ogcRUa4OlETuqSNUGtK8sQ0X3/Opjc+gd4dX9boxkTJVn6ggoDXWX/FFQVk6ZD6
cmVaxaNb6IEE1T0p752zw+UVyJciM6PrW9yGEPX6pwdCLcwpdccolINsDYRE1YkK
JrYt1G23dToPfeWPZm/gSV2Hmwr3f2lEOWWQvdyICL6KUdZvN53Lc/JRZ9WH6ZEE
3Op+EtFQNL8Ds8yC2Nbh446xgJI4Rcp1i5aykHE3p8WSKibPLNsal3DFTSnGdNdw
IItETsR6fPXccoZjih79wHegF2PErenvNle9dy1nJSJg5U+K+tyMB5fzGdL1qkdZ
HHILQb/VJLaf+QITiy0+hRaEGqGtZbFQbnoAOMbGlRIwS43JajtH7mbZ2pFxzAMd
VaJYHuc1IZ6ll6AmxiX5FfuehgXVE+pISVgt1INiWG1894hFyXppnaAeXslFAw5M
fQwUZA0K/bJMV0qOi+s/PhkXe4kxBuGVlaEMOjjxh2WJEnc9WVfccHvoA1DjQXSi
n6noFtFfm+aY8bQJIXAK4OS23B7wXJ2xGGCFxLTAuEn2mgfjqqZDDsCyuGzZIpbA
WZuYABRAZknc3XoqN2AaTfa7EJbc+msJgaS/x543eZce8LolrSMk7rJsLURU3f8i
7IY+Vg4gyuLo+ZN/d9dfC+6ytklcde1YDPoIg3UfJgdha87A30WbqyOMemWrVc8X
ItWi6p7LriibC73/LwCaX3GywEGD5D41CltfCR63Pp+FuxvfWKm18NArvtShfvaf
Two3O1I0D6fzLLNqTfj21fbA14lzyHGpEJwdPTVQmaxtYwKBheXTXpCNPNZefYj3
AmLTKQCEMRbCukAgzyuEm5eRgdg/LtGRiAwxGgvUYtosRD8tRURL4s8LqoanCHTl
DH6hxWSQ6EwFqrcxYK9ire1Lyn9SjyVBGmM9HCNTobLCjXCfZAS9rIhYADTFgS3F
OLv/XKBnSaFlL+ZD4eM/lO+7zOX9NxTVEeo8S+lvbIy7S0fGaht2jIVmayXLiv49
MKkfp2V+GGkb3inLYiswz6CZv8TeSKA9cFug0ekjJZJlphyl15dZJm6sIkDPc/2q
cFZtdkUcyX0BCaJ8B7+6Daw8ct+5f1cOnBMsRTnAaerDsBCUAgBs5H+yshFbe/3a
MIVrFvVY1G/nXIcuB580S/J7UScVkfPgAv5lnl7MB/Tc2ccgkrMPRLriDGIDmuOB
piJ4mfh1696jPhXb7CWb8RaCtVioyy11jcETv24z6wj07q8je8vzkJCHvWlsK1k9
PKOm7mmA1v32jJa/Sz80KriBZEvku6flbehgl1zRsMUIDFiiosyNwBeAyulSVprZ
Lkr/e7PqRS13+hPthezdPN+rXPqaJu9nql/dc23eU73UPrG15f1mxXkIpeYqFPrY
Vt3WYJvNrIj+HDfXyCFOzM3If+H1tUFKzMTR1umuANTxFoTJE7lCXt0eRRjTiu7R
DptaTVkLzv6OHGbcsjOHfZCD/52/KkSV/RYSpT6x+Qof7UAvA1Nhl6PnrTLHlEDR
z/564YuLxSdj6GTF2HJt1xIya/upv3QLsf3xtiBJP1WZlyUHe1WH1GO2tMIoCZjE
c7MDIZpUQSV7E8tSG/wFPXMhDU8pOxVxKPYjU3xBy2pJGV7J4priZpxX3X2MxRcL
Dg5xPYouXWA+KnmXOorT8gXUmxt4khizAJZP/ifcY7vto0N6gw4ePNv9Ac2Kqnjg
Wf6f13sJzsJVCvtkvik1yLiffddWPmQKfO7tzAAsaJyAoOOokgF3J+EUH2Hg4lqz
rUhZXrhOQx+vs/HcJNqLHtbUKHRaIQd1HShTPiwoiKK4URfhFvh8y4/SOxtcL5SL
KoJcl0IuCJicPk1+bqk41hXxfPn8MU4qgDe9D2zTy4jgcgI1AMqcQ9zAUuVdky0e
Dle3FkgBDAj3nSH6uALbCULP4bQAgSMnTIZDdjqm8A1En+EYjJkxdW8y+3mZ1VMC
ZZ0jeyZYZxYr0v0dbEm4yBhnspQKvklxZcB5OWuU+S4gyHNY60LQ9kd6OqU5G3fu
p5Z9bgNXEDFB3WA2aaTwkvcm0PGO8z2u1cG71drfEaSTcCPyWgn9V0HQ+Gz9m6mi
CP8Dte79stHn0d3MjJDgqqbhKCCyAOE8rwmzHQ7hTaFBONgQZx/0GXx+uHXoRByb
bxT80SRr3Xmk2RL5Bj1pOOXQEPOUBAjsLDwkpZx4XdEFgI/T/SawuNVDXSJZg/YB
AL+2092Jf4aEspMR0rlZyf3vff2JK8LxP50zc4BARVJ7+K3u2Itj7DFPJQJUbBZw
iqq1U9mlnSqXewwnQ7lzcA6LMqYTvsN7CSiv9ZlSOBEM8KIw36Ff/J+2mj8yKauz
qPHcu7wFOCW/WUSIrThWssJ5PUvbTaee/bf3bJhO8dklsDsKT19+S1aQ5Lq//s9R
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rt5Uoq94NUvndQpV0RI0xa6jMStzMmG61glGyWnzt+ytkML1I6A6G2+h+aZoflXx
kw9gYmuRhCSVNJHk9dW70jWmo8GmY32GNjk6h9DBYKrB8RbpgGLfMSUoS0l9PEjT
FDEDKj4Jc+AB6F2IOi4nxn/CKVIauF15LC7D4iepfHpGOhIVYZ597gVLiRHMKJ3B
M7tkKG+2pF6xhvw8qkNacdrnT2m/cuzzF73/Aqj+MG+Q7z5XddsRMPYpPsx96jQz
PGHaR5STaB9wbKXgelg0ZRIe132yGBvo/WYySJTnq/6ZzW4IckcEBqcxVG/PknQT
ACj+hyIJ35K60ZDIRHIMGUzDwRS270vvPeP6E0a3+vVJFMZ4qcerePOcqe8Xl/tN
RcCAF1wEMA2HDM7ULwzqSFpNpXiZ2CJUxeNOL88aRGwHTj2Y65zHlMuyH5wyOj/F
sh08YiwOJB/u48HzrCzg+j/EWcKQa1sVnm5Bkp2gT1JvmnNJkhqcjKgXcdLPkz5P
hzK3mwoaUOlU38MDWBfnPjkTy68ALIFBtKEj/gMfSKANjtVEloEbch5hGrKAaZlt
4bBQ+rNFSB1Exyzir4gdWs+jxUGGCmpC1kChOc8ITVHSTLSEjGh5pQvUf30alL7d
HOKsQeZwmfJOqSnVg8oZ90w6n/YcCc5027J9I0nmsRvQjW2vJjAewJOGhQaDfi14
ZmUCZFnCb4Hmi3TQ8Yvi7GDbuLQUO+ZpoiNwq4Rh6quFnul/UKX3YxhRWQ5F7mD6
r8v3PhAjZWsRQ1BNMFJbBWqO7ZnQJGpYJt60JBQ0HPGB3a/UuGEnLJQfQ1CPzoEO
h+QTD4zvYWN31ul6C/am9G53hZXK4lkUiCOBoR2x2P8YlG6MPpoyATN5eg8q9A3D
+v+ZtD9uj51wXVN1e/yP29SpVlc5r+ts8VNHWHNYwaN/Y/bYZKUSuEPCpBYaoiro
l5wFMN/j0z+Mv2c4W8rB43gJ8fOSR2w8+q/ufmGS9vSsusAKxTpPm3CRS6evlh2Y
+a0Aj2o6wU+aSaB4N5hW61qJ2zAyzGI0l3l2ZoGl4Uxp2ekBd21SWo9JyiLnaxfa
3BM57MJLT6bQsjm2Ec3bED8OBZAnUFICEolmNJB+o98YYlIf26TZm73mAQy8lSDq
PEayvtYaWdIzaAWM503TFDiFvzrL1IfVIdYa+ujdHX5A0preSceqS6tRXT3AEU97
d/MaKzAfEoCqx6EvjIaT9aXJfsX4GoLttYTEI83+L4tMPRW3UdIhcyWdjjaVnUFW
s1KohM/LxRr2R7pZjPvYV08dvX1+4dsOTlBbL9xwERNOZE5cmuuw0joZXdRm8/KF
W/9j+OYrtqTsT5KnIeY68eDI6LAjza6zlr9cqARSNMnCOWhZ5N40pnJsrEcx3tOp
jvDSDkvtVxvbEdE06cmB+NH8zLWcgu9kM4D4DC3wBcEneb1IwbfrZS8iqWB9g3mc
K/62Z6TUm3o3eBF51jhdHV/8LrTxddlrjrL2BrzmxcEgS42mYxyTMqR4xmmovtqN
bq/ubncdUrziC6+ZKuTky5et097Qz5Ei+JJx3Eb5L3a1RqUd7o/a67I3IFsmj90J
UEjMt9TAMi2mZkUauCnxpEKaMo3JRalEsDzZfCW6ixLwZ0UURDXY1dwl0+BhM0v8
uTUb69WqmU7nPAXqw2NkIv8VRX9SQWO/EwFaEjjsfhRY8DBgcQVQbIAY0IA+Xr+b
Kezz9XCsFYe6dNBUDSs5FsSoPB/IgpnY57CG6EajNxWPHudL032mU17SJSOsXa0A
WOqmnsghQnWG64aufapSSI7RgR321aNDsRihaE6S5QuhoJwUmjfXy4ujyjp6dexu
JgoW7nnfK42nYU40zvKhecTEo5mdRf4n8UJbMqNIKfKUaRuG8LCxumRZ184FYATJ
FFgXT2bWRxuj1vTqn7JNVKGdKu5iY1RFqUqsO17slcCg0LxsQEgrfdt1MabLZbAR
3l1gbWAgffUs4bkmo2h8PuMIYCDDCE1JwRFF9tsyD6gJ5xxDVkFMtFTa/X9x/jUI
TgKimN/a+4LEc9tJc+DGt2Zkr4adUajnyh+F9pjND78LMXnYes4269q35ksqaGLf
ZIWRdFQ0wIsodMeRJy0XrxU0ePt5FGPyK6KWrMoOCT3yZ99Kgql37Ghwz5fnzCrk
Fo8hPzFZgt0SU/4mj4RrM1b34SD9vdR4AkgEBM7I5HYdBVzPkAsVtcRfEyf23FD5
nMDhA6LuvyoIv0fyvZuLpzX8kvIOV2Un2lt/k+K1q36wuNdT02tLQDZeK3gyJBXn
H44ygkmCFxOW2VOaYjU5RwmzOCJL7IZ0X0c/LMisUODRoHPaHFRfRoJ3pDFs0Nhk
xAyKW1bw4SyucI6wqAsKJ9VUZG8quONXof7Z5Aq0M/sqwUNAsq5ZEcYIUv/vDLlT
NA7uCAloQ0/AlBYsA1McTBakeT1Q0VSdif3r/dPYnoQ/6+AONHzrJzDEVpwSj0t1
bwJcavJZnA6mdUES1CoXFcYAaqCvHeJpzFjLdYWqvwkHc4R5xQXlwEhIioPrDhoS
oSRR6t49huJsp7AbshXk4FrcylnsCVF1MRT/7s/ANWqTTYJEdXreFugXcDlbwgGT
5GgY1Ej3+64901BqlqLW9jneMuykyMzdiFAQnNNCmyDp49YyD8nGFDC/jZLG14mQ
1LhXP+sPyjWK7OqlpBSXaAI7gSq7OY7zOiXlqPX8gUJkjlgDyKSxNRszWkAlywik
zz7S+xmv+vQMbbaQ6SxvpXFuUlULb9HNjuOEZLsnz7GioiLkzEiJeJEV8hyaxudD
7xhkQ4SYyZLqDS5Bi5WdZ5Y7L/R9bGw2pjZsKbEcSckKhnDLq9tI0Z0WuX6baHDw
99ulF3r2aBT6cZrciKfKGs54Ms44jyTeO7t1lqKnxqJfsPCovSi7lKGbYA0cCxZ0
09xu2QXek9ma/7/CTxv/TlwvsaDpQ7aumhlSHYTYNfBP7jUO9PpKBDacY2KtH0U8
tNKB0nQPKUUyy8N6rgm2AO//u5aDbehNXnyNTa+usdzNDS7GyNNB17HjiLGFfDNL
8lpqznXSZ2a7homfMc9e9P9o15Nv+is9PV5o9kKmqknE7oN67guw9AqqKpsj2CwU
8zxlCdDUsttvphcg/HhY26SG9VCZcTfMxp2YqXetM187pfHVBjIIRl4dI5WByLsi
NzTTTBoYWSlnQR68DXI7KRpYL4xlVHPy5zVaJcS6qRXHjmQRvyHI4Ggnu58KpvHL
eE98Q8IH9eZq/V5dtZZQAv7cpzXwcLVQoo/kBFquUJTaITsMSczZ4Sq1ff+SBpRL
cWz0O/YF+qhBRipmzIMX0wExtv2ky/3u1JPtx8ddOAzZDa7kmEx8M/BH1We1Bunr
n54zUZzO8LrQu8OyF9NIyn1+C/IxoWNQYmbWvPNeYClQAXue+A7iS6q2JXWNyz/D
mg7imUGHfcUbuTvJBNedrPlSSRmi4QjDG22EW9bBgGCG/FGiAZGV1Jy9Mpdq+gQ5
Haeh3QWQYTn02IqPHtSP11A9InY1/9oJrrWlshIrF9evbq64aNDSVPvXwhXO0yOi
pTah6I8AiUtJ6ovNTOIUsiB+x8WaYg9djvFLNe0QzyPodjcF5VNc5RH1WLsPDA1v
rzwV7PPrrhuip9RZzxuDhux1pdyvoUB+GIkAwwB7r51LCRXo5Ds1byb91SV0vMqL
WYxweGwm0NMiUGdePNs0wgBQ1XRqXrf5dchohPnHjO93sF/B26tUUyCfv9zEPwC/
5BXk4zog1L0DfmlZ/1eV+jlBQ660yE5XfWwIHTbuuhwFVc17Oys325vmF1LyAE5c
OlDuXNxi3GSERwDXFHn2nV7/V64VBWyMn3jowK86Ez7kK1ZtkhFtYedKXArvkNa9
rDGf8amoVPQF2/8LtIGg/h8y0pLW21Sv6dnnBJOD14v9mwrNN7bw2mF9Z2WHY0GX
Krfk14E2yY7fnRBuIiCUz3knOFu7AoMTuooUMMS/vwbbo67qPlqYsKDHw4n7WFw1
fcw8N+ciZ3FZxFOnXRwKC3wOYaTahyEbeGaYXbXwXnYQkwedGvlXDI68FhKz8XOe
CmyOtpy6WSYp0+yt8gbz4POyljjGXqRcW/XlXp+7c58qczbq81chE9YiKmvAh1qt
de7ft2DNGXqc46KTFVPj8CEH81GwPyxN8DfdU6pgaNsEZcBzThHWvGU0KdbZhON+
WnelgWoZOq5OmY7MoeQzCO8hdkjHc/fbrQrb/EZnkoMt+o721zYpWKxkQdVoUfdx
Sm4mo5iZ4cL0rNnKZGapvqFpTEKRqPnYUu3lDNI5xsztXZWX6psok2dsaaFKgtK6
s5Q1O8dlOKTZ4wEKemhaV8JE6cmMxmJGzuqCQLquhOx4pzSXKR/EknOh30HZuBru
ac+ioeHEBc34cHLa3s0zPNumeLWafZe8UvkyLu2jeULGznmLCsRDzDyEGPBiSsoK
IRoqGoFC+YaFWNU3clQLcC5M32nW2ulHLgqbGir68GNjhV4E2Z73DECEvkvlKJrt
z7wgq26u6ReYG5Rp3qSeM7ffq5LDJtQKJejBtfgRHhGldIK3xBxorixx1Hj6CHeR
tDpJuVVf9OHdmeBoBFMuKw/QPXxQpRzLsAZocEReEWBOb76n8jWlmbG+iUFOIttW
WaKC6ONm2kzADw4iucqhX65u0hJBe06FSUq/tUbnVfEcNkMnguyEH1aGQcxeg9SJ
QdwK6qPzf/I23xjeA45bwrN5RLmCR25JUfzKBIS7JBO9WDH1HrD5t5KiXRoyfXtJ
eaGjgRYfFZtNfH9pJ0C8TIcqHY2lXX9oqh9vQ8wV/gNK0J1SlTEkqSp7S5mK1anZ
O6FTT9FmdcE3KhauaIvabkM3irsYqhKhZfq/X7Kb9O1OHEd2ocofSzn/Ah4Ej6YA
FjjqZQWVZmCmnytvogGkuuXeVLanbOLbiyIiV8wFpc1FapjFbsni3CMnuZrZN0Dh
q0GoFU+K0mR9ufbn3hajHXzwjrBFiBkrOUUoxyN8ZSdX7/0dJ/gLNyRjVaAPvFpx
k8oWGd7Onu1XBt35XavkLDZwKS2HUUmGKE/5pxNTYWxsUzE7EPwSZduuCMb6EcZ0
aZdcVzeBK3SEeyfxW3YNR7FAJa8FYOnDNztoIKxa5iPRWobHs4P23N1IYwnerz6y
AqAZ/vidSEaVVpdt7LNdAyZpIT+tWBCas+KRAj1iKY+V3tz+pNRTXH39Wn5Yvbnx
9yeZjVgcTe4eYvj2Y9qGzaxRvjOI8R/BQDGVsSTq+83CX7Hh0VU3NEb/d34cm1zr
4t1VJHfrZ7BFcVxiN1JCY4xVR81ryf8Vvzy9R+6z9wOJWV46rIbJ+CdhXUmNYMcR
4fw/BHDpt2nUozdgv1NC6ldzL/e4ZNn8zV3nvAbolhyBGdIC8wzzo3aMNztQb8E0
k62QHsSy/koPHl2fZm9c1rNYDMqKpqjPHahWaHCc4DU9gdTAcQ30TT1Y09fX928D
rJp1bR/BC+uvguXo48WdbkLjGz6adhaKfNSdv/F+VCimV2HVZhJqS5p/Rt6rdfxr
Al6fX64XvUJgSag7hI3IeQNCT2X4yrN3xy/x3NPFni1hC/1X8UxbYYFZe72IrrjT
TAcL4n3+HpeV68ERXLZSZNSqtFdF3FWvqu4Cuw0zFFY1Pigy3fLFIeXlEZE5rgAE
x2HtdlS2golFVLOG6jaxRYCkcVxIkHI/ylbid0DILKAlxkm5gLubsW+ysp8mkKO+
wX5WfNzkEYdvF6yzEcBa6iK/Fx2hYOiExnjrJx++psWviAVNuShFrzK+8olDuw0Y
396/dT9Diq6q8Ze+E9fFOmV3WR+wtWOCV1Wk1w0Z1AG9LFtpBvhuc78lGSfI1Q9i
ktm78Zs1oL+YNUr6ngEvUvCx3E2iztDEyoXeztbsHgX5bCkseiI0/XSHx3YENlga
4daCtbJAgeIo6nULmT9gnlfFCzBbIjulp/b2rrws9/fA6hKWR6vmdlQkRsqeogGF
mLzqGrbcGSh480jLmTocMgq4cDGiNt0afU1B6yeDMSelGevZEnLPoH9hcg8QTflX
SpchqWxQqDIAzUmlsxOO6jHxFrjQoyLxvhSzdktp89tOYNh0Ah9ko3PTLV37ypIN
ZP00tHY/uIGdYliNtPsnJ/BwWQpGcxHSAyziHaKmdRmH8pXZ8ZDWpAPC6asEiq0E
DNKdawvJnxwLtmjtbQTHToi+W1Ox5BJSF3gvbHPI/ag7dFL0yu6e6t6taW171mJu
OORkbrVG4jP3kbwPdJvy3UfEQFfFWhXBjpCRkxHStAnEWHorhTwYWTlRf9jk/SZJ
glCKhH/PJRSOi3pZZeXt2RIa5S1GPOJIX5K+vvz0lUxiT4KVdXohYznWg5w/oUZS
88iaXwncs7e2Ue3NZgfunbpwmY22zS2eLXTyPJymsLrzmsl6rbpGsRk/eaBjbZGu
wh85xV/l1QDqp4+hMW0SP3GZADKzMjfFplGm0qcChIshXeug0QeVsgGMejhx8xem
bcjNswbXc/8AKgY/aYGXQMtaS0BHS58OdV8Q8gYPUynbc+guuEI6XIEU78X0krJS
h9fx1IAHm/TB0R86u6nflpqWNEQbBFdCgXo018JLKVAiu2yoRhjz4ID6SFAtePm4
Z6lRSsaIMKiPJkZ+xftGxWNoUFppRqyWMNIQ4cUwdc1gdnd6RDZs0TAUusqqZPLY
4tVXI2DQT8PD1iVLQo+KPpHcghyy9CuxlsVW9DfWBaM93uw5YGilZjS0LFLUyjRO
L60qp8ZuVfO0ORChWDVvSG8OlahA4PqovYjzqW4877m5Ya18SzWvgIwF42mw7qC7
iY/zYiKjL/ueI85fz2mLz6Xw/NxShXyiDBgQuZUNWsJynH4RbHgaeeubtJ854npS
xqqhBO1wcfAoNEWTWl0fRt+mxGqvAvMLzBDWBLH01uOjnT6vB/Zpa/s6FahT7Vdi
RPOesSy2litCO96Nb0cP0zdCfbXkTaPCzZTbbxjKlVJ2VTTNjOTGp/+6sc5X4I/Y
gsk5iUeT7VYJNRl9NI7yCHqt4lE5npFdr0oMNAmaCNP5EkZspvH0a+sPKnE0VXQ+
eBM5vC4SznKqHbGucfIeQ8joMGeQR9tJxdhkDjIujhpW86EjOU3F3u+lHVqKyQW/
nZ/RVSGwiDZGmKBnn0ZTSmQgCKj9bnK7BJOgwSwjl5W1EXi/+7XRzSPvSwapJGMs
8uz2HJqQjGe8N0k8Ap5Doi6Ovf2UX+2F2RF3TcWDaWv5xw/LZE7+Z4Mnjfitog4C
oFURHnJ9r85I/jsgEsp8ILpAsNG1VJ/IDZSU8qFOBv9l8j5fjYoI4j5Be+CKqpIE
S6KQT1sSzTEJoBRo0PNKEAI+Lfv+VS2vvQqmlZkL1qsWjyxgJQ8eJQSYvDLhZf8j
gt2F+kG4lh1yFvuK6pQR/6xw10e6sXMP3gSo1pbZkg2CXjhwrBgxdN58oDncnUeQ
USiYQVD+KE8wqxQUZe9AQGCZ+x5Of7hn3uu4su9XhfDzvWS+PhFeS+vLIgIPyee8
mF+gwsdifTLUEIm+Q+cYig==
`protect END_PROTECTED

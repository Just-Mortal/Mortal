`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OTo5a9B6YCrm5Z5BTWKipkWmtnvMNRsOKhXOMwJXYhbI8kO8yK+GeJf7xVaogSZb
INcNubh1nxKrlA65sWdW4xDUZoG6QNVb0iOYgIMTWeKkxtNxmdSXwpUg0IyK1KHx
Gm1O1pXYjR0ODHGEhyhW94D3Xf0DzGkSsJ+O7XSDBzXS5tin7BS+jkPSukA1Qzvh
4QA/D+/4vulz3f/jHLX18S3fl7inDkoUOpa6phYJIqvB4gi64lw+i+cLy15dxqcd
99Vuq0Mxn5VzjnhFDWGVH1BclVh+OtY+b1dUZAtpKQxXX+Tu8pzxHgWTTNPESMZ1
9vXp2NhYgQxi09jQb5781c6v2lPJL8LfLkd8jwDuVenO0qql2AJVZxSM/BuHYWNF
UDQpR5ljY7vOCoXXCdm5L90ycOnpujgktrLwx4V7wnEdS7LhBNkIfyYKrflK2gwt
KjSgt4gvxq45SOudXBR1KXJpFbRio5Emtbak+g7gSKbgFkL43cVdgMvcGvlfezN9
EQ/ub7PJKf5jiK55AnOUAIEqpfqZfqYMaNYjAgtjm+Aa3kDCgF2/uGCfSRU59/rM
ot3NaBLtLEAVzndBVjWsE0pFB9e6VHy1LnrNGx2LbVTM0y9uuofpEW/yMUHGHWLn
maPlwP73bWh2PGjYfKiiipySQ81/nUEhfRHwLZL2cmLRJniDNoghGuoHovAd8xPC
T37EltFWutWgH9EXmfIO+ESZKCYQNQ//Z5Ulijjx2TBfbfN+9gBKDDmGsGay60O2
PVkkf9tMeL8lpWo9aCHANTXhVllk+dnE4F/BlSKEDewIh/vj1qUd0S0mFecHA7gp
IFB9QP8DK2YYUihQI7DS03Plwrj1cMUbXUcbrIRSD8Kyk9NrI9HHxAlTcPbXaAfR
kSZ/y9+6neHC7Q05wMD16iwtfou+K16f590vaKyTYbg=
`protect END_PROTECTED

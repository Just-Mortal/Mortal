`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XvyC5BHemFOH0mcs5CMy69CMv74XSErav5npxq2ygRV1ZwxloqyFov23374jkBNl
fISxjTHU0c2s59kbKvftdxZSypXc9KpnNltpT9NVYTGy6i4a1X3qzhMjKhCxSNl4
+uYFnjU149jfwWTAe9qkL6ANGYQc7AibRZFsXbo2nmeVkEGqRQIjhHjeuQsbAIl4
mKIRUhhdxXURP695YzTrxgpcLP1/AMkBUirM7dsW+wmfj/wHv5iZDDtbGeEtWi15
MNR+Ec4WAiFuwf2QdE+/ghG9sh3ey7YlsyxwYy9Y26An7dY2jZtp2YkPzQoTAK+x
fFNkyisFuv/Fqd376O6+dnhFCAhq3GPQHmigufm+RBIQiqmL7YZ6wgMWQ6E5ia7L
CDktJjwwsUlMW1zNIbs1dhoqcux6qa0I5xvDrMQSZ+EEOLRSlEHnezKhDowJAW/y
RbkOzneHPSeycrqQNBO71ZE7Ry+rmPUyPvvzm4ffoXLhuVNL2DzGt3PPgVYQK1OM
KADOPQEeOVLZ7B6jVUYLp3BfhPm86XlC+YH8m28YuFHB5nTm7pfa9cMoNukxe3e7
PmO0EkGuQTkVFqJxFccj+odIXEVxhYD+gfLCGd9KPfDfGoXkeiS0DAdsk6HaCrwD
PJ8sSottpp5SMhqIW+kmnjqELSyqhfQUA0/QkZSXEPVNtyTi53JSbIYboozaVEma
ttRdCzZb+ReT4BrojR/R6AI75S5/E+cd6VpzJs/UpiyuY00FKUw+3Hk3w5vRIZ04
y1/N985zd1ZbQHeQCnc/tx3kFqggYi/sM1Et4E968Dv9V+7RjOVElxTDLeM8douN
Cm0pFQgz1V7K2OyDhlRlv1XekWV/pmUQWgRtKAtxGd+Oeax4B+oZGZZ+VMdZy7DM
OxO5v4tkXL0q+CFHUOyiOZzAVP1KkVMsj2oOrpxQMx5l2G9DtyEn8TWww5ol4ztZ
A8ar7Hg37hVDtEzH7XwLxRq1Bia9eXXSf5UHDpml7JP8QLcoYXe+IiF8BBoZ+bFw
pny0fT+A1R6mylp46ioxbjXCnY75RqakUsyJvHqt4mI/nN3YEshPSzesl+SZg4X/
vuQnWL9CkvB/Ut7mNMJxghKNuHK14bT8sp/XXBch59UKgJS+tA+475DThucoCrQX
FI+sydFy62C1ZPJh3H8X0cFZYZsvB8F/qwiJ3vYxquouj0oIevSNOkLK6EBbSj/D
jfJijExL8HWkHG2YugeRpiZwMYZs9KCovuPv31HbGCGYJWcuMVLG8HtFweDpV0XA
FYHkzwA0zc4L3WQYNJ0BRmslBNjqBNB9Wo0sWW9uHP6BwUymt4Dg0mqwjgfzZNXc
bMc+WJ2CHAES8Tqog0tHPjQflnx3pqJ4Sn7+1xenjZjWBs5xyVZqRiwBFlqvKQ/a
7FEWkdTe7h7AcecU5hn3lruCv7UJOa1wO8A1joboHZTMbRX1SXAukMY8Tx8/U1ti
lgcuSA++C34RGTo34wmWKfg9aUXdPHJITrUYZ1Gg1040OIwbrVN8/ISjVOMb0ZXR
U1xgwc1D8q1/eS8hbBEGxoDDpHqAmc6O0/EaaZF0Xo7RFj6Udr0e7Hm+P33nXACb
d0V8KTrCcX47OIeX8pPFYS/LPICFSp3ZOy/pYZOTZzCPvHlYvBU74ZRBi1h5qmsZ
W7A6w7XeEUoeeYOEm2B/vfOrh0lZpBXB9TN5eeYfgeJGtGdeTzN7UvZf8f0A1/G+
IUMwZi0IHMPOAyi8PpORwCjg/D2IU1FzSNN7tK6+En+Q9QDA/NAkqL4cdqrzJDBv
zbichFa2GUd2E4A7NM5RVnQ5UNdQ8WrLfLTPbKl03bAGy5pWRKMoPxrtGyPijBoz
XSnHQxKhCTeqBnmxt/XlIVR5H7/8meJDFfbA+LA6w2DQ2PK+0/vKeYRoq5tPqacJ
AtPsFh+KfmVABjjY5yj3RgT1uQI4+xBAWplXazuaL1KaNerIufibECgtHRCF9EN5
cJ0Nl0OcZRuynp446eLc3UVk5pCvsv38iBxF/FRzi71cVceaKqwX3I07n9u71zsy
HJtv+BDRzO+y91ZhLkdaVf81WPf1tAX8iarhOYy+flAI9ZlYg3gnVJBREYzvP+g8
vHvTMwmEbSFHuT9sFVKb5gkq/Agf03lvEx2PtGrZ6ii9dEh+EZVMdtOVqt5uowk/
U3AjMnf/HTr6QZ+MVhXPxZyL1J7LWiDkR1Zc0vX14kUSnmRGjbkKl9k+4emIDx/Y
THY/W1cP2vdnnYno8PMIuXcUIu4k6JoD8E2eshv/bGuAYVFcBDvfZgYQcFZf9PZ8
dalTmxQu6YBEzBVtkLeCPa9QwJMrR9X4DyS6gGkBmpE8kGCdx8PFihH+ulHHy7sG
xkkItg7NcD0JIty1ZGjmkLmZfLKjbPrxmHi4AjqoOoTUZuWgqMDIqkMxzACe760q
LTV21h1jb+wkdM2uJRaQy5Bnuij2/XR04zbkP1G4dS+h3iKTDzd+gRrmBMX0PxhE
FOopfxjC8R4VNngLN0qrvjUn3mSvdv9rV5No9gT/BsJWy4tuU/HCPlmOZfUDqrXa
9fyPCLzg4bdUc2XVD9jOh9VbMciokTYHerddIwC+7p+/jvqVmcaCBHH/5sEPvhuC
DzV16aAgcnXiy6N6P2snR/WwsF3v11F1U0haxNAqFVVwb0FUEGsKdFKPOuSI5pUV
2fYKiuZ/6k2TkwUqDYuBguQlaQWnw2ikIsLIQxaWxDLyhSHKUAIc8CEV8rXXo22H
NNTZN8uPCrlVP3IC/SKCv42m0kKxJYjNPMo7DxVlz87qEWSAmx/xKrN9QjvfzdaX
Y82hm7lfRO/Q5C/Fscn0624b01srwQLUhwcIUSB3+PHIF7k8qU3IP8U79b5InvXO
NSTd3KSvBtA4ct5B+GMPQhJtAvFKVaYb/BNBTKiTNiWzuEu7BIL6q5svNJG1AekG
35aX3khpYA9H6whDPAH3rl+3udmuSGIOMkikezEo2IP2GC38GtZr2WabLCzBzbX2
ac8NN5Uy7+8ALlG/wwf07WfHVi24vdoKlJZgd5fT5fhZkO+j/yoHU/ULa8dZgV6P
a4ehViTF/IMQomDtViJ3qJLX8WwgZKvo04nNtTuFWkCe3nsbbMRZHu9B/tvh8nli
XONc+x7R6XNsd7pzG/ALv3mnlHRJtEbgE2Wu8GxVx/aKu6/kpQjHDCxG1ye35Ajz
msWedHCA7bsqZs3i4Q/clmpf52jYHuYYWjadHySqlU7pJk5plKRw+HQsq7EDsLV+
QHDbuNOMt0F8AnFtmXFt1uZoIHFxv7U4ZIfqHphMvFi7+9T/FszQCQiFeAMwywTk
9scIc4UaNtwChcbKGqjqp2adqlDnxZnY2ATScJhI9V4oVI1/TtAs8ZMkspgAYHNj
oQzIbc1FBLBHRTfmjR3gSQgUchJ0e+rqdzV2+g33m+9GctYdRpPzGkJbcwzHXX6e
jddg4gTFYhPn8zryFbqMgf3LnVStoUbvYPIYnAP1TsujqcGYGfxQgVeWaN/pGbrc
1XbHK1reIONJW2aDS9ZQvrDau3HMo6+n/7dyQd+jFHMYsvWbk3Ezh9KSiUZ18X/m
mMI2i/jCp3FGFU7VRiRICO1HBovafEfx0iX7jc/EQzgr0e0x5vnQuVS/NhTxtd3f
5rKHxzBNndfpiq35+K2vV30iL+myheZCEqBr8y7YvCudfi+RCQrEaekUaboJOIMx
oF7yHuUsht8gEylI3fO5Qza1Yd9doFYTie5PMR4T1NaqhF+4NBeJxz8/7KYLCU6x
vUk3TsZIPx2jOstYY3WAgEQE0cf7RIQfkettE8gd1vFwkpTv1B31gc5lfvMq/20b
URDBVxJShd/nc5p0bfcXhonSt+SNBJEprRJzNj3FNnCehdaJIHOREHpBEMO4rz9X
iUfQBmcriGSbxwOrz49kqTy0tMc5qfGdCwxURsvbOANvbs5EVyforc7whl7J7zW6
//joMK1rN1mdI9KTXVjUP8QL7tdsMEAbKYerfNf1yAQ=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qcaSMXan679xP/GXJiEWAFVjWB9K6h0au6klnnEom+Qzh688R/4FfA5wXZH9/trV
3GEkwiLtZj24pOovkklwUxT1nnDVdTZ1AMTjo2hJcdaUs9GvpfWMDb05cJRhqMdu
U8OCR4RjX23Hq8MzoLdbP4yD9Pz3LcfQiDQHOghf4o1oSHQi4V5lIMrFYP87Huap
MYzDLD3Tf72Yp9tGySqq94LM2+3TTP61a9jJlwdLazW+NxatfFaLWxPkmF57iL6r
zXD0ysHH7plGcmfGRXUrU2VfRTLEyuTHuAr67uODDhgzr0+wMcL7yhAJHNzYQ9pW
J9IpHm8UmY4bPtDfqyqsLo8gf0jQ0B43UXQqfvoZXUKL/itJexWmyEW+bv94nGmF
0Ndlq6WVX65RmVEEJoSJiytAi4M6G1Khs7S2ap+Jb7AFyq6biusXh7vgQ5xUrh8x
0/oBTirxdhT8rQd2YUHI8iwx7s8P3MTDBzNiUgf8NPvpNaGAExEaOf3zXUdnnpnU
FVQa4/9ZQYD02O6APL44iyy4gYroObRfH5FDsRvsdEq6sr3MgY0rTr/XUv9O/8nc
/06mj6WbsUlHWw4AxqPRlycvyeqnwXp6E71jRdjl3cqYa6rx60AuCrt8Pv66vST8
cpedvIJns4YwLeIA9a+/S+yGzM5naoxdeZbyVByxlnFg9rPf8KaPYaY9/OFu9fKT
pM2m6k82GT8oRvM1f6BvIY97UrxjpsbYGXWqDyYVxzigvTVn3sjcBtj5cCjcu3HQ
ZQ0HESL+4ywB28XMOPU2u5iYK0n/fYeILTvdJei6584BEF3U2wCNC2GB0pvSgX6X
AgXrUPUH2a6YOzljt9xE2hwjQ6HWoXxXQJ4wX1el3JnghWpaJ+w7erVmA7fOGxtY
/jw4lKcQnBLOw7uBdjfzMiYpSVHxKCWPhkyruSZpJeGhSzACxbmbM/Wl9X0Y/s3U
NJmuQRuCDd2Uj0yOoc2suVJQgzFux/TmFpQ/3LqQA6yoh38OwfkbYvQ2SyDFmLd8
KuH9w5NACPwtmcPaATDWWbcA2MCc6kAw8z7CtVH+b9GZz5wXOhPs16OQQ9gDhw6m
4cbFrx7rRwIR4m9lGpp26ORektJMUUBhD0SmL5mJFDiYdKeq0ojvMH9q95hPOthG
+04d3n+N4riku/ekCFf0zQ==
`protect END_PROTECTED

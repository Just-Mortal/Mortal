`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QR2B05DbE+mlqRnPpSvmW7SJlQ37xIaAV0US7VgY9N1fEY+If6sZpbetCx6ktJsy
RelTKZefIvpwG2oSKYy5wibQmSSldK8uLd1OPpjSHCtQC2UGAB2hT4prarvBNSfv
ms8xH4/8PFOgyuW++ly+J7/Q44KbXAVj6lMDkN8W++/xqYb1l1may7ddx5CtBQtT
MDz+kzRhHpRdlUUTKEI+hXMn4sD0pW0rKMzPi4txLnhrlamiLa3eqYGCci4kjUEY
Q01jtJc+Y/2iSKCT6FtHaiIzPGc6bd4P5FI8ce8a0PBcBruz947g+/juMCZvkTN0
BZMF+W7IK5RGBAJziru69FvZPRyVE0R7gacdkiJM0P+3y7PXNgXIpvcygYcPET61
59DcbsysX8dpAMhUzC4aQuoIZ55g+L7TMOmOySLQFbLLvcfcc28USWorO6lHyteQ
E0pFgl/yDsODciNpLxhmd+w7/4Qa5msMme0wMKmT9+QpVP103RoNAvIcJQUy8rzj
YbHnTjq3Rh1sOlu97dVzaeS9VEsjA+aU3jQ8G/9hN9uTgytouLKvRMC1nU2KC9Vb
a1BNNO3BSXyeG+AGhXwn5Yo//wYPUF2VekRpwcfkPH8D2PzqisMYEk+1ybFkMpy7
zlh5DLCugv0f/wWCmJsVmS1J5NkqxW9Ev+ysGCRyWb0Wcn/9sSRD6oSJVTjEM7EO
s5XSQZq8m7GaiMe971belCN1G9Na+b7RZRAwON1yJxEPe1ExjRcEJNtSjLBBM7ea
CeCVdwS2ofsILOk26tjZVWKPqBhUZbQQlLL4hfWxQIvm9ICAb7IlRygfMnLqJNqM
ZQDX/SoNwSAjkQDoxHdXiSPWwzUlzNhXoSrFR3JOcCJ3zrIXXhbWe4+Xk1PLxkye
6CfGg3kmWFgP7H7qOIZEGbnFlOlMay5BQqjNEAoMRq8ehOzPHeyKhn0b7GSYvpQH
Zwj33vOXHAncBXg1j4I7IinGCL2w7ByN6Ekkcvf75wFhFLYPGmigTAKSQzg6iB93
2aTfxTx5UDQmf2Tu/FFAi1dbiucbK+gE4UKuMKAgHefN1+fJ4UV+ckudIHGH8mh7
yx5hPoQhXAvwIl35Tvm4m9sq48wZNunpHgG7d14b85BHKlZQL+7scHzV5Us5f2zf
XzTml76oRGhvDZUwfJMC/5GhzaOsSojQBjmkTcRc8wQaTh0o5th0yxvz7OYVq/WC
pw5NK8WD4h/iDgou3J/j00kq6ROuk1t61iR2q8OOZcYVaYBtE8UuksTTJhKHgGD9
DTtKGTZmyuZHJL13T8WvZVhPHxmCTVjvf8y1YHH+zylzkw+xo0B1aInwIGm/K5m3
xoVW2GQx91rDRkis9mrC7cgNQZlkdVa4fiihCY2YMkw=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKixv642yMHCz7j5npo8jCwIiz5tHT0gl8IVmoD9Z8DE3CIJflqxMjh5jJ57i4uT
d7VJjFnHGsdpLbdjSKn2ctlqGChtDgOaNFKYbx6ht5ZDtGwU4jgJ0gHTDL3lvCwK
DiXtijqzuhvlyxuNQTOFsef2gOq2VqgPDEewVps5PC+yO5nBoTpvWIsZnZkmRvNb
4QLBUezGzOBp2a/qdTvDaK6hJdhbZWDDmPrSTRu5ub52O5BUkRqg8UAwqFrxVh9s
liBzaHFrhlpWD0HgKk1E7pl1WzrclbNFm8zYmMeuRF78kM324BsOmkQKdbBbFimo
CdrNgucBe7e75JTtbOx7bW6Uom19Nnk/C5qg0wkWeGCBYxfQWkYVQCoyCtvgHJhZ
2jwvtMUuWNYXnaa+d7tQX9cst8hgbiWu1Is9HE98OlAan5FbkMQupRkowebbmk9l
k4I7Rj1cPANPsAEZku1I6PiYLuZQmPMkoBORMWIzosIGztA2JTGEaWi4lAf2NEVi
uAlMoQOd8hWatJCRkI1Jo2cJKElWmnKG0s4kaOeR/vwjykpDVrPurWqaWdedY5T6
QSqdGs1wBJ6PB0RD5PoYLRfzafnqEraK4b7z1ztxgrToZaRRdA77gjtC7U/9MQma
ywK4RlQU2R5f+mR2E+pR/M9XY9aNwzdtnyUPBAXulRwVlc7rM3IKjS8h88sG4C0x
7ULCPZExam6gna/C+YlCpdtxiZlPCoNryhaDYwgbEdl+YEDY69wsJGfEQu8cg/5/
9IJ6zHapBivV805C3WBkKeYUxDfxinj13p+DBWDslfrvyR2qhoFZW0sOTJ6JivJ6
vCT/YqtG80Jg38LxvbSGksrFz+M7Ed4yUEvostjHcU6d3Ix72mlMb6fX7EgUbJJb
Pb3L7Px95GZDAX8cPRsZyB/VHQgLVOVN/2k0p7TgHDCn5FibU68AWrwxmzsmHjso
ymF6gSDM2B6/WCPOzoFUstKYKWAt9Oc0y3QEcTs4WRVBlA9ovQvFvrQ8bRsSfcNA
LoSuwpFYDIj/8ZZfyyyqB3q6AEY+utm61mFp2fdjSuwyyaowK+47fRqC3jHIzaC1
8cYDRsk9JDPV3W1KCW513c2dDcS8cDGGjqfEW3bEQzUPzaOeyAwvRaxG3CVeU9P5
DTyRXPf5YxJPKQNqrfsBszeO0ypt4mjoSJoeXn6zeQgsCt96Aaz/PGfLvbmAH3o7
l2WSpKr2q9uOcqlEoj7arnf1EAOQ5HFOCvV8xUejmmwfusKPp3rMsQyMNGpxap9P
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVKSqGio8dZ80ze3vC9lmUlYC/e+CLX/nE4/8vh5g1WQv0JewLAeXVAb0VeCJX/t
xyixoHyp5TniAmE5lLHFqA5OAjQhzbJxrsLpZgpwGTlP5p2Z/vBBfLxAaYzR6Bzt
nXi0Ip9MB9fj6z+oiYXcHr9VOaqIILhFsLt6gZcT+BYLhURDnQjonZVN4D9NYV3H
RpfTD/7wnxHQAXS3LUzk5/tkSWfuE3aebX9qjfoVaRfbafj4PaLm2RxmiPlzJj6I
IOVnQCXgY3HxCRlsquvypxfzdsQUXA7ebgMpBmep3mN00fJ0filwuNjPWN+elWmX
Re6htoy8mXplUWoxcZVNPQu0Gyw7s4DcNsulWtF8xvvmitU1A/rwVcqJj+UpR7ZI
LRB+oeDVEdShM9afwS+W18TFadswhjfg8rTleCo6gwmPBx3UbqFZsBkfkSu8Nz9x
+WaYsQ3TU1pxFBjwKbaabRlDr78NfDtBEQLdDzV1+ZqKODbEqYkusLZqHrg9a/fI
EMFUTC1/sypDXwutMepkFKmt7ZzLLc4GqF270tuidI3t5FNpgRcZus67rgMtnw3k
TvuW846f0LdDtpxMKdYq3DkKVbLr4pqx6xja1yQEcjDcg+qdkiGMwWNi/+mU3JNw
CdamEDTW8HTKC810NpIvX+SOVtAJeu8Eu8pjWe0MzGJJ2po9szGO76JDPKL8OzqC
Q5A0XuLwCTL2K/4E8YgGsbqiPaZmN79fb6LaCpkKiN/33mFUdXrPkQLf6pj4eTSE
iQAwb2AYxbuvep34jSm5kjmZDOERU4Hu/Gsg5cxCANq1AbIc+fLDNha9NdLHskgv
5ZI693n7wse/z89BKhveS2fYi13eX2wGUQWuqukkXXilLGOq6WT8kNNF/aYlF3Qw
XnP+fJt7gSQ/NhiebCSVRxwSHayNVi+uggvXUqQY2f2DVH9QCPSyCct2/XLVnrbV
7bSmS1K8yfCVkqokKbu+LsK0/FQlnNznfWxuKDoSVB9vpxXfHMWTgG78pYHwSrY3
AIzA6DJFmgx5DWCIdCNwhYy+2Lt3EUwBoEGEaP4vOEQuDssk4qQN6UIq6eDQs/eh
BLvHCkM/HmQ9nB31pE2vy26N02xnWIQosdmgVhi/5ApuBNTtAk113HPfUILPquHo
7KUpu7vKmxWXxX5H9Qv43c3xfW9tFt3A5PoMnhvHWSOOtqxICjPTmJy7HvwNLsHG
0v9ROUn35spaoBrSdd58fPxMaFKx1CuKhov9cp4VVN9zTh8IN4/eqxLwhZc7VnKD
DeFyjHuOAm2z7DHR23PNGCrNp0lzhKWo0IUoBrId2AgBvhcpjc8qzPlhfpeRkbqf
FAz0+3+e60WTaVT+u+xpKlkLXN0KXqF4MhU3AOpGfVuzulCl6nfICFYP04saCGCa
Y9pnCFedmjDVMzB8Xmn8TfUb3LdNxpSbtsBo4X6QwSJuLQekRAcwTmznl//8xDTZ
o2s6I1yolLKU8m7SQrmwi6BtJ05pfSJVcqoOAX2cBA/plsnISZ3FBJdfkS3Sig1U
vNmALTwOsCtT16C2wQjJlEbN7QaRk/Vge2U3HsSz+X6jNcRwt1BIJa2HHusXiwOD
BnVcEqiGNNWmDvMcNqyb67DKHOiSIS/pD4SzwHoMu2IhFDupp3Ufbp2UJfhAu0pZ
TWf2bit1VmkDhZ/sguHiDtv27CHfm+r2HYnIdx8UCFH3Jm5i1vzhfE9bVQRXB8Tj
5/rFoM8YQgBXt8OF0kJ/VktQ+SCYe8E1ih90782QDb70PlHsdk/qwvvV9VVrtZNC
ElPR0OJVn+NIeuYJsK29/aYEP2HXljsovqVH9F7dBgZsDZ7E9PJF3E2MyjAJbiOQ
tbLomcOCvTdMXjGFFAuY+JiO3f492mdawjMyQfz+QS9GU+ehIZCIPzerDbv6mTzf
1jGYL4prNG/rHQBTK9v9H6YS/Qu2yrLpPXvnG7GJdJtCLya4rVGQ5mubsHgaAkX1
4LrXg2aF52FXeeKb7sy2ixVxU7QKDk7KbYlVcd72LNa3gTtc865aQsxRdXGXv8Wl
qrp9sRxh0U0SAKCr5MqKLF0aH2own7DS4Ab3Hl/uQJsudM5bdpIADSs7egaZuZsr
Ru6P8XbX8kRMtGl37BIMmzMDRJ8R3ErbQsd2aHFUF35xmA1FXN8SkGt44QsRsjZ8
sYugA+5Nr24WvUvagxlUjoa0nHjHzE9AE5grqvc76FN0Pu/c1hoY2FtFAahiHj8a
rUw0zrrpUJqg4fhkAQZLKsdXwjc0aNddyV5oo7odOjFgbgnyu8u+/sqnSC2LuZ4e
UmiZDcGdWrPiojVnqpNQ33HVxJy610TyRWwsp762pbL3W74Z8i0oJVOftnt2jKtv
mPHmPZ4cNIslA0yL3x9SK+FJy+8GSXTuY5QqVbvz6FZqh9JGFeOyD6ddW+28uWRW
ecvyrMCv/hgbKa80A2bLKjFYrfpidLUX35nLW4xGjNsKFSDe7yqUpEZeolO/imsR
ur86C07+fCTx/mdZ5dNbqa+H2B4tXMytBA9x/veVYQGLOOqgMK70745rfVlKbAxR
R6hBdo6vXqVsxI0COhsT9WEOqrMp3dx0HDP1HDMR+MGTXXVoENNqgNjgGnXbxT5R
J6LApFPAqs/7hvddHFaOODhJWKhi3P6T5EkVDborKGfY+uVkPeEamEv/BnaqgsAs
URUme0BOXdzmCOC45gN7rA1r4tmuYfygdw2tBUOFwIgbRRy7fm3iAif2iiCQF4Mp
UWRHIIEpo85HvcQw5go58Z9cisB5GyZrvMKDai94U70MUkvbUI1rv9dC5iqovqhG
2tAUqQ+6gmIyjp+ckwVbGU6NT0RDQFur6ECiA2Zlefpju7C2SxBH6XafXDnHEsTK
mIdb8c57xD6lSgMD6Nrfrf9n1Q8w4oLUOB6xxtUJwJzs7DlT8Q7WubZyCjqcl6a6
xWwl0CKMTt/pSzM/WR0BlMjYUmg9GThYUPeV8z4O1gMDHHplyl/AgpBzkTtYNX7I
eT3HwNpXJ3pF/jCarjIxuaQ77hru0hcv9ulvFldtxGtZwZ++sxslCTIYGNlA6xUN
xFbUg65mGkv3ely0wwCN0PzaKNLRe159ESCjNguirKWufCTOhLKVF1jDPy8RFLaj
uOF5G7Cj99X6tG9hu7V78J/UC51kXM0rm33xkZfE8qksFJ6Wm+uY3X6vD8+gDVPd
AlOy10y31ZQq/7X3c53SQe8b9NoyD8PL55gPdNBXRD5kE3A+dbHT1CczJwwHcYHb
DwRY9zpnRrBRLc3QiutbyP2fa7VguiVoNDu66ICMHRf8E5S8eyODlKSZSlOoJ8Ot
s3OLGtUfviaOOQ65OYpzQ6fQBI1+tKnh5+2n6yzp9MWyivEP9cuyjy9g8Bq8CxbW
xJfJ7HTXSz8KiHZgr2K5OgyGhSWf18bTey664jCT1Zbtscj6N6mN5AI1NQNbH0sa
x+vlCNrPlqOyFviWR00+sGJKwHTPTiW3TPaB8V3nn4m4pCLLUhCvbUlBFOuMJr3f
vs3FZKvD1IPtTVE6Wvksrxz0RQMY7gL40P1NIo0w/QRmCSSp/wOqUVbeiiMRFQHP
KlKMFtQbkN28Am9cfWr/reOEmyFTtZmohPXEcuVqCHg=
`protect END_PROTECTED

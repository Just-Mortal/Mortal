`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g0NceMG6fQriXDjk1ufBl5Bjyryg1BWeWkjibpYPOLSciNncyC3ewOog/TGL6ULw
FybW+fyxP8jNqOor282dr5kzsNtpwtuPzUDQRNSFcyma1/tXyApt/3nfxUoLwGfG
ussdW+/KBnd1dpShg8Ef4qqk7DA46yg/uwkcqcQNgaHjCXNr4vmUw2N9hRCn6pxk
YUTOxadFwhRwnv/2xj2Xn2+jGmD2hjNSF99PvvO5vkMO6BX3MPP4U2EPuNrT4myX
W7yKbIzjga5D2FNOkaZFwtWy49jZ1J7bsasExrJj7Mg8CWBIslmTwf9LBjy9Ny3u
m0iHeP88Dw8RhR+CrLqyo3RgfzQQj/ZcLov6nmllI/mCEGUCl33UNFMDO2TS9D2p
Ncks1UMuxKwtr0zcxhW7YbKU5MMSQ7tTnMwk+6K2XEhRPb2Ok2BnrOaMwbTKJUR+
0tbbVOATfzSUv7ds0Q1HWb9q26V8JQcJ66lhbBPZgTGDjwdP9emu+f7MscOUBbX8
vQnsf8pYsnqXP4IcevC2a1vzGEkuaHNx5dCK7jWjdZoJ+e4IvvB+z4zokTOFpk+v
VokA4Bo99PvBPnJWz+KmNSpZSD8YYJY3529bQZWik4ykS/9m+7MAyJAq3wJTBwy7
Xy9bDDCQXdsYHbGBnEShDA00iXi/5dmg+S63qL+L67wiB7UeSL3HZotYN5uJaUCO
ZWM2TT2kHd9V9BqJROePMagtKaAsgr9xrUkJ01Jye8TbWNiEHRLJXgOZ1317g5o1
0oVCbQzcR2MC3jDWtm88/A==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y1RkydopY8I82ihAUrr816eJamf8beNlB5hDoNPnMFED7BRysBOrWG8JGC1SG4K7
PdjzFHAuN/mW0ZDp6047vKb02ONbF1/qmXGuDEFIXKkBOSNjwK8i8yKYORLR34pV
tElxhsJmASRCCCo47z/Jfk/dEPIkdQcc77ybNyY/C+QkJO/j1fcXn7H8U1mDCK6r
kXXTqX1oPPmaAdxupz1XFFA0T7wvZWYDuBR65KwSKO2Cx50LH6FPHXPZqDYYI7v/
wTlrZvehVsE+FGZaUGTkweV8KDX2bpiqFS3+MDzeKwB2LEUhYdyuviVaSBCGtKBs
Cu0znFJbIDF10DbzII0+bzg3o+8LiHLWuvs0pM+re2SkfgcawlyjxN+IZTgJb6cn
9ZHrQU8e6wKWb8lzJHJNj6GDbfYR/jZBwQBlaOGsxBg=
`protect END_PROTECTED

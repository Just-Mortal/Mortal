`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FyxfKBMZFXFSMEvITdzIIZVVRtb0z/rtif29XZUWT68tIbtmFdhzF6OHADcjvoR2
1xa16OKRMJSzvdYqQUNQ86gp4TRkTUuwNJKv8X3wB1ys5niatWmOpv57D8ki/HoL
dm3/IpVH8fx1ZnJzKtFSqs+lh1d9JeSkEbNX7AceO/MxztyCt2KR6uiPpHbuip2A
`protect END_PROTECTED

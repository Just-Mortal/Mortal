`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6I8VNsqL9pgpnAlTv8RByTOpLKnulYw9goKAb+E7gGNlc7LukGNQ68CfUJYmjpCq
i00ZNBeQFgu/rgPO1mz+pXMD267sfHBNNBihc/zYmXG9wiNAE/W4PHtyZftdDgwG
yrRX8R1AhLRbl1NzjYE2/wXByKJXJetnIOalkjVHmgkZuwkSt6AWDHa0yYnWyv+b
EJd0ZicpVHjJDAu/V+32SVohNrnznZ+jLt99SBslu85a5mlevqUp7W9qrwSAp/19
heXOT9YQHRjpufPwjaH1PvUKNvEZdnELfCNMVE99hEn/mHQn7Q6xG3hFvUqTx+8Y
EvCMoEJZkf5yZhDOCEY1NuODxbpZ00mwLRZdLTlC29Ughs/zuBToAuQwAW9kQ/dZ
eNhra5kTytQKsXbVbyVmi3Q1TUIN48SGs8bQaGQT31D2YqMCahUvLHRbrG1/S5dN
ywBz2jDHS/7jBERXxGlnf5fW6GOE6ylE3E8isRABKrBHmsv2JiDHyS2aDxilHoIn
XIZO4bHzgXHsooF+9/hmRt6mh+4jxGcMm4Y1p8z1aVFeva1aidCzbxJ/xcsEq/6J
7rizQZ5O9nyIzsPlqXITmS4tY1BTDXJnqMaDBMat5ShJ7BzMQLcETAjGycqM9SOn
coWuCJtep4WdXtuBwpyrTnNn5exQqJ8FBGSofcweR2ZC4hMt0D/yVrbu0ggdv+OR
dSoM7akOyPcq1lwziamu27oDH+47ohdOJCqycT5+9jdZEvdLa0BXClnnOWIpYTpt
pvdQR/JEr13/d5p/QVTei6+2Qsj2LzCK6kFoxVXY5PcclZ8VGThAtnozrxv03Pj9
DDJP7pKpH+YRH1uMqr9ot0gnu3CdFyNV9wd5gxiE+ixfyjyc2U+5jHk9NQdTVKmN
tk/xNvRutdRub0A8SS15zR09iYoVVNqJSZn0lWpueK3UxwqHXOng/BM1NOFS50wo
wdGA5QIyevvTKzwZOykhdX62jQhfjCWO2LA1m4VzbYkloxzVpzxSRDlHFUk/ZL97
mHUsyNNVWdYwTOXmOwXl67jczXpEmpOxaaTqEvnncJZG+nnSaa7aOycPRu0KF7vh
yaDLOg3S++pZTwLyTAQVzsNr1t4laDVHTWyKdXpwdIs5PgscVsBwOR1FCBps1IVW
wYPea2P27LtrZnn3uZOpq7TOGHBxYeuLt/uK180auAWmTIic/8eOw2dX+xptPVmn
RPGyfzSiZCFynMZQ6DqPBw7CVkyZrwU510cmtQeZ9wNFvvqEtv8t2qI+/fitRiyb
sKYoLhi1cIU1HyIrJ7JRG98jJaNQFJHhLtpfr7L3v/J3xRfZmr/twAoT67DUBzry
FhuRcA7Qd0AacJIpZGnXShcFxRf5nTtfS5hOFX+BUNCXHZdt7knSK4qPVL4yxkYn
+JLAEWUz3cPbFtcM88Un0QwPnUEXUAk6sI9mYL75qO7wrqhsLujZp9VBGFW/iYVJ
fyo+USFaQuoRQiyVLVUdTUgpPYIhm8FfFwDU1lQOBsaBQCBAG7aRVdXpOTTr098a
Ihl8xC+zt/C5xPzW2pTd41aF5Pssh+uwN4I/j08/5cp4xPFNUPcpGsvYE9RVbGm/
4Cao/PNGBv5KS+yjF6LdQZbTP2Fq2RDyeYuM0K5nP3RFsdB0XjI1uJKCnMo9Xlhl
NscwbRZiv5gEdKkM8BLmpHKiMUgE+co8ZzJskfygVJ+EBsh3BLDCscnPsrW0WMpo
Xnm+SjYtjIQe0cW9mRZ8e6iWo/uw6FspHZlTXNTxIZ+0u7jPoztDlzBimdyW7/X/
6IE92cL6G9MyjptAL3huBnpbAlEDz7LNzC4PYido2yyfckoARpAoxsvac7z0h4Er
rVEjMpIHIRMhbrZtvIr2tuHPZgsAgVJVR85KM7MYYLkN1blXrK7o3j3avpajcFzU
/DIi/9EaJwv8EfSGGbIA8u/XSOZAH1w7at4oaORrI+almpkPHtaJrr6Qg0/SYmNE
bIaFXqyiykpmRY+ZnHqJyiRIJ2S5r1weC+OwyYa9EEciuqmbjYgSLdBA/GlH3aqX
7vDlPQW66KT0l7MDm9l6ZGvvFUlpPZ8xgmmuRgNFaWIqGCn2/8R6X2WD3bsmCp3a
qsO4il+NA1mA3bRik88H8cm5bk9kxIEP7n1tSM4ktboMAkfdZCxnNeRO7jCwPeWb
awP1BcuTFRKzTyewFrJEeKHI16fc0aph9tJnmwG1QeaHU69JmqjxGwVO1FzrjetV
BvVvsBm64f7PogLuY8V1nM9SqHyounMH1p4iA/d30trx3aFx7m31O4p9maW8UEvP
K2OvBqLfUBVWAPqGXfsZUzWQowujeFEALmKZ7wVmKPd75j0VIjYvotkqC6U2uwpi
`protect END_PROTECTED

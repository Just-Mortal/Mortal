`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wLLFuu56+D/FwZXcyJLPZ6boOwTo3xxW/mZZi0IXfhAMhjxDFHe0rCGB6aC3a7PL
SGBnUnBak9w75lqesOcakq+UUiSO2MzCPNqFOrkLJOEdb099Q3u6uvTI7qBkpQ4x
p3/oX66EwIKN07wK/V4zzH0cjVescIBuaxIteMpsXImMriVDXOCRvmUzhB8ZPOmP
7JY8vmI3cC3OR8siraaWLhEACswBOmwIsWGUDrPWHUyxcB2pkKjtAnYFV8iEm8+V
RMqot9PCcmff1Iin6SYCb810MyKYK6f3f/hgs6O78RrwwRhgvJs68A8KKTCXAJx4
6u9Jb8h3UH/dHEJUnE1QHwLRDRJVFnHCHTTmCiWtD0GZQO1gd+VUO4p/KCURZn2z
tBnOdv+bYPJkTcKhJpo9VVfuvWxYO7QT+aNINQp18gJ+e8UV88NvVLzSomEjkSZM
bl59io45AYbo8Fe22KNZ/paLMNfvF3CdwawmwgG+hp24e7fAXktyEPFPaV2fv85X
uMCr5Ou7rjiROwPAV0QcWHSLvjUGCBBi+Ey69VmGmoo1Qc/OSjljXo9XXpCvbR4W
/0or4ZrMrg0JERPsvxGNsB4iCU6OCPHIegFmKPMm2cRbeOBLdzqyQEXM5B5IjjkJ
kAyJronMaQEFlHO/+nBPiI4iuMxJBkQRUIUTXc2QZhPGI39pnv8Weop6tD6W22XM
yFuno8d9sSV2bHK+BdhTk5rBfz0glZ7tBQkXuqgx5cBGm2IUnN0WPYYzxPZRQwNw
DSG51QQc+SKU7wxAUffvkces33Oo9CKqWPtcm1X6A7N/wjuvs9IGSqjp2jajg1Vc
DgvDXh1fKU0GDvrGWAcurNZkqZ3JQ5ib9eTHsdL0UCpC9cCQp61/1nJO/EPqFcBS
Jr4pITwL9i6haC6snhKpbTQ5LcefzukMSYzJkxowFu8v/0GNz4B5h/oEi1HRdsyK
+VVdomWVAYfNwrIF2V36KHMRO0PSKIAtorenc2RbKCkIn9yLq9IA7YC5k/kBaY5+
lgE/QwQUrewoJb4ng1nbynPa+rniMV7CKWK517ZAGX6l1kaCHd+cgDhPkr2j8rdA
qdvadsdoM6gQhtcjFzyPKWmCGVM+aqmNaFcdsyRV8TENC69FWyyX/A6HTMOsige5
Sz/5uKeQjfFBBvvtHQiCf5fIq2/6nPDhITq5m62pWUIyllyfNB6TO2SNB8lkCtq1
tkT8vssz9KVp4+WPnEmu1IDLu1aid+BjO7fXshB+JKLewuD38OlERFAqNDLSh8A4
4Eh3s2I3vdKbLUSV4AlQOVishuBOqSIca2TAcy8KJrr/czGNuGTh8IFeFQCXxHao
r66l/pgKtqxcJoNweWvYCwjdrAx/q0hMocLY3oIzozAcM7y3sRdMIUblNzsmb2UW
8igjNLsIkaXlABAwaiHwx15ZA13c2prmJyQwjRrS/mqccut+4S86qHulCo5+Bkdn
3qjxyVlAXR2LHnN1eEMC9YAwhz11eJ0nyMqb/G8SGU5LaiMCLdX/78wzr+MVRyhm
dieKIdk7baO6DGyA1EYaKvybfaEX+WgtfIL1WajBwiebfw82FxofdZQeVan15iby
fJMNkDMdBNJ4A+lff2fgducyLiqSUosfAFgq+oi03mS2H2NaQfH+tRcYlaCuyQA2
XbyJGP0cP/Y/bwvm5ZPoD/aixrNsWNwlRs9CEWplxMbO8gS6AzhdvwSITZMgkjhL
XZC7hdz3BgFKOkZervBXbukrZoaz0hEFnUhaRhdxaoOw7hyq7fWyKw8CRdrtlq7S
krRE2p3HTE+pvSWfLzH7ZiG/iOwMTW3o22K+1HcWzfjJSZckzu3gjpgghNpZ/JBg
cTOE7IKtYT8VrTrQqVZsN+Pb1hyz2ewe5uu0QBFIgkgEzoWzWdRdt0UTnGcVgB4W
dsXEdPpL99ps0gbYCgRS98w2BI7hRaHA50tuKInMepn2C4fbQWug8cUBfVge1nVG
A/SgX1t8xOPLPofiWG4eRwlnvJA/DIVcSR2d3jS8aJ2hXpP6tR57Qmd8iu/asMpA
WIakYPcHCYpl91PYgEwJRb10hcFQAIYG0Iy/lRsrBc56nsvZUlF2Ya4tcZa/dcCK
VfrbvR9QUbym17j3pHYwQz/jQ1lR7zwhgRWTDRszo5gODRyeO8+fg6wh1XoqwJcD
CjCxo+iCYZThfgpRqWr+RvYCsioSDzKdWkgaqwETc7yvVjGUGUUwodU2L/ihG3cS
QaSZP1hzVHeuBPS6CGqC+oSUhY1Y1a1NXOKHZJPNl//4HHec6HThuZkko5OmcZqY
ImUsaYZTNWvxh+K2uVIaGNhFZ8JKBm8yTDAo3RNfvHwLdnQfRrz80oggJaNq7+ml
yKNKL/zAQQFngG0b2j2cMdGdLbw0ofyspXY6jxE+GmsWANIsPQus0Z1gaW9tQMnt
GdivWoLP6sVHkuBIPtGV21d5mCdIPRhpdt/9Lost8XwL0J4KSnEaGabJWJ83763s
WCTGAG2bAB5gXN1aRDxAk0GtoR6lofY4U1SZOOi1OqVX0pM/PiIMDBYSDUolaEQr
6d5NsojA0qeRSRW3BqfVSLLnwyjCSPnygpR8t1uqHjOZzletpddeF+cjhJuEAzuB
BAgVtLpLAl5jG9MzHqoKby11h34L8ucs/6sNy45OQ2YevdCJ8ZgTW3TcxvAV5eC9
LbeXEPBnHxy6qbfuU3gOLvHPZ4I4ROO5lj0l+uoFbNAOQ1NtflL/jsYNAbw+ZTDU
fDc2ztxi9pL0i7RjaH0ZTQyoGRYr73HwD9d53mvp1FnJWC+zogjqSxw6VDIvPrbP
OmLpXQAMC489U9gQC6Gw50sSyCRPwaVyx37SKFNuMkvdI9gU9cQrmT00HicRXBBe
CW/heG9LaVbEjcykFtLB8J8u9Cmr1E9ag3CnvzLtIIDirDsOsYODI6Ux01eQahwX
+r6/4tz7vOEtpX0Mk72JDMMxuEnjzLLn4E/JExRqfRMkfEp5VUa86aohM8RvV71Q
CDIM29540vLsKVkMm2lfy1yeb0h+q+M2DYXk8PxlahSBmOWu4fptE0oIMMYDHdvZ
ETdzsFprxdDWRhEhrpjILN511y/x36YnJexJNwPimI+bXDsA+KpntJJ2GiHmLL3M
UK87Mv1kSR0uLvgjgFt2w93LCIMDWK5usmXxmDk/OfT6Z7yTlopDupPMhOzpzdm1
mMRQsGCHHIgg0EwscT2X4pznFsb22uxOdufDwTCv6M2TvZS0LVt/+eiFFzNboNl3
8+Dnr7RToIZu4/GB9bKS30JEHe1mFPOsLsH2Mcuo8PP+Jsl8dQQ0tkS4oQuXGs6Y
a5K0j+JmD5Gp1eqtx1qO91/8bl3L9vPc1Cbf4zVzWrR1KFkRSGgcJVkAuAWs8p6S
wK4X1UOz41Fm3JLADYGPocklJT7pAkaZV36NWCj1KOi4ykcm6UC8S0c/PNPikIIk
OWZBWIVy9YF3k14hWGEP/bYS/tVqfP+s086WQ9Al1EY7iv6bVjuufCz0SsnEo52O
8/1rBiYU5kL44GLtI5rUyJCqwckmLJxNfSRnO1WHCW+HQeJOPnsCvDljHAq79aDo
DEjThw0x3H3z9OXXxhy7EaszeQDhw49IvSTvKwPXvEwE/Ri7+GVkUcQ50m+PEG4I
sKbThu34slrgw+w+/RakVucLJu8OxTGubCBrUvwh2zSOkQaTT4Oe+Ho/85UYQkZ0
dPmnQtd8cGbb9k+KewJ9l4d+20WsyG0nbdG/FYZ64nHlChRbVlF3wS6YlKQIZSJ0
UOWai+p3u0BXAxjCw52orW/Y8BirKDZH++bi7tqreEtbfisMG9nsSfQRdBJo4G3N
iMmGKL4hNU+iIgSh5kvSjUJz6R15pV9Vp837JIw5IleR0979bKU+FLve0+MFVNux
rKQeFJer1aicqNo4hQ9iXdWGTzKwFOChPK5B1gRwYEj0TRMkvL6x3WVJt4qRwABX
DZyKigN43L0xQAzucU1Jyd8fh40Lp+5jb8fjqZYeQsmz/usE2W8n5AVyvgZ53Ncm
hg7zklVOp5oMnPKnTXbg5S9Vy2afs5lQ+BRY6diNLMvxe1ylRvtwlQ4aILzAbiQV
MZLj63e3ZlNrH+SIqWpkZQxRpUKwPdUhfzEv3eStyditjUIHSKzoFuwM8QaCNEbx
R2xTk9JQ6LO0E/uTrrF2N2mBhQ21QWjNyeiEedpa0e+3xYW/i3GwExm08QQq0phr
n6apIpgBNF1sLw1016CyyvJxlUwSvUN21cjua2HnP24El68Q3TcUr3gbc7v+J7aZ
uQ9IZnqK9XHKhkd8Q4rprp4ekmOTeogzR5SytLKi98Qfbmi49TSto8CZg8ip8oBJ
SiraBLL76X3amU8LY16FGD1fmorrMbDn2oGiUgyN3QszCtrZ2nfC9pPreb8qOzZK
n2HIFj+xMQn/XFw8PhPukObdpDbl+M1Jp3hZ4yqSBG/vMbn+8MLZi27FzIpucaPb
74QBSwSbeLSJGrjKuwyj/rhoAIO54jaaqGNd0LyEjI7SKKLPH9QFOGfaGmCwfX+E
X/Ci8EkD+3nVXWTF2wRIlQ+b5FV7s0vlWv7kS3b+mvoBdcg5EuH8z2UmiTChUFFv
pQGD0VtqaXzyjtOgE75yAu9Glc+VEGe7xI4sWizqfZgVXbMAngmmzH3OaCfB0ocH
TCMwUvFerbu5s9GrgcW8EPF8lR/qIUceQzbroQCOIHgwMVhzfzHA9QJElZuEFkdc
x8iYaeVoIiwNf4OPGasQAD6eU+v9vWkr0S3JovROJ+NKL2mslWDD/CXpNcZ1FSJY
Mhfqyh8qe+qZh0tlESF2tRMS38lVe0qWI3kvXVvlNtL01ZKseJuJvK6FvEW5xdQY
eX7lgIbtrXc19bQ29yHM+gWhw2Em/PBTqkendDq95pkP9RQtcig6o858q5676w+h
u4tV2dkqenRzMkRXWS1ukb3Seqeu3mKa5/9X1S8S9hnChWhG4uFgbwPHeQPE/9pG
0Kx317eOVynjqExGu35D/fjDcRF9rKHwS7Lu6EOVlGv9KWCNLeuF5hViJD4P2JUl
kJp7I6tEqakLxWDH6VIm09FhV176iQmwq0jCfpG4A3wzhpBfC9oP90aYW0UgS1Nh
Wr0IVCCyAI0g24FWDi+qLZ8urW0slsezN4asIQJdEskQzzzntv+LJg2E7fHXE8YZ
Lg7KhBlVnPNc5j8cOleVdmMWyeOxat5G2KzDRKjuYiH6G9GIxjDim9taitUGQ8Fs
WGGNrolPJPAXInYB2AvaEVJPGBVogz5Zm33q/gZcIW7l9byTnTAP5W263XFud+3l
dPhN5f62ngV32myrUxZr6ob5iFUMNWUl4URLJsxJDsDhby+WM38ynrJc2NMzSuLa
nwgYIMSC/LIxplEDH7id3iO5UtZX351D8tWetqDUP+y71GE5PQGZffP+aC4olcOH
R6RmiO0awqRjH7+Q30MHrGXcOQkTaUmw9WluTM+/pzUGe7wOjcs6OpEskPl1RbKr
920ioYbfGpK1fzq7bV2H6IY76cJn7zJXcw6F88x+Zx4b8l0ZPJTSrhwb9cqHAWYS
2Oz9Z9h5HCFdg49m/MSoRHVhMl89fM7f23vZomD9qawTCOUjjjLUpX5F7JDKEbDJ
+1fiqgBYm73tBaWxPFiS97rzX915k70tzyY/QEgmQb0TJm6aHz0zRyaEnTDfnaU3
l+wN08bgLeWZ6wdfxEstRCkj6g8VSZGmkQGMgNt+eP0A2KARakYA8KziRn6MGlf1
XF1AkhkRcLdlYTEbW9WRpSoHmPVqrdSIjExhA71c53Xw8IzYgXcgFnFtJ8bkmJrk
OrlbZC7OakTqvBpyRACACrn1r8UAUywiXK8s4vgMFN6nWflCc0zITHHrTeAZxJop
qGCKGw8USKrFxoowdN0ubZaX9zVJKv9H852/eq4PgBYC7zLYKz3I8EzJ7fbvzLrh
vl12dCWUM72f9Fsf5e/dz9C3xTkYUg3vybmFyxOYCRVZ5zq1cTnCL0N/2KNhiNmL
yIU1rY23NgGYdESeeGHmZx3tgNLxwRK9iro8ZAgKnd/JmBogjv8BIm1fB6TZmdBY
XisagMqoraJ6rF6Ck/LZoMTcvEqi11uj+97fP8My+R2NwuX3+rXznr45H3k+naI9
32X3fNQxXlgRy5MgChExeJaP9rO47L38st7kJWK/tqCTJUi4XpojwSYXL3doMzBq
8rb8CMbZcikY/j8JPECF5dTsxWp/8Wcyc8GecEzIBcEFEX/G0Ktx8fwvLv4NPFRG
pT4HwmMLVOWB9tk1I6i8bIvTxjLE5l4uHcEji6s/wMr/fQBh9u41kw7RMb4EOUCy
6XgmvYIRzRPotVxHunIgN+zPmmqzsrIHspTicTRzon4u+0kEHEBlMnp89wyQy+Sp
wWzt0IBXD1CD/ojX4qsQ6dOkcI0mhmU0/Kh+xFlz5X3zuVgdbROGNN0RYnA0xP7B
8SG84ujnMpkLnZpyyXJsHRv1/maqOTdynARjBfYIPof7YHKGJsSeMpbpl9h9Ca0g
PN49Ckn2kqDh/TEsg2iyvSWcQ/+9ArtueW1sfHpG/Ce6kIDMsJxNnn8aBlQNLzyO
6SS6MCclgO06Aoy1TgXE5UOaJrMcO3L2DT8d6nzCYbsJg+TkaK22i45OHvzv1HSv
4SzYn3siVPp/kntZdnJz7RESICGOQeRWn4Zkhc6xTCFMrSBb+ireiQAMg5TBLd83
hoQqQJqf5OKngoWJR1N2TZGJC4UV44P5kF4Xcj8NeF6JyeN/S4DlrZtQmGeJQmtm
NOHmzEC/s4XIMh5Apkz/Py+4a95lXQ1D3+htgbgQeLFqdtQJ3eTGPCy5wEtqFnvr
we0CgSOLscEmH7XOvi61M2BLm/TJQD/WO0VME4RlkI/tOYzVPQ9koNnSUy3+GUhn
E8p+AqWofzlhKcpT2XqTcRA9T6tBboLiMSFUjoSkpL7V3YTtgCrdYencXJJXqcsd
xkfYQ6QoUolLOhhSj6mxFVuKtecKEHg1PMGX6ouLafvnGxUTgfqL8jyQE5xl9PME
6Nr7LDc/dy9UwWBRnuARLsgxhYZipjZ+KOdtWVJjF4ffzQoNQ5VKB487LYR3MhAg
O1XN5I1cN82cnJyXymbimbMzyL7CC5EcKKJZ918zI119sXbeGLF3grmVaUvxSOvh
tm5cjtM5tlQchllXxheSieZJ/1cIb5fVccKQq9rGJsmIHtD6FSUalEOq0PQLZSnG
y6x0p1kxIuzxnrtnPTq4VHgwz4+kKLHSPDCFkmQ2+uKOFKuQRJx0z3Se5Gmjxp9q
aRsxMrKiib25pWj/GkqYfRPuv9Qc/E8H46NL30G15N3rXooFmNeVaSfXAyZ5VE3z
YBOfRRVzuDLidv+LXASJWLTkcyGVEmwFgMo+CJZqnhl9u1DPhYAB9PWCIM401eK1
3lQ6kBgwV/Yc9vJAetE5e/HX+CSryJe+bfK8eScIeuzEXPJKyrse4Y0qktL7a8z2
lj5DKXJRXyJevrTKOHk7MmbWl0G/uOONagPmUlJlTNZ11vLokgQ0k54293zcBlbE
eVLXK+T78DcfNJr1ZjuZFSpF+6CDeoPYRClT/XUK81iuMkOCh2FO+IpaNfE3wDh2
3ifZ6HPZudDzdIXFuP79wX7drxr08zaPo3WPPHbNCva6lBxURSgQTM+se9F5JGt+
qr2T2lCihFixeh2vIu3h65CVz3AplXEStuFoqT7Yh1BYcIiU8+ZNdSSRzPMPAiUo
j53Fit6f5dS0fVjN44U8/RuivWurD7nsLsYSTPYRzmhi4wI7TBPaeeomgTqQyOtf
PKTEUg+Xa/wH/MQr88Eq+1YfXT5PgMxR+3BXVzz5NPYEHGOzzOHIiHL1N3Y9stdo
/rMNCTuOpuarR2PnubcuHH08ytomymWi9SwNpMM/tH5I2nOtyyqy9sjkSuKdwvVj
zehyzgrI5PzMvnROPW0ocpIgTRii+R4y8JuY82N9p/2D9DgfwCyVUaj5O8bU83LP
dS8tMCYfQ/FmZIIi40AkGn8deJwgPfKj5zr6JsHlRamFntlGuAKWpEwFXqG1YD8h
UyNDRnBOrAHXUTQ2CHA2eAdlmc8fb50GhqULh0U0abvll/DrFku4sF40x8dJlMoQ
XKFRoP2A06hOhF+fnFnaUFLWeJVxKKmDzndTlJz+ZlbBzEOwhpm7zMf/Q/AyLyBX
DDmCMMNaP6Qfq7FmeKwKnFY4Am+hUPWVZxjQsL+iofYFtZrvSs6LL4fsC29A7MB/
AOjU6UhVXpwfP9qrszV7VCum3wzf/6LB6REcseOI7aVNhOBXlym+2wHmrNv9D0A2
cpc6tOU0sx5P1vXYP7dhgDlWc++0daobTm1QgsWjLfUpe6+IV5wkr2ArLZPnU341
/tYmTcD8Mn4Vzem23vUySE6wiMQqWkFAtbTCHhwCihxdk1/T6iAf5nVM7fmeSrAZ
DPhXWGKOXuCzc3DFLRJ1HR8AFgObuGlNQE1ODJxezyK8q7DWKCrd4jFm3jlYYczS
ThBZ30K5PsqoCk6K5jC1aq0ZX8J4FhdsXTTOB1dZa2WeHvwdxNOl8Trxxrnq9WWR
+NL35Gqtwj615wgkWAC3jT5svQVqDfcBWi6TJSCPDH9ZyEPNcHMSAVuWDF65aiuY
0sozDynzvsylm+nqTgtIZlDAVV9J+ZLmbp5OXmbUSA35G2WdlbTg5w1sv0++aFeN
kaycpeppE1F078xTI3gxTMTJE5yEy2XbEBjIchOAsMBKuQT8W3bWtIlnmfp2jIzM
y9Ly4RQOzOHNoZXI03g4vVJdYYvyUyEViqzK8izLC0SPTt7XEpDZbJ67ipXXm+JC
IbnuX3rk+5qJzQrKPI8BtBckfLwg4jrT9XNvrETD3akc/E1VmcZRXmeJY5IAkGbn
4pjWqYeqBhXaFCScGNl0lXtYlGh2bc8sLmUa3jQiWoAap8wIFWUbgImIUc1HYT0z
tVWCWKzR7E/nkYEGIEpmaH/ZIll7JJy0S/VO2rEgXTdsB4WWqq9A/A9cjMzvl3fk
51EWxNBiuKRB/LkZbXysdvVDsOWMLEpTKXZlF2EcZ1jbZNnRrNPb9Qyu6UBB3NLt
Bmf4+uxSkCnz5QLnmJLrhyApBgqch1isHGvBOO7uGovBpxAcPmIoK5LFh+k8tP07
hoXXRFHfpXia6mOdqU5+jLITQTaYR8G4xoCyEu1abwIgtmwqrinEDbDGtAmBOAY4
pq1+JnLeGS01fqvyW+snI0KDoF6s0sSnP2nqR+77+b85lgLHs97GK1rCuU9DcB+B
4Sx/kToBSTPRl3MkGNXyWiq8WmxQUtnt9JrzMG/Lkygpf3QOUa8Zh3Md9tfuEJd2
EuUAGr3nsZPxNHv1OVhDIwJjx7q9/Ns5ettpXCBzCIQb9n+YHwtgLXiPPqOeSnfd
+j0RcXpQDJecSfcQb/1PWjzsIEoIXhNB2p/ewttbbK2pw5jxMCDtgXo3xxA+qvhD
XTAkJJ9K4kSCoIjiLYH/fFqKqhgNWVTduh4Z9W+YIoxbQYsyK9pcN0LzptbrjmLz
oxoc4jyxU8FZFf19YBzMfZ9iyO+Tx3QidoCLtBZ6I9nabny7cPuqLL+0XoTRjKsl
GtID/OaJK5HJLjMenF1s0zjKUokYKfbl4Ki69fvukEhZCH7Z+EqpAXKNBSU/1USo
S3JjGI2gZ3LjSaKD3zL+q7nUQbriOvlx1n63OgGWzUpRls9awTOD+e5hcfiqIUCN
0s2USTppa8oQnsbeymqXkRHHwYxZYNApDrh3taW5i2OZpikX5v5hWFTF07S1pc+b
6xIbEPARGqv6rWQVpCi6KGQMI68aGZT+MrQ5tCVZ/CglUPIEbVUOD+vsU+BWWOOX
6QBNgj1EU2ZRlsblxxyqNNu/rgcdK4gDBhcpblF2g+yZ8Z0m2C60VV1MONmKQPkz
qeVSx1pFuep2SPDymOxuOCmy75bmi4lh0zYXdLyPenQhZKNFYhf5hs92dxp2jlOq
yVAkqtzGsmIwyGCJLJCeFW6doI5NbmEngqzai2niIz7vqIkDFeINUKTz07Gjp/s/
L+g2HrFTvggrXRM8Ly7VpVbXI7XSMZQEc+X3dj9BTJq9II1ucUzPXL6ieBcYHg94
sVOeToBXWcB2zPlshF64KDlQpX+PrfBSgIfBW013Q8KtwyP75yY3ZxRQX1hshcAf
fe25spJDIvdxMvj0sFH9+eTE+roLKudCvtFhDphzOjamsI2kNDwUQUclXtrtSsjl
fnh4horsamlvPK0vNvQVsMN8gHDDGD0tYDScsZ5rpEg=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5lK8e2fwfkIdhH3oUNsEwsgf7+cbbL+23JxIDOE14mjogdODB1/lvVm9YjFpfxs4
ZkWvvkrCuv8kXvGWN6rXj5vx4UkZB0pUOrgQlgiQSgwujoKedFE8Or/bDu9cRCix
qKH94s6iFIJy+/m1jKvDJC4LZuTb/7b8KJY/pe3Ysd7HFs9i+BdNoVbKEIcc4hgc
Byy+kCvQ1qhEz0r0y0ALmQJ5cNe7VfVa59hK3jAo2vG2dVKy9oAd+8pnIAXO3xe2
M9DADvQwZMvmfIVqdPz+IoXNGPsenzGyvp8j6Owk0ggueQCr3lK9wJEgWj8q8ztC
aMmabpqgVO5RpjslIoYisLKZSQRJnEn2o447SwXZ2z3KZsSmqOLRKXGqXuvEwwEw
tLHn9iPKnmKz8PvvbxoSFOijC5/VAoJygqg/8Ff6vGSwnMflguERXa670rMuFbXp
rsF/5I990xPB+rB+iUcx0DV4faA9oQcmM8BW6xTw8udTkiZr8jYO92wHXhhTYNe9
SMtdk4X7n9UhhsC8LodmocN1Hd2Q8jreTNTXgpKU8t+S+CKufeZ4YQSERymcAGdB
n6mKg8PispIYpY6EnX3SPCESUDPGQJpHetSZ6onhA+VAELrsvsQqjVbMEHRf4Ad3
5cTA+Ujs1MhYc6uaQHF5CRRJbHz1+CR8i3282cWWtvIw7rDC1VROr5yJQhI6CFse
jYNLeOuGFcvxXgbtS3YBwvNaKgNofIZRnp6+rtOrtgSypt4XCdmT0WZWHHDjIAqo
2CuSuoAuLTFcCKUmrrg9oMqMK81UFN6f2IqN8+nsePzvtK8q22YpxXLwIhZuwq3y
zyrEpNPu21Rmth2ko+IV36OiOKm8UsWcaaQPH2IS7WogBeM0W5tx0FCfo2kiawO+
twJHUXq6HlGACgv12n4vsGXHOqtOtoQK30Os2o7r/QtHN9RVu8jQV/FZPTomOO4X
4n2BNyQqqkWUPj+K3Ek0ALmXMx7iSVEkNzU5Qm60T3Ka3SUPUW8PY/48+I3vJtxc
JJUerzCrJZnEGgrfSVw5qi/rdHxrHU4suNlBRrd21RbY/NEmieBp97jzTzx0I4wM
qaKuaBgaDfq+fRGhFav7/pthk+WW0Pa/qzBnjDCcticRGbYHxffcoZ1/lvRQekyl
0431RTNtU6wJhevSpeI48XsX7P+hwA/702nL0cSlkWSj5kpc5B5NhrytHEZilEm/
04x/nDzk4CO+S7cFqdua1b0yFWTr1YI7G9hUX4BpemZRA4Y0frQYXm3LvYRBZt4d
Rogl5Mz9B81Sd/cIWZ1yh9wkyNOh0hNBzVt98lcXLbRBRjYILLuUVlL/IoLdx36y
LBOmzxL27coLDCHSN3i1KBzDip2u5rNwFbOHA1FwAT62/zITYS9Od9uk8q6OiDOh
sg28zNJrGL9SfpL+pS0Sxcx/53VrUy2O8xUFTzIAWyllM9LU8C4NxyoYX227CL+M
I8tscuFUJDRvHDyYNL+cxg==
`protect END_PROTECTED

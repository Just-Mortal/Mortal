`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NeF18QalmZknqRjmiuV3yFswmSuk84BsdxQ/v4mPF3hR44snvPiZquyQi0pY9+f
ri+3e8VxLearA1LAr8Qc0FnG76joiImtbCjNcrEq1Iy0O8P2zXlLyPGnlJO91XMq
gPCZzAXSTq/k5wv426T7aziHL79dePrauA+Yf+AqYbXt42zjD0tMwocSU3aemz0T
+9OYEO1tYPkqRmRTB32z4DJrymcyI+G+mOVfQHuQsAg5qBRyKMCwnkmuwYA6Em92
AgHSsNe/HvrFgp56YYm8FRVgk8nvr64dqFEGTwJPfb9L2WMWbfMHxiLH3XK5ETKe
BSeS1fbkuEihob27qnBwTGaXjZvMA1TNvoEV5FVa8/Aj9sV9zwZG3EsHb9kvLUPf
8XqTmUQUYNtHzH3rKqFRSi3xllvIiVOmzE8bAdzvzPhG7pAmmHxiauN+SPIKvxNT
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWzY/uITKryMkJsmL8ftOvPhdTwZBwL5p+zmVSXo8gbOPo5uptMu0F2+35K7d2Gs
L+KPZI9IIvSjbZfYrlx2nGksroYeipFoZWLalb9WG4pe9jqI0hz3rbmYMZ8XbV49
J1wWp7I6jBihS7/bRvx8Yqmq7XOfME3zXpF700alcGU1BUrpUo+/PI/9EoxYQMtX
5VkrOe4ovhORKY/8AcroCpQLH40BYt6RFzBP0XPs09NYx28PlSt2RixC0SOnWYSB
wCwQxfERTvnYf0leczsXo1l+HQorD0Ga0n7uEURKXvso6AxLQVJpNrs/38UAezzq
XvYcO2lAgDOdK82PpCmkFdPHiMJa+qXgyYfMDpPy1yEd+vdKvX+lOfQy69uw95j5
+ULmnHS7TkTJEt59cMLuBpVByYu4SNjrt2R6ii8q//Vdjo8yxS0XHpipJtlrsagf
d2RobYlomumXlahWWBa6uAT0KONjNezl9ezdZwgM3p8S5IfLzkyNk/3xrDW7+zSe
zYX4U+cCHM3VGu1c2wYfChvJKOmhW1Ez/CcwVGFDkiAR5C9jU3FgPJTJhpeuaYPT
/whB7ZQLPHlo3H+5Yvhva1NT/lgWtMInVKWKZsPuDqFvcadAkGUFoMRdgfmaN37x
mEp2+3Vyu88Srdy4om8+R7wOj/wC1YPX9WdFHK7vKYNkdVuSSBVeuIaRyOb1sPmr
NsDLH45VGJ7HFuHRo0a1lt3pDvi0xMAlhYp59RHnylW8iXR5ou2mPYxHDiSNVhRr
pH48SU2+UHaRXBW58wmloN9w7FmA8pyvKkGh5iGQGkkiDmQR8nxGVb2YDI3VLF2P
5Ypovth72jHRwro/o+cLvrQSzycovShhzoJuu8Z/YRPbaIiRf4B7ufz8G2dFIvSo
36nHvvXhqXtN15kY/vOSj1dpJiXOYdnSpBZ4IZJ9Z69CDymg+yEujMEC9pI/+o6s
pO/FWs4I5hhY6jHYcpQ/DJ5UWaDAgDw4Kuk3f6JvToMCUHkM9rsjxL7NWTJ/fzTx
1kAceYFpbhzgJOU8pxmz1uyiJs6ybPb6RyAVWB6Wxap0a3M5aYsV2N6XlzpA2K5q
xvlSk+l/5Em23Wrsc0KraKHOpDracL8RjT5T6E8GGDSzXDUbrKb4cDbP+ERkNZB8
FzM/OVdMH4abT/z0gYV/wAtaoXmtq3gAN9y2RdRs8uY5a/f/XU1CgPfZFav8tu6V
3VuT6OoB4Vlmp+nU5LYQh4W/mXU+Qr2kr5jIfcW0K1eG7UdM/1aLsE47NDwJLEp2
FU4wf/DGqdWL6k3l7GiQq7P0ACsdQwDhHz7R1qSNGOmwkQZf/ySVIPMTC60LGK8+
y9psSZIkZQqmWsPfTlmToiYTWhSsoeQ3G2ezRElDTFwbd3R4blEaXYbyTPhvcfrM
lhLF7xv7BYzvMFt/H/iY0mRLruL0p6lCLO85QXlb/7Vz2tORzW7scblNPPBw0YTe
Nkh+H4/3qI9UZW6GK6XuBa40z2OyAF/bDzcQuZJX3/SafSvqECgrEDd1+G3b526Z
m6SVTJiivYoxxJv58bIS3LNZoSUdQTfU+uMUsE0p697UeuRNmPrQUFMMq8ZBiqEE
BSg9sBipgBv08HITz60Of5MYLT/xtPAJ7+mS5ldEGRHWVaulfC1NgEfk5oBR9Wn4
J7KgNMcz3Sn/nwwQDnWA2csmBlLlKuOqrzhbACvwm+Zo49bvaFRVnzRwwCHCDW5A
0xsEQCYNNxHmN8C7N9h7oCiMQQ8na2ZzGT2tm4MPaCB1dmiQguEOjvDdwcDizS2d
+rxnQY991mC60Io8XVdNJe2p8zm1hrdT4zuMxnxbYCshhRiVrADz12W0F5NtXzGc
jUB97xZtpAoD5UI14NDHsNup/zYXKv0qMCDwaHlzyn3K/c2f1YkBqRYeMiMPmL7F
7q8F4EU6oTHIiCyvAS68RGfTduZOQj+0CHb/kCNGPF2W2pSFNTBAFf4m/gJ17J4X
IYoO2994AI+EfJX9OuxlKDnzCTK9rdXG1d/BnYBec0TpIWmKZ0I6uHdZev6oiRqd
hAZ/5A14PkxjkCUOQlJ0nKdZU5fFYXnuqRK++hmPUNTeSHzo9Z5vKzuo1JXpt8d6
5RcHsPCEjVV6vt0sTk+tD0MKZon37oI+7vty3occbtG0qcN0EUUdzW0+n/tWDkNm
YrLd7dilPvlRNItAlS6fu8HaKk58Ajq+hat9i86lKscX8T7k9zZQMHmDoAirTx/T
T8n1w50J/QfIBWVDgAkYa2ioOeT+25NgvpW4aOZA9xlXUss635e7KP9Nxyidxx9D
0vbK6OmJtFAN9nGixyQRYczpvlUujMYWLTb3lgGWqR/XjyaxKZEGmp8olAgg2CEH
mvJh0vUuCspu5iRLUBEe8orH2RHpPq5j5BpSN8KH0MUtwL1voSHmnMh4rqt25ZlQ
AsET0IQyiTJ2t/La6TKyzW914o3epFNvPuunjCnflkjxJOVtLfHxPYqfDiuWabSE
yTcJxP0CHbargqbu8Ec7LHKMzF8azBh9R/In0vO0Pd6XUDrS7JosKzCxq9AthWBp
tgsc1ez/Eu52rgUcjqr10oh4qY1TSgCrP8ibg0QBF33BN3bpKaFAfdXzOQC5btwg
+qyoo+/JuzVMpfxI+MWbboFcSkDEGFfmNzYzBz5qziRAphMQinjZjNbr7P+Milsb
KvtE9jvrl0M7th8fAphyW3nQGEQgq+vSpSdC8x6RPt0fA2DTwGLY6QyaFQ1yF+nd
dS0UGiAH66M8DK08rnhCARIJ2oREpAObvZTJEYApz/Fn/sN2vRLpaqdPS6OlF1gK
jnwng0yubQprvnRBy5t4HSGCyp0Eia9VwERbOaYpU+AO7lbUjIFF8wJgHurenZuq
XSDtdUNvGnOSFNf4gGU5dLuhx21sZweSveE7wKD3yfLqABK42ZiVXPudjkaxozWQ
2gIP7SDr6D5NOrI2+Fk0jAVjRYLyn/fQpWJeRFPfwN2krE4iXvaf71SlJFncHatg
FE7YFWovygeFfkUveaq1KH7e2FtOqSM1dXT0mXPed0x5BuCZC8YMvaDEj8pD0l69
KR7tSaws2KoL6Eg85EpGjxHMryLxRodGc/MTgXWxz9BXYyIMokLlSZMEfi8nSw8d
e3sZgQtDUr/iQbAnHolWCN4dMwZkLEeTgpHymraN1aCrVCRrwwuCWHv8xAf2mI1D
tah1CRu8zzsxsoG0lD52Iws2T1q3D7ivZZe0vAIS/Pj8DXDnueOrw61NnhNSS8hH
k7eds8ZtrvvIUwmqMe3DWdr3gzdnTlypa/iA3gSbgjM+TJHlcmdvyrIeMfKihCXg
cFaRsMCNDlLJUyou6XY7HiNZkUAiI6zGtIUt/haAMpRRATp9WdTUQSk9sJu4OAiO
MYEfxtbhf5FceOwPasaWAw66HOM+dKtMdq79NnhmRA0CXFrbkvWBI9MOiqqwlVEQ
HUI6s5jEkThdkfbbHvAifmRi8USs+oFG5EdqHq+ZeVCZeojII53uvClCSSWMj0Lr
tgSdH0Ns0+1mqBpLRmvXrLJKEHodVAZJrCKv2gxNZAkkzjZ4JFJIO13i4iK5eG3w
EgXixOAlEj1e1KQAS68jCvM8/lLqprqw2J2cUunVIle0ta9wWFnS7p65/+Bk7k73
yEa3aUKk+mZh5WkUTOR+to47MWUWtForV8Oho7oILDYhLbEXUDBojV0PD9l2us63
kCcUkwiLlacGrIYo2dOyGyDLGjyANK/RDn9a7U/Nm9SPP9XXC9BGtGqDYZshVNzj
w9aUSQUy1ejF99rfSG8yzsNOIlhr+9HDLvyBXASw5La2CkU7T3JpS3g0yUpOCKb3
fc/ieWRJEIYbd+V3P7TwDhTziGNSzZHf3BcT+aBuALXQs1x01+g9Q9g1aF78k0Ef
SD54nn5sda9GV4fJExe/SJ36g1HhpS9mBUsrqT7IdCPn+JyCk3YaWV0Fjbmb2SaL
VUZAynobaYE2xFvYRLqA+Teu5GYA+/qwHUERdhWUvYdPQjXNzCepTpVHmfb89n8+
KhatnMlxUg2AGEj515HFEdlOW79Mrf7pX4sYqbwF9P1LdM1l9mkAZbyh2C813rGy
Vy95VU44X4j41Rkd1E7nyIf29/NRVy3xs1HJGXgWHFq2vUlAibeaxJPBmLFHLNM/
P9fMGh7qK44XPrg2CuYOlHCfYQeN7wwfw5m6e/uXAgvQx7EpRHcZN7U8DHHq+SDS
llnnExgpT5p5DMz0LoCYuzJwTQqvqpzSkgqOUPBht/ZRNNqVuUxT/hkRG9aXq7HU
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7LQdeMmnhQI5oEUnAdEG3jpC5AoNxz4SaS7Oqx8jW7743l+EJ6d+Peyom/iNHaL
J6ipkcGhL71QZC9al0WdVu/35w4iYThnGkiMa9pmGWN7M2ciI3P73VCLijmzgqj+
TqDgAFBUJHTdRC83g3/1vLMdr1QmlyQE0lvwMwQ3Pvc4wWY9pGNIz880Tz3AIHCN
RTYoS+dofXl2p2Akm0F/waIkiqOvhLENM5KeZUhX7gA0aoEav7xK186dk5MkdNeI
vYI2EirkPaBXTdWUe6jvtROXUi+t+DevJfkvdaux24shwTs6SY4z1fXskOWuSpF4
8JVrr3+eN4y1yJ+V6ihB64u84h/sGFKCogtVXmlQal580DRIn2pF/GtMvD42+Q7z
JU3k0Co7Dnz7hl5EUbaXWyZOMUSYL3odAvG18SESDrplScWRN8WBXXxTBPgXZexV
t+elpfokZtbf+G9cdhmT8iFnARYOZ9i0SURkHbzjX+1BCB7XoD3dNR2Rg2CTNbry
WPWseIEA0EjOehF3E5CDev0ktHLqhUrnU+v7VU1RPUThqS6+sd7ye58VFPum1LCK
WXAr0hIKNhDRqDae7R4KN9Qd3xcduHF0vMorJg+CGfK+YDwvAgIbSykiNOMoTTAZ
DYy8CGATzxwvLjxpD/qR6ISs/XnkPpD68Vp9q3wUWi/OJi8GdOCiCpeSalmgV1yE
rGvWhBEEsameVrrCn6CLgBt0Rb0vsvF2cqQYYzsE8V+1RnF2JHirjjarUdDVnhVb
hXfCMw7XJaoYRO0xBSqpQUsMkKh3FPcbZFJg9ut1wI1g87lROmZ1/1nA7K91Rnp+
VHkvJ7gBPLLkK7iNHYVhYQ55NxlyofPllt2Z/vAyEkAiPHO8cBKno7ARJgSQsOES
zswR3b1PMKjadnAYew8BqK1bqX/wmNeggADP3CV9QiHostdQ24UR7IOYgjcAc/we
N30i9RkbO6qPyBuRyEHbsUj6jVcMge2ROdKzhkHV747lEk6+MY4L8P/PVQkQFr1u
ecg6G2ZpQC8XIeixramuOvPXN1ltTFwk0w0NHBbUghFrHOqmYZQrwwWWNsO5Sfuj
Zd758Vkiw53+YM2m1ApenqvYE03QOx9L+H8ILPG+6gk30v7f6hPWBRjf6Hi+xmbG
YEC1EhAAQZz/MdNOTvGlARHCeBjHu19umKTFSrTQt21qkmhtnR4UILTkBuIqE9tn
de2TU6Gi7Bemd7UJO/B/l1PwXrF11ORVv+kykxsu3Qas9wqM6UeuMY/+NapcaHGe
ZCpOLlfNKo9lnJGincrTN3kMmZoQN+2Bi7gE7OGF31+THwxXK8cI+rArJ8IT89Nu
KYQo+tgy44G0ol45T5J0W0HpoPF7rc8D2eVFO2gulx+dPfaUDphEwsiG8gcOb2YC
vY4e2iMh+QYT2AGE4a+9AkKuZjeIalpz7EsEhEWA6zah+SA1L+ShKoOizPruZy+A
Rl2jh50ZZG8+1NMqMMx2ubqDvKRcCU8ZAshuI72UcvwcjW9q74KWrDjDJ0dvR/EG
tDDOIfvygwE5GKjJntZlLb+ZiIRP7FE7Yu2PQssDyYhGatKKEzjN0P7R4X7ljuc3
F/ZKjHxoORnSWqTOXFeFiHWrKRktgI8DPvJT4cKGAtANJO0bjWB7X+PGqk1YO4pJ
m329nLdZBxILlmClHASWZisexq2cc/SMbmjeVlAL8Rqd8t25IVpugAvPg05CPsYh
fLOOOqKfyev4Z8d/bvITeiBCIThppLrPI9OJN+5RxRgZDh5v2gBtOcLZkQLLKm7Y
dOjbwhdAssuYYOuuTXHPpnKc9Y1/Lwdoj0rHAlAHARtIMgvO4SsTs7eO0gEEkGKC
ipRXdDK6oq0c5gvMJtMSRTwVEWKYy8agPcmGX71OQI+te1mP+vzw2mLgHnIw8GyM
XISHdoNsa5sYnNDaVQazzd4pjY3gJE+wO7nxNwp9zJVpWeWEcVXRnuyja9yxp3Nl
XNabdQMuvLMFY9U1CzLSzJy/5FUwhETwSTYYdPFOuyZ+BUjDDAaRxl74ZqK+jEOG
xkWwBklm5+yDkYAjhw9/TAEyWhxKfwj6H070WXbFK7na8UGrEHeoTP4/2dLjO4PD
1mAhjKQ5KUb7q62Nfy4vlTZQVOR0KfaxDVilnjdH6HehRYg5zVw/h/8runHRmcdo
ZggLx0LZqV9O4h5ehj/YfbT+4OBpI9HwlGu+jXgrsjZFeiDotokApk5bEYUgQnz7
pnUUp5Ss6GjIGSfFQ6QT4E09OYM+dOCSikBEmZPUy72euAzQWWBWrotlCUgdtdYD
2Tx/OhsSPfl7GJjZKagPRUsGuCkA2+pqquQSNFToX9tivlYVzl2lpeMMDtyTPF5N
Xz4iEWu55SbhM+iZhEkaOdOM2g3rDv4Bruq9sZgrXD16x2jujKlmzafFyuoE+OLI
8lPBT0UkSdgfrn6c3jZ8F2EV13FzB/rG+od/pCndxkIkYO/ChKTiA1ubJLQMey2+
7GCToADMeuaDfwQRW3Q1ZwGVEqjHZ6C98cpL/jOMVTg=
`protect END_PROTECTED

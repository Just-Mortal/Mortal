`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qVYAwCmCOEeUutyXQF+8NFW8XbreF4NsCsSFMzfHuqITEVtF1RugbYShWbJd12Dc
s5/gjreqnGkVPVd5gddUXjcpGj9z3Hg+VtcaTC/5isEx4fBX2Oy/G7vc4mnF7h8Q
Qm4ok92EdLJi9MTzZS0BCa3bt4cECrbvegJpwWyjIpvoyuzch6B1E8RDLwWebIkV
4AM+Vxuu2rlZzTB3vkqTm6+LBbkRMgEWMY3uEVyfw/yGcxgVEU9s9jggYzxEY3xR
B3v2Vyi08QjEZjuYpXTwjSINQxMu1vhEu023sKjTktLNcckN2mYofKLYaq4waufI
jmA1FghU6W7/K8uq3yevfrHzoaeIO4lk2MMHmrLvhTQZ1gAlzQo5h1ATm2mLV6bf
Jkq/9I2GFV9gCNyu8qvA8VwwomWlSGWhKbhyATR50HBrreoaP4d8jZZhIcx69err
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21oI/Bb7HqSJm7RqgXA7q/NMZLpfAtRptfKLapDkk65HiBYD23SPFon8lziEKkxJ
uGa2pdiPQNcNFMAlmp408+g2HhxXycnNs7kXsIgLE/+or8ZfWGyU8v9rGEwm5EdU
3PVmpS8Zt4B3ZrvjeA2Mh6klEVgTcJ/uttmqxHPNdJFYayC4z5meUtDQgXoUtb55
2QodzPlXLPKNaMc8hPOFTLvH75O93CHx3aW9gvSebgUvwkgLwxT/KBdtM2OndquI
IFIInozVaHQAsjtb78GSbN8dq72VIdNnVjBmf4ILMPFJmkmd2y3xOvv/hOM0frlG
dPnD/aRSfFef2R97ik4XDFmTj5r2vJtOyhRNmfIRpw9ysW/uXsZXZ6nroyt/oSbw
Jo0o1GlzauCrV4U8cjkaURLiOcfqUjYRXc8okxgeuP5vgp7pVUDwc3GpmNbd0g7j
D2drotoUkwqiC27C7kSbtxhd9yx9oIYy+rnFVHE9OEVG7BcsG0MS07KXGGM+OOYy
aF0oR6RTkZF2egoe2gJtvZWFSpMoD6NwhC0/yKgIA6eQ11d4cjYAVznKo5NcluW8
5slkUr9HvBdLsd+8L7pYmF7v1MTR8hemKjeYVt9LUmuOV+diYaa7ldIvX8yA/RFX
3HKZpfUt/p2jP+/t9O4ddWqn/LMijwuT0PCgu7K63jgtq+H0jsgI3Bu+BaAsrTx6
jm2T5mV/olLVIi9YwJWN4hDWT2IkratFq3FnYJ/B8Afc8wqRa4AcvISXPFKATBw8
tSXyWaPHxqS+YJOu1qPm4aIowm5I5WE0m/LUySj5ZufM9PYqdjYaJjSicuqcfs/U
YQfy9mvUdcE/+y1aJDr0YoccXpfn6wrF0L5w7pRn0/yESnBlXKDdFxPdoGbBiGT2
gggyusnVcc2Bqoh0Bb/6LNs47hE5Y8gHAOlqtjiP1OdckrvVel3m5kAdaTJMZO2b
NcfiW84x12XFzSq13TgUivwPV0M7G6GUFUZKeoOqW4z4bJ7mubFOREucFK8z7TEZ
cbe+JwhmtSGk6f6BwZCxapH4fP88JgQW+wmrYQc1ESRMDQ891LCqZGdAaz+VmVTs
+aKVroTBkcgh/r6k+ozyQG5Dqo2wgVhdrwl8KNTXVt4tzSRRFUr3uXYsjI+6PDkb
Lf/hxedMlODyNZ8SMFt2DS408Y6QfgRMxW5ZNEOu2ItwrLDfV1WzccjChV/BhnN6
UQx36mXwLDhRchc68Flw07vpTjbrZOexgxNSs5Om8hy7Wx4bLblRqoN+IUQhcBBf
oYe6gBFFplfvYxvYaCPpwj+BR6Fz8oTcW5Lh3KPgO6MecsWZDk/CeTrFScJbE1sU
OMaNjg46Or/O77e+Hh+CZFQ9q8/TG3zAg8FUIrZI22LlET3Ao8pYdSuMaP1L9xKn
E01v0fbXCXZtxwEfeCxkcrU3KdtE8fD0TiKww9CXSRNeC1hkujLUyPdFCFOPYlvn
INHnCra3HU2GOaRM61LCLgtdOmiKU7I2Ad4OR3RUNHKcqrvcornwa99zUDa1QAOf
3vffMRbp8uowZiWu9LUu4MVTYZShWfGS4sF719z66W6jicJtG2136DhHbOrOLG4r
GNz+SNvt8+9hldavHYiI4QyKXMNwGRUtZVStEnLsrCY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v0PaFDa4XCwMoRPP2SyGZUTLT/njTDcR5TgdX5X6+ZE26Y2DJeo9hCAxtWc9zWGA
EeMWxavOenhZwNEdtLrzbpMdRCCoF19bWRP7Kdxl77EJER6A4zmkiEPEPa/neOBS
Cnft2VrB8DZ/oo+5fLurqZqRcTQTYTqEvzV4UxJ5FxkH7BM8PMT/AXfeUvJK7nVm
EcpL3BNO83+aCwxFDq+lDiZySY9SP0l5jURuhKvULEzJgWE3+xFX+pABx4fGOU+X
p/kWY7q6TgXFQsS64sU1GkaIUBXyFeQ2c/PHU/kH+2aYkIRk7CQplnh+X51VMiPm
Q0MGLmGR4zrgXrx+gmicPEHekzwMNYsiwHN7002toUlATpOsaoIPd7Iziwq6EyTA
qG7EW2X7FlM+W+MzbUqW07CTZMQjhrxwVJSe3c4Z0/43P0cAHdZQaC4+H3xd2HBl
hB6k29LQFosdTQsJgfx/BoGF1m8OwakWND9co9OvSAQHKK5S9axWLjwSXOuP9jpZ
t80lQ1G/JV3ejm7c/YFO555ugtHsyCjJjQdG+GbBB0/IzdZgcU6jjhJ4JiYAKQtV
e3xqFS1Hq6+6uJ6FOID6tMXwlFHKBveWiQD3G/naGkP0TA+mxarVSzPjO4Whgddb
2D4rXs+dbgBYYHA4D//pa9WjQU9cWJX1VCALB/614i5kounSX/ViR99FCfgHz67b
9M01yIYInSb7hV1kyBeWkXDjQENkGR8IMt3lCyFQTmBuGWn1LhlUxi+sMy2zoTrP
oo61guaOhIL1B1BrmmHhaVbCJxwQcp0aPSpLEViKZ+kl/Mx6nQbnewJ8c2RUPCia
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXHFT5QrmdJqgAKbF9ha7gb0CxI0Wni4sSed5wcgmBuiuMwuR/gwOSwTw6XBBAI7
ZPtmHiR/w0nOkoTgb30CL0snrn4zRhSwXJOQMmBMcglQh8wCZDEgGLapScCjmoHt
2Z7LwR+PjpW3GwFno28KuNDLkBxlPqQosVG3u1W02hm0dTQZjp7njxxhUTCTXOB7
sPts8XiIi9Fwg/DbK54figqXzvfat5bHP2eQQu/rk6TuQH+7DG5kneztE8oHi5Ok
yKNOMUNqGA39hJOsR7WJWkKFEUKVXTYLIvRak+D5btZG1Wur4McIn5WjEfZQPlTi
/ihpgT9r/pr5QQaFXUeemPwzh1DlPnHLC/kNCH4uQhPqPuQng4K+sImrhrYhi/0M
8J9vjm0Zp5JeW0ibg2eu0vdydSWw+rc4Lf2+RRlY/Ii0KvtA89Prk3hJtB8FX+XM
yq10sGs8nGq2R1Ob4RzjXzMJLAq561/0dj2MpzDguqdFPdrtvGBhY0J6g7WBoQae
ZGDgnl+1MAhszBPYvvuE2HyCon6UGw+CRE1EkjPSzcND+bPBJ451wl9j/3SgCVSA
yq4jbecADN8FTfyvoJqGKC/1UKQi/eYeR056oYHkPMgaK9F3CjbYAuoMFQp6BZ3q
VTuQZrQWbhRG5n5WLiiw7ubKwAOQy/M84gwsQHbQMa7j1WaBieGg18NwHg80+yI0
O4vWGLFqc4YGagl5Omg6ewiAsMcAPQHXmEybLUXER8t6KkL/PGI51MUzlrJWj4gd
w6i1n6pysNYwkyXbhGEs181iLKJ6SHQg4jWu1WGPjQKCnArfkAmlx4btk/meqK8l
08l/BuFoTJyQ47Q8o2ITF1TJ+HLOM3M9MhoYdJUsKh1vyVDr77VUjs9NJlta2JYo
IyZDb4hFSqPm7LgRkyYozpu2gNShzqn+H9p9GH/J3Bd7qjvn7J2x6ao0zLOask/g
/IsUZ0FZHP8xbNsO/YmM5vubRDWsEAnr/4XV1xmzIrTbAW3Mc/Jx90buFqmp1yd9
F9YQnufRVoF35X1lef6MOIVkhBLApaV0SiX0HiK9D6cerjhZNPlopXrN5pO1DOjr
7su7bTwxX5EjUCdqDl8YpLWnuY4VhFJkaHSTFJvEUi3ccYVFSyQeYl+mZx7n4/ZP
IfPCJdOpI1oKW5qHtYCc5Dekt3fCpFbyptCiuzMMcI1t31cBz7kEOlRJ2qPI5SXm
H1hUcoRICbFX5/LqvkbVUkQ49KntxwFIzZ2FdfjBTWya/7U2zI4ZP9o3ssIVFthk
VBWXipP/dSpcP6moprrZa1XGhsLmpRsl8Fe5l/tog/c6yUVGQsRpFfD/izk0upw7
h0A5mqOLio5luTUo0DReuk96UMLpbwUknfVuSYzYETjwd/q1jbEvjDAYfAApXJv2
SaWINqrFuwU1cJlNBnji9qZ6uosV1AjosKKXVoAQPe9OHhSI1pwXMCPDEYRwKRPC
zS/fipcxk+6BoKF76HY0G+vEseDU38s5jHINniTRyEbGBiYAfbCWVhffE3HC/fDN
yAkGYhpKhwi2Xp3mRFoVUbN1UF2Gfq3hX8fYA1Rbb+dnC2YlsbpuRDFaoM+Q7TC2
eLTIVIBIY3eTI3Cz/JB39FlbR2YwUYER/aoD5m96el8Xp5Sf7a88MwtbqVmWoV4s
UBrenorFl2f0vmcNAbi5pVPY/5UZh2wiq2h5tFXmpM7QnsNfGJZy1BSr/7XTqMZ7
baTPlTvQmF3XCtTOt3qfbM1rnWqZvQuJ+GuiwQM4/4pKJxQxmbh4el/MSoC/cvJk
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FsSZktwlnGswCcPVPcSIjj8T4RsrwU9ZGzHL5qhoy8m/pS4UacP5rW8NnoWwAVjO
jbuBp7ZS0exrh2nCAdnfo6Ybfw2fuiqKWUbsYYeVzEf0ibP1tPj0zrD53rL1y1c8
gmyJDHAL+sRQ0am+yV836jbF0NXN5b3y8Dxp2r4IWCfdsmL4wX2hnzihXpW6Qmgq
oS1NNjQRHZIeS3XQhgY0100Z/DJJDxtUe4jvDn6bZUs17SHqUShX21dfVKiOl8tF
qaO+NiXUrMRgcWSFECEQB2I6WiAlAAKBNe+Gd0jNRZV1mqGfCqsVHuBeAnyi6HRD
47EqhdWiSkFLiTCFss/wvqxdISYRvEUfPiJQSnld+Al7wHqXzastZwN3WX1hI5jb
VzWZItJUZP32EqZqnc9MX7NQkKDr0qyrrP3dl3b3PFUDdgUdCbrtDtbb3/SIBbHf
5L9ziLLT+64uYgSPwmjtwWnk9AroBDuwDjXqR/BWqmFypQz6d/z4z9e8irmM6lfn
nuOftXMhMNWkX5rqy/1RibhXoo7kxE32NpV7u6clHG3/UCcPO1IaawxIYvqQ2WVC
ikzDFeG/smxaVZEdYYzOkBYP0lTLnO9EwZzmabshNtrIFQ5YIwyrHBirciMDO7D9
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9QqDbgMMLaZMFCebdH8qPgTL+8ubdWT73t1JoXWKwFjeWdb68Ret5813xxyhGPg
qDsT+yK7wfalDKcNeSaLBPEMzN0Ny2sFVuhsNKM2M9s0HHOMsZ4mR+u9K9mqlnHY
sZgJvSKCFMXnZ7/Gca3Ey4nbVZ5bfy9k2STpy+g/eBQBEfg2BS+FU/TqApJa6B5o
BtNN88IQjt3ElEy3RHhw3RwehahJ3Xzyt68H6RbkPqB9dMMv/YJ4VFCYsyFL/jJt
1s+0OAmFX3TKZP8UiXTDIGhJYIb5iUeY5VEJiX0ECW719DtwLjp9uWIw+X04mYBd
Noza6nIAhvv+K71owZSvMf6EM7S1r3bj4HTIUib0akNK56G3G+Rvu0KqJRWQqldK
ULGRca6c5EdpCFk2bvd1svkMzxhSOZe3N3Ha25VggRqvrDrK9X6Gmf8bN9kM9efb
qhFV5T8DuvBFmqoN2Ty70CO1R8wkTpMkgvDUGSWv5S3rb9zXKM7jl0ja6Y9cbNkA
ayV7rOQi1gs56HZ5aI4XtSHQSS57XLPs6pPvYcpp7mIIM0XnLTciwOoi4jM4sTjw
D7DCKrSiWIeZ/XCWlck+IHoZzNadnUTV8Odz1AcO5EjfbLc8LpzyJWdDweZMcsG6
LtzyuRWMTYeVc8KMndjJdsuIvUK9vhg4eWEqk4h38LyrkG64s8/ApvAMBdczyTgA
O0zIK6iR+1zMYyzZLncOX6SZDMFJYPHxUuiEhRwUqnrjoF0lRfEuflQD8BHVR78g
OWe34o/N5/LXB3nognwZ8y07vXDdB3vQ3p05fxFO3ajvKqYNtXFBeBK5JOM1F9Ol
Im4/WZcSyuwoEsgjimHaq5H4i4sGFTIFwBmRgJ1oaXBpsaBOeKxQEct8PMHBY6+q
GVRz0+/a1lCXfzP8VmNbo60/u1UFS5u8KA5F84DyZEWN1zCqL+8Q69J4urHmSYv/
KpCX5DAETYzy3zMtTdyHmq4mULPi6cjgHft7FCOAAVU0kTLrPrcKMc4a4DQj/8/Q
KIWyN9yZpcgupEVyZ3Fzg5nQZkPUB1Mk0OuqHegMxTi0XTy6Yjkca/YkP5M8+TVt
f/esHlVL/qFYkqAazpw3mOD73orQHXxjrVCAGquLgaWucyxZwYdsa+NnZOepcNLe
G2YszeufwEsdZkjMjBME0INyZ+x+CtbcgSYF2sxbIOAqArOwoclXEvtqTrueUvKu
YnoM5bvKE0GHGkkB8fM37/dRnrPTCN3qjiP453VqcIsvva9NVUWwRSsAh5/vqVeI
WQjVSosBdjXTXgh4yPvedLFvgEElD55WPHYmcY1w7dUNlh4mXjJ9UdI4mVqWMjfc
7Gu6AsZhSfmWmyorD4H8rkO/8IzM7LQ1mLYT9IrNxRodC5tLIUjUeMnA8dkX9c5J
e+SBhUOMK3mi6mZvj7CQfVQZVnzHCehxr/hCfqPZGNzcrYzIYGO/ejuammMQVBEG
W7sv7EvkMyMzSb4ORyq4uuxdPTlPV3hRdKdU26VXwVLPmfMCdJg4+GBKEEtPntLK
mIhd097cR9v5mY3zWhaZo89Okj/7LHopJnfHiD4vWDuGwRB7Q1fUlBR4ytq3dGgx
uMRX2qlQUzUUcG+3WH7RA4YJqImDFnaucAkk7xxMF78nxzjKW2dqItVIstQYdNXd
pDm/fdL2pnL8/exuKn8G6c8psg+uSJ11qHKCGMJ0nSktnBDnWHHvz+Cv83npAZhO
9wIlO0n8s69w3BLzz5jlXzoy6yWdKPEyOts7I7ZtxkbTPrpl3shWnnDp+hjqBdwX
+IOBXfhpSW1vYm22EgW5H8Z9LTmMfcdf643SRJochxe4he5dFpFmiNTm+PrJ87ER
5z7b4X6SOOcPZeTeOSkFduJuLjRVB5YuCSmtGkcf81Y0yW8y9IhCK/FvPTwbFgRp
uNp5htW6t83JMhgGzAi3i+uf97RXCXFpaWroXG9G8l2+t98XN5tNMDXVP7huipjH
eW5HQAsbFZMrkXpr2kOFGeQqerfNAD4GYxkE76kXcP5dLJzd+xcD71im9PEw6tUA
OcF1pQzj7cJwzzgLB2eZJ/mYgWMnjv+6bfpR0JWPWDDSOGiguD1N/tffj/sU0Xiw
E5MZyTJL2F5ocbEASULQvTPv92ETh3pTy+c2qChnA/9pmYbKOBJiDuQkgJJBogBs
8YLgUXsJAJBBKxXOtEVmjtucBioUz/u4gKSUU77P242mNWw7BxSW3qpp0Gavwmy7
B3mh/Nf8qZM9vOd6bteoD4k58//1vdxhwivrE+vuM857QI6K9HxaNPxjdyYb1lf9
1H4ZCbJejuW78Icd0cmh+dGwvmxS4HocY8eJr5CCd97VkfUC9Fh6F0lpFub2wAQ0
t1Wg9mL93KeXenkxsJ7pWINWexfYgBsk4B7Q6CE6xl9jad7UnUi9Cm4TK5pDE4t6
Kg/klu+JqV8j4Ginm6NgH/hOU9p1JSpNNQM72U43TkYNXDDuFcteZxrjjgs18DQC
YEhxUjwrd+jFZRawNv6rajrnGli+7G7eNaDnXRWCRflOGfYIAXJ7gjIm4hN53KKP
oBz1DJmeF/gf5SKYkxeoxHUdW5uary+ZSbP0G0jF4bYseb/mgHZSfUIx+D5wlSWm
W7UxpeLq6n3WISHxqvgovQ0yk2xbeaGYBOyWT9ODtwkaBsKbQyTyLhLbCka45E1j
ZnPIHI/p1MMcbc/cM9nGSBhBo+hoI5FjHrXJ2XDVzPck/7fgIGg6VcpehUnKrytO
SjM86W3T1P+L6CkyAM0KlIcj+nwkDwzxmkWxXmDjz4G7TrWc2WD875CqRWZ/bh3e
2nJ38tyzBjKspPjiPsxdbpJVv8t1/mvNiOQqOih28Ij0yMQSgv8LJ7goZp4Zku0v
Uc8QZQ4HnsO5fZt+niG+ovETZW/NcHVYF7WFtJ8GJHPyd/2x7+7GKyQmKhEIAcET
k3FBCodVBnjzBqH3yCcDzhiOyje/LIzVsI1FwBREuGEDn5HUXZyN7Gz03y62wKR/
Fjbg1jMtjbVc8TGbGEnAnfOrYK4Hi046lrUE+iWZ45azPOvWrYRwxZ/W+Wu9lRlm
/PicKe1ocwTGbAbiIWNIUn4khE6RBdP6r3UoytKooPoKEbq7JqlhRU4cyjpOdxBH
4u/VDFCoIooPsW7UUjGwqhEm0Xfoz9lbNl8winbWkHXazftaf/WwB4pFhdTCZCeF
v4pCxpvnbuj9QHyu8FucpzM4cyFWRlEyJjJGHVXFGaEXJnVwvg2oMgKt5Y2c0Gd/
EkIa08pCrzvINugh9N76cN+j4WMzFU4PL843yC34MzcLseofyg/qvC9JPDclvqlE
1KGG57knZpe6OlxDn/+D9iq4Ec2UpR89m38hi14hVbdS6W3OZtxcVZvq34EbWPL/
LuJjU95x1ms7BdFTOrqRHqmunIrsGGk5O6LjRBBGRRcDcgqJUWr6vdgT448F67u0
6zo63KFCTS+nuwJO4rHvQfwRZxgs2DCMuQvXyWKop4602brSrWbLw+ujh21fEC3c
VCpEp7Hts2xDLXnTwSCzzyLkMdgSAQy0uUez5kzBcXiZKm2pKziEBPo3JQEeDwmL
f7pWwhE9RYpJMriu0W3rIsEh1ZX8zAje4gbVMv5Rn0Z3DA8qRgNlvsklDc8NLpbO
2zJSP4YvFqBNPxU6Ppf1Y+IirLBXLybgsoHaehuU63OqqJJLBvJSCC8Zhb7hqk2E
Hp1YtSpcrsNMzzOX5jlzr54v83eqZo4j+HGDpFnzQWgnZFqRcian01uZQ4gB4Lcg
4I2bbdfkGWzq6CAJ4xCNSk2tk4lkAUKjMIGKg6RngIzGEUE+yyv4ap4PEJ5yu2VB
TewVI1s9yRCDpL89WW3YjAfK/MzN63kiCacnuO5pujjoM5iSUZ/AdGF8/unEqBGp
vnyc5CE2DgQ9lYhC2DZ6oDNZ2Hic7Os9EvtqNIu7lFpIGEAG3kofuG+esUSXjNwq
kDUtU6l5xZyYwhjiRtuzJ+QAoJ3AN1Ci1AQnYD08rP2ha41C5q5BcwiN0TnILGge
K6sZQ1TT3D9feBq9KpH8Mi9B6VkcZpZ2asRXFpWLagWqvjsoYpQQF4qRpqC9D0A1
gO5pjA/+nHcgtrupU2yQ/HW1ldXETnQxuyDR9Fn9AGFmdzqmuACvFXkjPfFIl661
myOZebLpUDxsthJaf+YWR2YXGelFy2GKs38CHH+5kzswh+yHGgQuokxH7194x5GI
2tnhm7KaY9TkpnP9Aynk+WbmtSino9P8IlXeKnGyJwePiMmlgYd+ImOSyofpiWgw
M80Vo0IdnysCF3dCBQUy/R3kX+JVSeJDobafdyL8SI2SjQbN+5h2hlVMilos3Yf5
wIu+PeXgcEAhQa9BMGv5Yi/IYONQ4OokG4qlUI2+YIGo9+suyJH8aQEq3ly2ItYk
sZc2QNQ7fImCw0HDnyBEKFoGCUs7P3q9K89S4TzYvsTTjBMYEX+dz9eUp9fcTnBQ
eAx3n6NfbA2qMT4Uw6bUuecg/5ctMVO/zZQ5jDhe2hnmome9YEovdg/bSiuR1fiO
OUTUfzp1JpSmXhL9Q93ImSpQeYeNJj0t4BMSNR0Jknv21pFzbuOvHHE3zBMYxIv0
mTyMo+O7l8HfAR1atnxgPQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4jTxo/x7Z0vt/3q6nbXxW1kfZ7vBm/VbjGfSuGgSMvr/B5BCUjsFNQOi68tzE4Yq
5kij8XO1plPVyqYcnpgZTHObkij0+m7QN93nAD/ZmhD0DUVnWSCesAhIKveF4b7q
Z6AcIhYLwJ1RkR1e7AwtRTJCVgcSKEZUOS+VPS2WFs9ea2nrlNeWnB//hTbQXUkJ
gFH/fjTOWhhmPjov6FQEDNEozNBrSqpqAR0JWcucNhnQNi8mtSN5LBkJzSel24Fj
XgZYqE+2gIC5C6PESkkqo/++OkMl6JdncnGX1Yh+J6uOQB3GfZ7AgjIp4izPPkCQ
nWzMOIPMgS2d5/VFtPrkXXULo3FrUhemXXvIlaBhr9Gt59PtvpbuD+MpzDT/uIFt
3D9r8Ay3wU+Mj6hhGAVaR8Ijh5lXs4UYkYnZAsF/cwTBlLvCALUn+W81HiSmOjeb
qKXIh+PJ6cC9X1YN+heNXfi43Ke9C9xXEGdvgHsKC1hGk0FcmVFAYSvRd7xKm05b
o78k88KXyHs6lra304tY0nVr20LWCCgEf9rCmg9msOScx/RRQTxtKBWb/7HXF7+P
wYqZLUe39taGV9djHL5iFx20N1xovh8HBpN1YH39kaiQAB6o+VLnyso9nGDmPhLp
cMLD1sYQfzS96irTuvAxd2hsuOc+Yf1pUWVNPX5/toYMSyERuNa+WBQiFGTGeEOr
Nu0L0BIz3IAl8WlUzcR7D5SkxYurseNa3Lv/S9N0j1bYjknm+r7pCWx38/I0bjcw
i34pBVyV3dL8wwNblyDosvHxV9NxmSukjPU5ceXOfaPuXmC2fm+1bDW8hS2ztksw
0z+e+ZatHo0DDxDwp6PnzLqjtnQhcwO9GqOZjRkwnLyZxrAEsmU7pZ8ljyzcnbeQ
iI+4iDWVnKRimfwkf4mW9zi0FEZX+9L9aKR1kroD6U9n0tgFl9+UuCDEavk47PUd
6IR8HEUpiitCU8LDT5WQx8ZFUe72vTX3YdHLXOJNRWgoBzylUnqJX68s/SJptnon
52qiZ9nR/pMDR5DM+JarWVn2RC3+lBSFwXywiGlH0QEGMuowgV+Bs1FT74Q6DElp
Kkbds0JcaUZsxHV0lVvyjLmtXKUEXPIWMXN+dnEBlosjWLegGOpiHq0fzhEu7src
VHqQ4G7gT1FfcRf7nZpQD0RbuflLC7Flg36+NC3KlXLO1TBIEBZCcfjp80NWhZFQ
Ad62IwVbtZCnR01Q/hML1sniyNCrZimd1A9Gpzy9obJM7a5T7pIk9foE+pqqnzUi
ySy7bdPcOfMBNFgwKt2wvPZEofULlH6njGxbkf/vCM1cfrN4Nk/d3IGhoh0Wvxbh
gI26npqDHG1jJrCTPgjiFnjHe1a9aBnjMawsqzOsXL8=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nN47jJWcHNPNmuE3diEKsKddTBl3CvQJj709DSXN+KbQIORd5oBy7EgAM/SzUqCA
lKM8dePclSXhEK63wCBTkmKIIhSXsJMXJGH3dFll3kNwOyt/xBK/m8ZKyNGJ6U4t
bZGknYD+bYvIXbylKshODImsalzPubYiFL8N2iyLYUc/bBTaioopoReRfVyQw6h0
z6syPm8BMHDXAgVHfm+xAnK8QPqJnq/if0jhAWE9qyER7sMy1X+M/mMjmYia7yN3
r+1G7hpIm8DUO4XmpGS/3Enh8dWz6p3NdpvLJfcVBnpciPNs1Kh3BSxXPjZAF/Rt
3U2BD2vT+5T53sG58E9dZZF0Lkn8abiPsB7umZX9HkUsGghD/MMz5eFuCKpoL49S
M0vfWQWBkLPEqjPY90AFiAzF6v2paTFWSSnm/FKRPvSY6qJPUKoEAY8NnuM1afrx
OQNNTakKwEFS6QY6yYTrC0NQZRgjlyiF7xuFk1kFVjHi5TWM3LpHCa2dQdkCYQq3
EdD0s7jsUncKQe/xxuKj5h4DNawDlnvjYgeEGmz3EjXUZ0fox7xw4O1yudHV5zIX
ydlz3OHSVgypl5gBz5RP936H3ujsNZbqg1hWpH9O+BG6HqkO6/cbfY9utoBTHLBD
It6GnsWhrHALImtKASqWmbR0kYgduP5PbturLe+kdaYD/siCvhtP+kaPN5AxEM4n
R4qwx1fTxFPdn7g3C4sbE/TohyJGLOG8cCIXl0bVKpcVGFPkvatiYcUSDPQDoRB+
2voBu7VUEJNlLAMVjZIrmCZo8iqpyPREHyrjt+n/23dh/6Jba+9QGbaMg162mgXP
ER4wMTWED4q016hpUdQf2E2QyoByzi7vx8KJ6mArDsAQgTYpfEGx29CFfFhIUuZN
MwjuIduuXl5CS6mrQ+cF4cRsWh83NTHZXY0wvkIkSQ6ucbDMNdRyKDd1gyl5exdl
PCfzWsVRbpZbjFaTSW9HXRnk07eVpLCfxYAtd9vx3loZLSQ48MpwNhKwoeL6O+2S
VHO4SjhBr2U0qkIGZF9Qoag9/oG3yYjYaGu0IBcshzlj97h1I6SD3EIQ8wpEXyy5
LqVwAI3Gb71q49oQcBBtzW0/Axp88Qo43F3loXdt/kJmk+GLKcmfuGqvaghbhcfW
JyJmpuHzvVANPq5D2hp0VfP+0KRonQBIIYARxnauyfxRKm1Idhz3G4zqevK1EZqa
LrRJp/lPfhsVqJV8yEI38eFtFHNQQkOJjJkWAX7nJU7Wat5CQsCHnmH9Pg77Rvny
VTAfGRz1Y7GH6nTgDCRranJuk5ZKH33SA/8aiVQtr7sxBw2tRK/7hZOestjT/4jf
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wO7xOZLIcw8QmBQVmpx3x19TOqhMOsePRoL8iGdP+GzxZ1t5fPaOaHmlFIgy38y9
u2j6kB+IitrwNABV6jWDT7S51dSZQV6qYCKbTpilUJr1Qsk1SJ9fkkrpV4HxYShu
uxYZuLFXPf7iHWtvSb5gSauz/U3IiDsOjOaM2lx8xCbWKCTvPzZ+Fdbfld2Y7tPo
wP2atIDFpLpiE8v4d/a3ekx6kYZWEiQ6XfgMawnwaB+F4gReFB6lvAPS7GpsAKYS
lUNbsq9cLcd0X0oc40D7QUoCU9bU+N7v9YuvJrM6VvXorI+781WubAB+vxeH8Zz2
MdpQbjpJ5Ep1xZ+5DY+MJCHoshihjsMUOI2kK1eZRUFw9Ijy3WEqKFG6BCs6lQ+3
`protect END_PROTECTED

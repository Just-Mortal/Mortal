`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZt++c9SIs+hGcCpqOKMkbfhZ9LX2nW4BJ87Gcw+UNiZsp+RfTFiRK+rzfzkUUwo
dy1qTMysCgHw45NnkUDJ9YS+QgUCtKKAAi1OdtApidR8HuSg8kgrfV31uGmYEF8w
x3yCoRosFPh3Hs+aXYHl3LrzvERAvMGukZBSKXKexKFwH6z8jabUsgjZCKqfjNjw
Z3JkcoeOrSyHBzQGVmHVxxND7k1n+Xx5MDT+XOwLotH9WfHd6mVoU7coSHqRqWUM
9UOI2huqsFhOQmMuLaVyaD1wiNIKCwb9JRtDv1SzOE/bZHmuQtd1NguvCjUNFQn+
mVYGm/5jg4ujTlYcoDKDStANsweG3nQyDoXZMq86JStscRwfNkxqfkNiDsSLdzvn
aEdk2hblN2emTrYckcih+F2yc8cLhdQRt9INNHwuim27mZjn0ZS4QRLV4t9AluCn
zi2QPldpfsadErM9QATIV3PU0HK4PArTIVswtoegwDwJzxvWPtH+F02QtPmfjc/2
5a7G7DWSbXgv/bVMA65LIpyMlnXb06kUzlZgKR/9Atdyqs4nNmDBtb3Y0Re5e6rY
nZArsrlR3nmJJjxWvn4kj+twsN3h2PoqlL2gOKA1ibQYKL9I54sGuOG8K+Jgaywe
Krhv23o018iJC6eII5qkzCppIuysFLydWkNmI9fN+pUylOVk6sR4NGCJ2yCGGCAj
UJ61vWGsryDDHGw5RMjZuRjERGMz/9uXE4n3K/UY5khL15MW3Mx5Ev8YI8+pz23R
BP5QO7ywz8ivrlB8DoweFCDerhc9PY5ghvL4ctwEEXzHgWDutI3yTRnqC9CBzI7L
1D3ydpGu11Fl87R0EqkqAjTqxfRtqB4ROGFfD5QbDV0oEVWJumEqzhiRUt5ck2LU
e3PU6phcplhqNo3ZBuXYKGmQYbj8GpAH+/mYWHJ6WuUQ57uSAA5AYZQq+HWNRxmn
an58oB/qF5I1+O/PucWsGFGGDnwFe35rJgFUkq7aek33nI9bLDpPq4rKClhjGvms
6J9kl/Aom8ps5Qm9HKOksGYUEckyJaBeYGznYRjAU3pH5aD33fz5kKy2Rq8LSN8r
iGJzV0bSyHiHtVhP3FJLMTo0bFl55x9GMhd2vqQ4ZV9kWgyrBSPhz2qOnU0Hz+ld
aFjDRmqDKfW4J37zxpZQIEf3Rlk6pw66L4OS7+k7wn7ClyMBD+iVQPR076h1LLwB
uWUK+OOdwfHCFZ5SrpAgHvbjTBJ/Nw1VcS6l5BBovQysJKK8NsMpLko5mqsyLzER
l2jQR3BIuJ//npeAbnN1a39JuDPojyKmEdEVKUZIjfZxbHOsM3SDP09lJLHKG0/D
ryg78jdxzDh5Ie8SPIBBUhkosDAdW/FTdetYh4uifTdnmPcKDSSkEzcyoj5Yf0QE
jnpJETdZP8hE5lHVxlf2mHHTabQhVrHq0vOCTuQ6igd8qMfKO+2DSwiwQHnt3i8c
fEk29GBQm9foTi0Ibp6Wwhj0IrsqdjN8DFOTP1h9uLy43eKCI/8amIxfnQhH3R5F
+3Y5ixdzGnEsPBkU2/lIkJ8FNW4VtZbwKxxO3+wTLf5DuCD7WmvO84VrlxvMSPQZ
g7Y/wYtFn5sexYZBSsbFaspELoPkOHgQMeM16QFd6fR2589stxd2CAx3uzGH792H
sjIsbh6kLWAat4xLxtjJSOjqa8+Is4SclgN4GJ9CjHbXi6LJFAQCPzfkWXy44Zil
JS5uGQ9picUvf1L+BSFGOid5mBAJsN9mlYNs+oovOuz05otManPATKXgTKHWQJTn
bqnEaNeF6r7QOIalQ4j10XKa8HkfehTSWBkjlpM9GtXPsWuVEcoxTW9WzizQVyhA
Byv3jS/+qPcTdozvnulLGuD6r2asEOVJYkzZmgDfvDDoABwTGdHj1/d9CxeIznOC
+awSzmDLmg6fb8bD0JtNhir2vBc5xrM7vQJw+h2zsxi3GOfMh19Ru5kLX8dJ+fxo
wSdygPk7FIBqBgIKG3/ifhuEnm5J3raUb1X+9FyA4dv1eFozLyYZO69YFxAWH4t3
Z6JWJmy+sQs/09TCZyMyjfrx71AHHa2ITKoFWVPgCSkI0luzK+pdgDXQhvsa+m6r
KjZh117v2UfvNJfPMclkiR399NGn7qyLV35PSNjmyWk=
`protect END_PROTECTED

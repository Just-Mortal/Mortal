`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IsajeXcYsUXRWXXpH9wJobaojsKpNZQwKDs2EJBG4gCV1ylmq0HYcww6qxTaAAsY
qxKAIOVXLPoYy5xt998vlz3oBHHfBnyK3RzsogbKGl5bKVwGEQHig0Z82w0WTVMD
HRo4oOIYCJpemS/ltpUWr+3fFvNWnfmHRBLJ9cQBemcvTSuuJ07TCfXHbpe18u1a
QODz2bnjaTzCYP3jErmJnv8sDb8QsKJIs3nW/RoUAW3o0cL1sYW6XEWe82Jxc+tm
/Wuf/BnBHdoa1N+sUFhfhEbxzLJU2YKG+TUnGEKnPBjGWE7Sa6F//dnLgXk2PAnd
HT9RZArGwPTuLrm0w1Q5GhOiXtJbzfBWbZ6mqaWr4YYBBPS2NbFlfIBHTWIkDtjW
toEyaDBFEFj4k6GWwafi6fdME0TvxF/488MFVOxXzBsKb7FbjgL4+xEmJ+z3ahnK
DUyran5iClBXQJXjhrL95M2LeRlDQV50PRRJ34YtAHFZrXmvu5HE1IwPHaAKpzus
ppXJR/4PZdV2FdyyR1H+qjXBISiWHvSt56tKA0i/lzSu9MzkDhjn0Vj04Z0h7Fb+
262RP+9xMnZk+VGvf7qenq0AnVtwWSiT04rtlHNhwT+PrF8879T3mFUv15xo/LcD
qQVqX+8WKGLmf/sBfv+aY+8HkEDAlfJC2hQr2CGlgLxZgZbWUy8IJ3CtgcBxDLl0
DL5l/I2Dj7GQkWoey+apwfgZ1uLFSS4feM+3VU7hD5tlz3CVIyYZMDxHXz5Z+a4J
cU02kPEVfyUG7ntipW/8pVnMuVwdjaPA1HGXknQLPafzvf841CY1N5p6KKlfxBOW
kz7TnHcZ2+WZWN7ADTsCoHTzbhqtfFzOXsjzJBnZ597d52+dtYLNYUVApvPOGS6B
0czmUWkx1RQHQbEQ5pC8fkwU6uxfGDQemgre+6tmguUTCWjjf+iDFuwEAQ8kqFSI
Mq+EwYbrqK/BGlpXQetRKcP4EiE8F7SEwDC3q/8e9Rnfm84pZZM9+z2x7DL8KRfT
U2HIXiqroFa9YQgF81Dx33u48t+AMSM0Pw3GItW/6/Lx1YpQxxq8Aqo8SUnVqxBK
kQGpE1C7l0vHnoIGdyGrI8yFbTZy93drYmrnEdKJLiazYZgbEcqdRAWtk+RBs9OY
q2+k7cKzITnWwg5Py3Q+fQd60xH3ysiHLaSAhYI/VVn/xeHMpR9wM/TlHs/P9wTT
P0OoG0DHyiEjv/bGU9fiB8ezRIFv5UZ7wU4tE04UwSt2nOwrRdgJ2sau/crcMixK
mRpCahAdf5KWnq3GgRvBMB3rrsLIFXGkooIUVNxBKdTdHE2hO9EsfGoNhH31JDDf
dpdYaqIgZSIpQIUigU4jbINxmYKAa6oNLxmIvZW6HxUtdZf+tWctB3m2v6BoKare
iKtsUYIRgNxNWwfhPP1OPIzKPA75DQLCpMr5jDrgNBMWwqcws1BKEPu2hizyvA9j
0779jPZJhPKgIcKAoFOkpX0bLt+HkdgFc4I9Zj8IIYHxw2t1HTBOG/q6U5e+lp3E
lcbUbTlXivi+kU3szr2z+dSjmmA2Des94TDWobU1D4jlViKXF572HOo31vH+CJIC
nRDe07rw5BnQuISJCaUu9bpwWbp9XP0MZw6obTIU5dhL6BJgR+rhb+rtenVOV2FE
xmkyOlDI+X9jMcKoh+4tDtQscpGml4vzgqlwLjUyqABJYiifMxvDTDzJtBPQheUk
a+T87RECDoTQ4dBUabOyeRDG05uqiDblBzn0MJ+ne68lSwVC4shLKWfiS3knFZUs
DMBQlYYz1fD3VUbyY+PdYlPGeMX0oOxp6tJD/tcRzn1KPJBFgTmmIMqhEMUO++tq
ucdgPmpVAMIXrDsvvQh+JjueXiP+L7o7Ge8cwDBmuiL2lwoZOmlKPS0mY2DkE3GQ
uKe45LwcQyeFvyFDXCx/pZAgwLsKkeUCJA33WR3IdusD94HTOdQL8BDru6dqdRdB
dpT49PU+fTOSquaJkUZehJ+IN3MiVU+n+6NE/kdDupssoHn+zShgQJBtcijrD93W
+OLfkJ9h93Lv+9AC5MEEWbrXDkJRBLRIkJgcK0WDrjB5YnbJG0uw/dB7NNCHcQth
HD5+tepXCtMpYnCztW2fu5P+eGFDCs0LRh/0DA0u8asAQvkTA19zo2wzEHVTQtqV
Zh1nJ3loYml4V2fcpPZBcip7vip/z+lwRmiOWRJ9ibreGbu+G4GwXSj2sUJ8U1RG
o1GnyboAufoGBil0KHRml8rWFRfWJFd3InQI6/jKQPrpdhz9c2ibyHHJ0kVZvoHZ
s4+Bm5wC2/hDbj93V10RzyTgA4Sys8qi8fGanlXqj2jHFBMp3Y7KDVqLgI5OeYag
T7IiaYgf5rRJIECFm66uf/pdJtj5tBrYcH6/o7GmFrf/rZZTKZN0MynpnFeQhjh9
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rn5OfWdWAO8sjtFbo2v2XV/wB9ueYsjjO6plqcJ5A/eqanusCpVxqyZkoBqiVZCy
zgQ8L/TPP0Ud7/01Z03fMa7ayWqiLXO+cUqPMcllBigSdPxoExGWVZLLIuz1IZvN
wfdQDSz8JiKw/bxoADt8vaxruXhN79GpwO0mQkPfjqz6rFWBHJOHdsu7BkSSLPJW
lpDLKf7dsYR7sBzPk/yzBl//Kv98qAiDVI2qTYv7NnRRK9Xy+v6yCUaAQSu1SDrb
10jzQmJV3VvsjHpXjTEzQj7RoLom3pcHWZUHXjtWlmt4yq/XDqV8RQvHYcldhdV9
UWZG48wU3xtCJOlNAm7aIqUtxnM2GOrkVlPhZ66qFuuPzGi0g9VaGvFZe2fDLDnG
IfelR1f88r+pFJFlJCFFI7eXUW1Ae8dwAjlEqXEQWKYKRLoOcw9F3imnR1cCI9MT
4oMMCDUYjKzzpMuniU3x+/DMDA4fZd5Af4p3Bbt9COCqA9AdB0vPxABzbTaPr9OV
7QDn5s83vShxtrECDzs0RRJEz6vN+uHm/5CRnDb6c3QUujVOs3d4TsjyKBuLJ0An
UyVxAQI+2Rai+W3t06WdQnd5Y+mnpiUgsPOF3jxprfg=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+GBaD5EGqdTNlCD1CeXdWoHs/XZhNacJwEQ0r016tgpep8Q9a2j0JMbu75p7mEz
IhCTC/+Y5hikhI4k1Ifl4Z9EeBOkUF6VV4HGW/1z3+YbF9tbutnfw8ISxPfzgnF6
73JtRiHbKo5gJf/vNiUVKuFuySJvfDeE3C6UI/xZR49Hk+WHzOz2jXO3PxOXHyaD
UFa3lZXAXQNjrySYowJXwhXqNYwKN4yhV8znX1nSDm8Rw7VG094SvS+7nhK9poT7
DvoObAqY/ZNDtmQWtAWQid/N0bQtkbzOsgBzjQdG4ITnRwYDkYXHbwB/HBbNVuLM
jo3dDio3QywV3xENFUwCgEiIb4+DPLfzGUTOgEVT3CVst37KvHaCbz051ilpNotd
YIlVcxTgdCmeLG4f97OwCSsOue7gv6Cj6Efhp5rNGWKpQxFB79kEuOuTceCUt1bn
EoKo47Un34J9oUE1/yQpzyl2ehRr8Jg9uS0sqcil6alVNZx9JRxbKhQBsjgOsU09
qcDD1c3DKr02uVxz5gMm/heSUxLC7Zu7lc6RL5LdbkU=
`protect END_PROTECTED

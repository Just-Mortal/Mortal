`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2C7p8biYB8S95NS2/uYOTHFdh28zLKuNhCZwVPoQ3EOCGFn+eBNg68h+xwG6XJa
A4vuZxNqeWPy8Fiw3ZLFQw6t0FRGB6JO/L8sLzP6MuE2uj6pyclMIB+lCwGImHxo
pkdqW9R9A5iTwYKb045EeKvWNU0zKggXJDeo9NaTlWH3jjwvzyYpLtdDVfqczKNh
xguge4fO2dig5T0CiDCvzDK+/AL8Vc+z8/Wlqz1iH4kdM+WrumkfGaOV/XWU5fuq
40qUWb4aopAHFsGIkl0lDUMD4vG55emFCx/SekVtDRghK8MWUh1meaLnw/P6kuGB
S+CuzkgUOT3SwiKHzOuxWAtMnFr8nWNVv8/uyjRuP1qfLcocs03vEl2iParK80iv
nAr/hefF+9HXNj0qHADUFmpG1vZsWdmAxEMgbvQN5JnQXYlYtabaFhvr09x/9J8Z
/ikQhsxooZSCc0OPg+iDejI1+cgNhUcz+UWZshS+tU7OhT5mUQLGUuHzsy8RI6Nb
pQQxHZJoZjVOSw67KhZ2ByCnIZJcPrbjXjqmm1DPCQ9W3AfI7O0RLRx5VvFxCii3
fWAZfF9y/gtOG5q038Qnvtd7IIWY/YznrRX0d/0bf15XRhWdIS8xjWpsQj7oSTZA
97cYW/60v/ZFXaguvrdCRW1MhkvOsBuMoW4ZYXpqEZioHfVKi+c/54cQvFZuFlNm
mFElZSoOthbClZqmCQg+WNH/cByuuhWQP0CXOXEFtZgiWg+csthNxtKFqN6V+a5t
T64upLpUHQsdPMyIEX3d3pjmmhE1fOGP8uxmyzEovIT0BBKvzsy4c7Ft1BN7h3cs
+AVzZML7qt/hizaybV5e00AoNXUG5CZd0pRUuHEmEA8=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aEJZzUmPrQ8grSRecJvwoJTVr640de1Pfw8Go2Qt18AqvX/3RBZN+bXOruTqi4Tc
f1ODGgIvmyo5vvun/lZVWTAKI72RHQbTWRdMCaR0mpcPKANn/hHkAMdqg1oQcaqc
qUGPX0WRa8RR/c4E8vu7kqmUuMDmdcrv3ERoy4OCYB7ENNZ166RcQ5hZ0iaR8Xca
p9+5OsmJ4ESEvZvXyBRglw+gDkL01swxWDuk3NI3xHff2UdhUMLNLqNoms/sNXuu
joLeFcW+59hSdgsetOTKkpWbaeVesEGNRPfTgPHXy32F6sHXuKXG2ziPgNMD+tLR
arW9EazSZiSHxXruJxlhNb1Kimk6uONpgXhGR3mC39Zn3LgsSKCrr33o3zdntjCu
u6BLoSctAX9oh8jKZGjxEUFSYsCf2hqC0flz0zINSgnECRk3IUPE21NTRuRtCFxq
hhXucMzfunc4M/f2T6xr+Bgd3AZobzac0z0RZfpZkm0EJFA1qmbqlCyJDf1d8YnB
JVnoIuL9zx4qChkMhhHuuugrQrZp7IixIcq5tplHRf6A8LHJrxRfhppySgMp911I
V8hR38d1Se3k6Vk+FCm5ocbmr/fEWhaDXhU9z3hlcq5DQnU+/afuuQEUQjTvGjJe
c+WHfljqIwbDy+7pVJJm4zsOQs1j+86wX4vwMyY0vT7Hm+0nWH24Gk/DGuQkuTS6
KlVg/d900iUSgh5sepQIimm9FMZja01EK9XvWcFPqHdfDPwi22e2EwYZp6U0mdSL
tkfYqYA/f8Q+dZg+6dlw2hxseUUpecuiiClm2uCPQvGJYafkB8TqUyoSbvwOsbiA
sPDoKRtvVPqKU6OTbm0WYiC4ec3IUmmGrYiIhAv+xgrsS+khQJYutuWb9WCau+kP
pyWRVBYWHtH/teu7hVgpHnCvD8q3Tg+wLTfgRlG/vlygTL7DT3G5TApvh655KEU7
D8PaOfIl9hkAIQDjIy4rZlix5jU8goTWKTwOQ20Smup6Df8C4BQ63kAN0xqVamcN
VeK4Ha79XXdz2/rQk2OOBMvgtOiLqQmg+spepVTfkeTMBR2qeJtmY+UNg0Ld4GZt
QRpp+4HgLGH8ivUMBYlJnQ5x4vN7FQyw2C5CYnT+lYqnWY3UK6cRCugFVWhuuBIv
icvnFKQz8mWoEZiC2eufg87tDiytK0t6T5E4Qj36185zF/M0byQ/nDvvyxIuyOxN
ULz14BehkFyUK37Gwf4Qm9pMThXwV525a7lHVe6qF3o=
`protect END_PROTECTED

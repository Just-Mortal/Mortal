`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WA7Z+/7Tg8TunrzYOP6uUhwxRMuZeIBh4QKqadWBLszstO0/cvOd8LaA/0VNpmON
QJXJVKKooTvrWbh+lQh9yaEJwUCsEBre5TxlhSBZ1jE9JMCns1JPo9H+eQZheSZc
6u2sEQzASby+uodjnbzxbOAjwJHAQ5B7VitNF/XU92DiEUfEOdt7WWCd0j91w8WJ
2n9yUcsMcOYIUyfmnODLBReoUgIut/WHMWDQ0w+IM+C0qxzfQa2TcyUUT5hEr8A4
ZSa29TB8UJVx0unfVgVBNJdqEOFhr4nJON1h+9DK2bFkaz70JKa7kmJIWyl1OsUl
pMxxLze7xfwuiDLMhtOH1h0+SE2WK4l1xSNFxWmrAQ81/LpFH6lpf1z6fn9n3sjM
2XGPY8QuF5G1QtSnLFvdaw==
`protect END_PROTECTED

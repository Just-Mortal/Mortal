`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XxZfkoxTZG19T21/7MTxoF2vpmeIVnGIf3FwitLig73qNOwSAkswPHTfm68mFNUE
d7XAGDxHx4R3Us4mmYuYEfZrxpyi26JqsTDLiSvcGwiG+p3LUtwgmFK6nIpexaG4
6UYXtBzlZ1jXNwcwPPjplA2QwRnGnaVJLTZr449mJ8ogyEYE/NQ/QXGYMS+xagoj
NDcrr1QSLffppcPV9Dfu05pdkZtwfNny6BK+RrHQfBlMehonijerVUD/0JcVn6pk
vaUW3o+rcfoEpx9GxMN473a0RRmWoXk0j3kR88FAdTtVfADpxpidhLU3cVmztw7I
fXY/oLEzyRjSu1CbwouYKkvjzh/u+OeoDxlnbo1MYNTrwJt5rkT/MekqbYPvbz/n
91knnKb8+AA0AwR+LermKoQAY/FYVQBn76MB8jXgy46z8b6Ird1ieRaapMdLvhZz
Vn/2xiGL8m+YDXRHrbPC4eMkPupJPFjHHIPCGaD/za/vHH2mGzm9zeZ2+Oqv7dCA
mY4LyTM6l7Q108IlnaMY44bTRpXkWMI5Nt/VinPWIS5aJeyz/6mydUFy1rWGycjv
ILAAM3kTCL47FGRuzXFpgIm7MWx4NTZDmMOGHo6Q8pXmMskp96CPNozZ/bYavLSM
nbEoED/6HseNannbcEt4EQaEV6o7Ok2oXluulxeq0AD0dsMuS74VXYWpB24ksXHG
qlBp4HlW/qpXQatV8G/UmVXZz1GF+s+3LUxz0HXgo/X9WadrXXjlLd7+TacQHJB8
GAT8c7RDJC4+sbFe/vpLt0kyYNtq4WmjgjRo0vJI72dtl6HZ4sIKzeCrF+pmjvSm
RlsSFQmEP04Wr4QqkktDZ5+8ad3wPZiqYElT7rodo2rFM4W4ujTiP7XvyF7UZbFd
aPe1m8e5io+gP+/d8/cIVbJk9Ci8K14m7ZCQpMjImXGeoOKZI9+T5SY61BCvoWyo
RBwJtlNj3vcMQLJBEjdq9GtuzJxX7+UpBpwsoqiQLpXzMKidHwLg2N1pw59yx1e0
+JueHqANI8oDH0kJNDU4Yn9zuKuuKKlLwwjF/BUXuZ3zIVAK46T3NI/Uc2LxmngV
JQbVci5Y+9hNsnYgZJQpDbOwrycTLrL+aO7jrYS2PFAAWsfCbs/hdyRJT970mNwO
46yYL01U9vHzxO8lmm8zJ/uv8w2tebM+x1/o15AqZhqH9iypn1FgTupgDuQlby0S
B6B+6sz69sgc05PIz9pE/KuP6E+T7qVqYXsUu/BOV4U34Aaa+3GcCijvvZGZj/S0
dOIGZedaxQgnCCWM7uDUY15+gO1pI/Iz9ptqpy5oFB4=
`protect END_PROTECTED

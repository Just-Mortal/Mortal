`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJPOlQLbSYE7Y6XStQCy6DWKFKhm+Tt+awn+0fm3XcU+UznI60Ml/HIpl+nDZtQC
sMjslpTIYaFlR9yONAVRUB/VPT0S3bK24sCfwm0wkDg/M1TjSc6H3NmjsHNd9V3t
/nuGOrYRy3NEPX6Yw9qgqzRpo/V81LmRjUqpBWwzKEHRRsUkFTN3m9bOT6v7snpt
Tc2CPiELZJ9MCs63ahe/7prynwUzD39S5ER1iDnlhwyvD8XesxWy3dwvNyuZFbtW
BYwbvx4ArWx2gyEWC4gkQ69ZOOzFDICDM6agvmPyizUolIVCYsPjRv5ECfz0FLKS
UT3FLjq4+kUThjJQLBY/1W6Y/qEqFFrvNcWP/VpuJ76QZmizgqcZGB2gycfzTfXD
QGMbJkrM+dcYbqz3uE5J2sKmlvlL7fC5eBc/YNP6A80vGTVOWwtrSKlpDoyZXoSN
6CD+B1UbGEeSrgmM0i4hzQ8XJekKjerjEvaFZwKpHFj7LS9bO9M/+0R8VB5xs1gC
ETU7opMUgN/JAsXfRfiJakvSMFp+aSn2LBWngaQiHGk/XseUg/n01dp7BNr5PSi+
s2BTSzhkvYSEerJg3kL6nofUneye+Avh0UvunAfc7ujgkwZen8EqOHD1NjqGc7Rl
QZDQpMn51qjCk5CI2ah5Q06mYvGKwERWe5j7ECqBZkltzsJaQTYXfFofIaAN9SNI
m5+jmjgnzuSKQKBDzepvBbFRBsY2lqvG3ZTjkjyXfI+U0RrNaitoAPrCb7kHneEg
s4/nvdPkoqpvP3ikZXSy5GhZFOxzod5P1etP9N+NYPUJH9uskcry093DHpA2mFC/
Oj/BQBO1lJzG7roZU3Smbf+OtIAf2i+1wRHFESxY4aM=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
feHcJ6dA+dxB4mcBTqJY1VwDn6ZjKo/J90uiaOhPCZpaKqOndNHaDBFJhV/2ZSfg
fzN8ZQABJiz2iNyH68X1kUI8l43534bwqAQWXGgelPYURi+nJQCD6YIu+wQM36Ra
YZoElnfV1pgGvhUOLg81UZ9iBnhRiLRJowoQMSvoftGXmAi60s1PxM0sBLqxu7oT
XQ60KWRvy2VH0A+rTs8nRdCVWOiHycxbdRlHCgr7gQOlp3jlWu65kVN/A2hSIoED
JK2GA+ohOnogIruKW0dxy0TRdLoOv9pQoxJAdjT+ax/gB5HGycIQ+za/CL8JGrWf
1VdtdCW3dXLR0/PTG5deRL9kGIfzHrgPY506pnZGg4cSQ38QQKM3ODZOszaVq+vl
2WXnnShuoDIhcrrq7frSTv88uA6nkb2+xl7OmX0lPOFy7o4IumcZ6Hlyo4wIBoS6
NKFtbcN/Jethm4NtpkSoWsI/6xnla47dAjoCN48GFAvBMtRoTXnNSfHXET5M08xV
0xH68ygVWh1PCHadGn4uP9PjRgL9kj5qupgJEJCOawzKj8AGylXfuvG9tsV+zRJe
uIc366oV6XF6mxtivWSa2xSRUiQOFx78E/gyIA5z+5cUFN1dcWH+WULTfJGYT6wT
mfYdXB6WRDkdZho6TGJvBigExhckAcp1uKEsx5HHWUCJkjnUA62xOq7XSNS3JFo+
tx08gEpuPMXM7EewbcnwkENsTbC6MSKQEJC6hbEOmaud37N7y/WReU8tviKnjkX8
EqMUQmgHUUmVMcK57S8YFEpDNYrUkdUwsrUCEgqPbYp17MUMHMRfGRGKgEhklIIE
uKuZI1Y9v6pOsW6iT43uos0GCbDqWzNCE188Lnjwc4U/Y5jr9lnooAFIbpAJyfYX
4vCgO4oKc/NpcMCiqbSFCerRKVaFpUtv3rUkmhEV/6Z6so1PnhdGsU9mpu1Iz6H1
65VCyBdvIIuidzq/iBwSsMpGADJXFZc/2+HxJTsgMlw/HzITouyNbBDRvb8znrRf
ipYv6koBK4hm0y7IlumKK2sisfz+F1bdcW8HDKFRS1Lrb1NMC/aoI1F+btAnhT2P
NIrPnyaTcfj5DSuRDxp5miqcOasSliM/DT52EwZkRPONGEbDGvPtckPXcEVU2Q+M
p/s/1wpP/F3By37HCnQkMIpaSOxmdhPb4LoV5fSLD+BIPMpZmqLhU55vf4BFVkpX
vGfsFdD3r3LCHwYuxvgFwRDO0kkMAGwFWJmvR1QnuLrGz/GDVS3XFAwGVuFk5GGz
CLopfc1H3+4k+JNNlw94GJwE/Cwa5Tahecfrjukq2oxpLJPD5BiQL06nJJGx4/ZW
MhMCw9VqgJgo+pX1/a7PiqMkl6p45TdIC73dMIEAgYmke1JP3wmePfNgLJ01vHMv
V851VeunsgaqwjENguHD+3VFElKo0kDaGnU/YJ81eGYLVkBVVBYpW4B6rWyqinEj
SVcDiiKphdNKV8RbxPNFLxCAUGM0ji/3MTSgIN59qQlo0BkxNBxVeq7qENocwaTy
fjqPMOrA9cbKb3mcaUaO5fJAMNWngJ/tBnCjZbv5/khEh6Eyh6CRhDI9npWYNLzx
NjNbuuhVUDy+WuikvaiJ/yIaUnFtzf8K5tvKe5/9wa5yv6juZmYO1t+JR5Mej9hp
P4R/ws3zG2/njBkl3yp+M9U+NRZCkXlE8nyadU1/rCR8eFtI8VLmA0vQhuu73twh
rgb/oXm536RtuB/yGRx+I6HTEip/lpgWfohvEv4HzJKQyxs9QEqjvPDogQcQFctw
YSlh4ziTndjD6JCu8NlYzAGJepkn2jB7UEqXT4yHLYog7frljlUQlqTZZS0/6Q2v
Q+k0WyGjLXkwXk+O3zrZBJl6QRwYlmaoWchfhICGQ58NhApucd3PIE29xlW8Ir0J
MdMBqscyuaq6TOGExaVcHUK8u5THxit0puCLfFFj7Zv9z46QdgSAjQzaY5zn6Ilv
CMFW805KlpVBP3h9fxNYpzU7nFhjCiyyQvgfMs4QTIFsbNnLt7AB+qKbUzFg2sVa
kz2AcB65+AHaFpcPLf43bO0y2zCz3di4bwIvGwA0kG9xwaUFdhcprIsBkJ2xijQi
9bLIT628v6cUjw4iHXsOb0VSELNaLKffIUJmC/vawS3D23vqDcVGBTGmRBDYlQm2
SuFQRvUU8tlimZCx2p7chqkydZfFNjYcAKN3deLax10iKrRGEqEnMuI0Cs5tvgZJ
QM4w4acvRd0Tlk+QvtYtDa6uLaFDd1x2BcA62uKrT7zZQn0IwEAj7T7CmZyifPfX
y6MewXwK8zzpn6Qp9dRr7Xb19atM7CvJfSj2i9PKlCLIBvnrRRnWXfw4lPenIZzm
BXDoXMhMDxyEB5WHEWNus9iZL9/Rs61iDzooavn++72nROqBRq6rq2LaJvOzZtIT
n1A6HvXXeOhKBi9EIQho4Bop6xsChNV8WgEjLCuYDvOLA6etEJj4IyciSFiuizho
gghcEzUFUxDKatpIt6kaky2xLlB5NVMHRBs5x0gS7I/3t8LR2S0IwxnyApHRCGi0
TCh2pvaluSse7jBZjrtLrWTsg/7XOtCcg6PqLKb1Pd7jwRwEalozgy1zdEpJiB+o
Z9V5pzspeg2eRaJalgDmvIhTFOKiKZGvPM7tXYJSkcYm/56m5QjjlZw4c+5p/jUE
EBLbLYXWGhrrQ5+jO7iiQLmtTAZeHG/lPAssIf7QRWtNXM1NaRFbilWY2HqAUDUX
9Th0Vi7M17nDvrlpotulyiU25k5zcQiZkxSfn7LflWan524N/9uOfbTMEStr3yBz
nqAhT135MwaSgQ3wo1E7ikU2Rndcx7RRB/tWElHkmBYkljsNsz72smM4xf1XsDPk
h52RSgWzanfZg8Q7AOwZlrXMJoenHnQNT9E4qRs015gnj4Ot385pIQlRjT1w2NMX
jMVYplIhDVnIABAPLoTVhRz3lSyHo/sKxwaWixBVIUtP/mJg+nqU7gWiR86Qmi8p
+KjG45sDtsRyxvGJ9yZQkRPRDv22EOa9sChSrXnzeTqkFd/RNKNQw5l3wOoUka27
wkfwX7CVBAUE4g9XD+58GGCc9diu+GDjnoflOUtB+EhqKOFCOIo5kpHh8LLZArQA
DSVbHnjcoTMueuXkFnAPnV0fJv5Dr7NNjgsGYq1uP71gYg/WLymz9Oq+ZIGCGiHP
JmTHIzUT0N5vRdod5Wtaq85iAiAN6KK6aqxjM3bWZ87tK3nUH/YuALxmzl1W1C6s
UJmZekaffyQNV1HBq+5amDITOnDnOzkmtPVswv0/Gokq2a9mLRWbw2/NR39Dp2Ts
5Bxi1AAWhaomsRkhQeoEDvtvr95Q7BHSBwrJK/FnwVG0fSljzK20Dx06Zgaq7sLM
UAZIIFwrdhd6CbstOtp8HsK0dkAv5dTpYNiQXVFP3P+r9OS5/i0RWprRkbNoD5JU
vlVdCOtZKk5nTVsQcFdSVkxyc80H3iaWk1Yj1f7quDjn4X29R4M5vxD1kdH84XZi
YGrHfBEhzAlWvE5NqrxSLpSJ3+YB0byuCAzTRCcOTb4OSQ1sB2ajg+6+y2fuajxM
0bx6cfgZV32PV1LRh8xH1hsXGpNlpl+OJlMub4UEbz0NuU592dDSF52K708xG93H
MHyF2lb4NlG2eveJDQ6KR/dX4dAB3tRFq5gG2LfCSltlYP0pVXg2Jm7Ja0l3a+6e
Q56Lqc57RQ27mbBm/RsVOJfv6BZz6BNLe53+DfsYsQdyrj4qmXA55oao+h1d+Im/
CA7/JTbXe0k07AWrIm4+7DrIQK2TFGMop3Fx0VD/SIlOqisweUEa7F3F8ck4lw6M
e1QzNP3BgOwLEY7GTPPy4RtSJFuVE4ji6tsRWClq54djzAXBgNuDd6f4jSNvRq7V
58P3oYEZQfi/vDrRP/iXHrFnCT0v6lIL3vz5E4vTJH6u3nmjp1UT//VXc/Eo3Jdc
IlYsPpBfizRhQC3xR0FI8Jz/dIrAjs+NC0MIoCKV+ym+PeZohmnwtl3kB098bpgQ
WAnFRwlnsfZGZZySCuAQe1sZPwqaYblXP64Ba6IYFUwjanq5qLqriD0kKaN+LeQi
t8YtjLFJBJWYAFdYyHpy+rzC95NHXlzA5+h0yqsZoqDa1W3fMszBIAXMlSKFPF0m
sla4nAJYq+RUE5SCsJ8hncV4M0npMUg1NOEMIRCpv0qbg+y7sWcVuZwAKzNExET6
mRonLoNYQs8UZB0L5FkMtWeyUgFcCjyefhy9f2cb/9wURLcSPJNTvE1ShR4wJQKA
IAKClOyZfOYdcJqW6BpyZOfEs1SKIVW9QT1guqFF2OhUmJ7fyMnDmRHd5yOcEFX5
ACbiF5C2XCqm9wHCe3Sx58f730bkBthJ+u05xGYXC8C2g3a9YRmbdjO5oH76v3s/
0Dy32rYUoxfXirpwJVoDsK/83AwMXy0bJboHuAX5dFin4erdDCfOE5BNiv2OkEhv
HPaWnr11DRsKqkW1pbYGx5wAw3X4T8o/hQCB1ePEdmXpq4jXMJBrTcWaHV5aiKTA
jigziW67B1Eslf/jBKiW4OyiVQYuOyV30dMAFPjyu09+2dnCSjkU9VKqVaKgdc6h
kKvCf5gbQNGL0+YxAQSYoYIGEH4lVq9dFAtOB5ea41vsxY68RlfLZwLZk4pUsTLU
ZzE3y0z81l+7AR5G6/wDag9KfDGmdKfToalhLZl1kgLALiHlYQrz5RIXRsNPTfLP
oYAZbaKbD7erNblQJY5L+kEYdiqZcfRLkLjaTUP6q5TuLfeVgT5TQfaCdPwPJesa
N8cvehU7JPIANYQrbBGvtTCVF2KHvmPbwtMt80e063AMeFm54voTo/EQ6FfXmNi7
YBk2b7D6bhFeo+JvNs2jhD34J6AMxOd2iv5j9NluBfpekKg5SvKRfGMEfRye7nFW
khKynE2pzdYYXIzEZ9/pNSWc/hSNIdfodfpEU6mtVhzZvooEvOqjW7EXQ2hnP174
K4wi6bGmEM3328BFqe32GIDHTSZlvzQNznIcQvotvgy54z9Lmf7WNx6njjHAOUrE
SUvOsFJM2KUz8qDjSuX5c9fksbnKzaQQnL4eH1lQ7Kcth1TVm/anKbHvs01KMivm
Nlw+bs36Y15ESTEmdqjHIHLtAp9/GPunHH6tPZ8GlgJdy7VwhaOky+Wwq4AekY1C
TLMfpueKjynNyrXDqxtiaN3rKg9GFEvueiq+26ymNf9ug/FUTSGH+XmrUJZLXT3F
LST7efr3Kop0a7HT/EkM2YvT/s7TGmE2XDJQpfkjE2ZKcxyM/U3sNt+GadlTLRBO
jU6GEaOsWGVkfTex6OATmpJbXV0XDRM7es2H2c5B8AP5G5cBZ1ji/PNDLN4mRYVg
a+m6sEaZonfhjp8hlOA2X7bQIbBz1lneRw1pJzUPxoVFf89mEoQNAaEj49HvPf2n
RUslevpZTAHA+QHiM5CjRENEyIKqSMaem8Cmd9juouPiuJzfIpcLhkwKBHQ4dNg/
33qdfLc4K6UfU0lySSA+Je7o6/trEyXQ/OoEdH6CkbWimTvDO88r2rP1kOTCe1qL
fmQs2o/4+QspVEQ1rm+tLCHH1q5D9VE/FQ62vmPzqYavrgTrbSECs8nF+z/mAHa/
MeVJadV9y/nOohJobFMEVEMDY/d8AvDIl9WEXvyn+0C/hnqY4Br9XnpO4OsSx6qY
kJ3B+er5dvuCTD1tofOaoCRBfetJzQ8bZMIhHApWwPhQ3DFXpBS6gZqGBfPfSLgg
p0KYY63OfiHo50W5V2gatnddHtNENxefieGoxT7LKpzrqygtTwyxYiCsjRDLd7Yn
GoFmCMHwxsibZsjCsqpQyNyLj1b3pELqDtTAccUDDloNZnne6opmDnAHmHYQTLet
owmpMPrcSOPLVLoyC0TvXIPJyhJ9zNzI5aDwac4RdU4/3YAQpkcpfNARtaWOkjPf
9S9xHUoBqtLsg7VTRe58yNUMoNUjqt+fa74hezhMUYs01ROVrwMdCe4LZX2mFj51
Tq0erKslk/Mdj2f+g7Fr6DDVT+3YrQ7A0+4KUlQISd9fqbSUlQebnK+seYWY5FZI
0G9FjOLZIHSI/3/2y163zV4iuYq9xQpQw/8ZsMNUI7uX7dT4YPUL9w11hezRpXnI
RNe78QWLihI7LJAtj87d41W3wTKXr4txZ2cIUi26jYAyLbAQV1tMB16FDD7XXKNx
9q5hNoNx6Vr67G/WPJ0yVtp+pIVVYTglfayXFMBEJv0fLSw6aZyRuLWtgpSMPvT+
n3TGJUj7ama0W5oy37PJ87pwC4bxkdGhmUu4fN8h9uNgDeI5EC/AUys510uGYg9R
VoEYWAdlQZ1gH6kBRa1YDgONQhSCVM5SPiQXM8BR8blaYf4Jn+nV9Qn8utT9YeDd
LHE7rTPbJKzbqB4ewSmltUammGpCNsqnVFyqOc7HDVgeLmH1VW2MDEYlFIBfH7eg
24GpqJiI0BnGRbnuZ1agM9mbkJESM7KNjGiahSEo+F6ichYoMoi5SfHkPFrAMI7x
Er5CuYx6F0O0M8V+y43S58orHSo+6fbhzB5q0KvMbnp+tH+d2MNCzY9/jA3yf6um
AX9GZ+3cQ/Mjn++FNQ8zzGpMeqgazj93YY9iuGGYd1lNtQEstNX3DFDG3Gg3IPKs
zPNlnH82ULaTboWw+jto3uscFKTP731cloh9jf86MVkauYp/mwDi265CZa5A7evZ
uuRneuOkrBz5dAbPK/MP58BZMTx0/0K63yPqUnmK2DerfBoH5G3CEdrpjNwlL/1V
AwQfHTdF6y1qzhjsGOZjSJqyR2etFIR/18Oj3r8dg4JPG90ElRLvHGSFe9DJxUDJ
x9OMk19JlFvSjRhCk/FoKpZpuPMTn4IdEwt6lJGeJcbvaUZqd9ZJVmTJVgPb6VUq
dBss3mijBfPTYger2DpfWZxB4tdxNqGa6VkK/HQk9d8ptB3T81UL9RQlahvNSObZ
AGrnwJSMLn2Z3D7QUyXYDYUkRT51Cf1MKKZemluor8o5HtKbD8d9H+xzuQmH3LrE
fWNh+ImJAJNMtph7uWeGeCI1/pnMb5Zrz3YAYRAjjV+ZkeLvPR6E7frsparOn2Fw
VmjG148w04TOSbQ/4/UNfUPSMqrWOOUb1MwjjRIGZGGgu81x9lN/hdEwWrSYJqX0
wndFhz//q7pTmIEq8Zs0DOG2Px96VupnugAfK5ffJQUVbgL4z3HqguHlnIrtAPtT
+mRV47x4zbk3hGpEj6bG5zskcM5GaaImspyn5Nx1gvcAhbaXsfng99FtPlnuzrv4
PnHMbowXtjxmbYAha/+4JFxu0ucvm38rNFXBjx+haH8LVld4KuQJ5GCtQSKbtXWM
14X8fLJPdcfd1Qc2r6OTZfBt3tQdBmvGj92MkLYnMBlJnD+hQDtUGNNuOP3f/s4z
CoO/4gXFFDnuXKo5BlSIAhV4NwnkqbLl5s8XEg0ophj7jpX/hZuNe0NLkT1oFe7t
093qF9kgOWwMQtVDuNX9WnfmXTrRi/a645EIod2Rez7UPFj3il+yXRAD28IUtn/8
PG+bsEVTjqn8g7YG1CawNF8Z498/yV5XVb2mA9SDQnB8+tPtEJp4DQFIcP7W73cH
J3/zp0Ze4KMYoK5H2pzovsvh3A2RSwc0NO+EBu1pGI5hZg3BUgKIg69Ss0tfojzZ
lfqi3hu5u44u+VtAlemqXi4qzHb1ycqKL5YPWGlrzxd+U5cDBk4FBRBZAfq43sdg
BfmYvtXfyeq+TYT2DFXPmxrzIVjt+UiIhVEmJxA1jku7gionFMZgD6yC8DTuCBG+
C8olkTjIi66EEfh4HiXGAM/SfPALQ8rMg0pKUFWxu1fSkIhgJZ5HNYoCqSmegPLA
g+h5XWolQ2kqOYdym7Ni8IegbgTgmOZk0w2NJmfHL+Kf3WHc4F4pEYyJfBt7RZI0
Nmq+pX98yc0uXePbhj2afbFwT8QLJQn63syPezoIh7WqZe/HyX2G4K/xhxdDz/cw
yGoo5mkFUuZNfCH3QUhP4ZeRXYfiV0iLN0BumVf+cvf6ao77Qd5zeWXtHL4Tj5NX
UUUwnQEbYQ/eQ76OmIL/kTSPdw54TPXHEz+Fl4Est8FbXjuEViN2mtIBiH58+GSz
WQM/HX9pAD6gjDeZ7TqX29+AtatWNEyUeAWVfdmC0DEvZDunH2w+wR7GRgYhaN5j
JJub05rGWIw2S0I7WkwopVdRYs7g5zrVAzToIRtteUzGTaEyK6bLYrTz3MxXQk4W
9CZZitKp0SKDYQMPmavmyjMojv8usHGurHm8rGFFAHFp4QOKkPLskmP1rtMyhkgZ
9PKQSrwDlXllYjyJM3G6nrD2sL2WtaoKWXVfm0bn68FB8fFKaSQ4z3VGsqRInKh1
6MGlUJhgOSoImhGtBy0JkCVT2SXkVAdTbWU1ctC08bIFOzkz3cVN9Ntjrfsn0Irf
oNyrjeawTnmyOzBMgDQ4oG8VIB29NvCEoWx9JEqHx5DOKDBnEt2RwivKLzEJCXct
N3jbFumlCieFF1dLxeqD35U/Gi/6EPqg8n1NqJ8VvPJsLuWe95eu6q/hJy1Y1Qry
fgOXU/daenpqJv4/QEuhZdLe2RLT3mSENvygj+TGd+miB4vopfU3yWeSE2Vpyz1J
MEK4f8voD32n8nfw3BHNbhPmc0wToEYbtQLsLJVT74Xzz9OZLM88MU2ZgdMlhTVP
v24aWJWxYPYO4spo6YIVTZ5o8y9rlgbiyo+ILHJCjSq/CElzznGQ9NpiTT6wHuV+
JhSnx9/sP4FsdjenujQMHeYu6EQ0VYPsgLPiR+3wviZ/YM0KEBvibSz3ecTcYEPp
u6xshcZJozwkibTrBtIpniamv43PGK2g8DkbggKywAoYEJn4QMKaytMMohtPHY1A
Tydgv4Bdxikw/VFf5U69k0IddlrNoCAz/6LAHID2zvvmiqqGMewnMBKEMEj9SDfe
CoTdL/f8ssFool2mbU7XMGtOZNsJnv+kYdvNu878XUskHqCNaOSpmTRTrSqfJ7+d
Zcz4iVTeXWIEMVnDXMwX7ZKMSFHJN+yNUrfbKfKWxZmEB8Nxa0N/DlN/gZ6OljEX
sn0eQ1Y+ytcKR64gqhP5CbG1edtojdKDYCtLU5afCJet024jG4yEPA3QioVIwWZE
tct7lBL4CWObN3Y0/gnTegu4Xn6VxeKY/8y9TjgWaApfzwEmGNbu6QDifUqASTyS
AtxF15dX35ouSNfXRLzD9SwyPegmOJhV/6k1daXyAIXHx3VOiXoACVShTl9NqhWT
o+KWIKSX2hoD9YqdjR+WPh4WDMkQxv6MEu8tz0v4gLBjOeOlWFFNmBonNG5ug+iI
9cIDsWNW1Epom0ILxiSYGMugw5FZicZPTa3BVvaUmrsRZB9nkrbV/eBnJvaGJ3hg
9PvKSxWyY6KwtS7o6XLU0k7wLTu1AaaxUfkntXVdOo/AlNXXi/gSYCgU+8L2vme3
Xmxu40ftlVInkANk5CQ2bPnk5OoQnIfUYgMIh0z4JLz3dkCRybXLuSMTY62fCh8j
/E+oI3Xjr6PlLryRctzXQ0DQxVzJqFq68wGL4VHk0CCw1EHae6o8axZAWG8+WlpH
Ifk1satYf65558UbDsJe4R68NatrtxKMcwSEZCu952vs9hErfwTwdphbKUjwh2U2
9U3gz8xuozw8lMGrlP31vWjyZxZWHhckfxFUBKgFwWQSXS1kpK+ov27YY0pksY5O
zO3tuieu4uE28gW/z0m9mrefPz/Mt8/dSWY1hT/bgSfakvssKzRC1uZxv8MWrUMW
iQfj1yahpfssRm5taYGcRrb/g/5yiY8oBHI6Tk8j2AwfMFzq/skDozvL25smza0M
8zXA80KU5w3k38YUaKinZuf64n836hIwhmGBrWUNM3ALPlab0v8PfNWcsx911eIe
XQYNZ7ivVo56WvZ8e69gqLd8rG/0Jtibs4u5CWvxVIwh84LDuRfrEQ+QH3d1Bt12
Zvzj1Kar8G/fbOZ17W9L6ckFbe9UzD6mS9+4MwtyZy0RopG4n2AOwArZFs7S1ISX
4kjCE4P5p7Wf13XOryFb+YPMvTbBBX7suCjzeCcBgwP73um8hPvirgsuU/pJHHlC
mHZ5MDADA2tR/rS4AdO2TkvO/U0uS1BSUCFOLokvExbzFobk0HIUkfl/qkt6ivmL
Ty2ILFTAM/CmTqNNbn5OJt65GS+8Ux0NE0buumKo+lS/1j5U8sCOHctyjQS8FV6V
lLck5H3uNanpFgRtd7v8pTV9Qb1rmgGvUNsNnLvBTC14xVTRhwkV+ls7Vp84Q/7B
ec8vjyRGVyMZAjtdgCNM7XH7F++I9MhPjBVmA97AyL6G+Xw5DlKD8MjStlTUGghn
wC3iCmVlYSedWn5p4Z9IhZQxBeugwq7/Ge2lpUGPP/M+PyvMgY/bKeiYrerEHmR3
+FQM4x6ZIdZ8wIMtwY7xDoKdBEIOUG0C6g2OL4sdgNEZ+3hO0GN3BVR8kR0+5Lqi
wnpMDQA7JuUDLLzDqjWROyjVL8EJxTaYZCywKbRdUz3+RP4JvAB/+Yi1cJW03HKG
rwAB1By+SRj4CpnVkMLpfBHSL51tzh3IiAQKpHasROIszw7aR2Hf1XYa4idwUCQI
EWxbn9otHchsmyOQm+tDewQWFlX/1wYsGGHuXzl+UXZr6l56cIVa2Ltp8p6JLLbW
/yzPO+LZTFodutyY0VHjL2EPo8A+AEi/hM15CSGAXPidwpgadKkorN+AhbLYhHps
hMdWpwzvxlpBSeUUheSgSrTVUYbNVgpGTqmJHSs7Df1YTye2uvbFBuX86QypbGSA
53lwsKX0yQl+0rzFWWexjg7aWp0rMnYnIvV4zRCtVqmIbCBRTGV7VQxsW571VT5L
mqvUNQgi+IWRQLJxMNv5V3lSyHkv/K0Gt8ex9OLkRmz2/tGYcpT7cYoD+v1A7uEw
W9DBbzRYNQhzGyUy2whON1IVZPDYlu15fp8/2E4Wd5jBtjbZucxKKy8Kid6jgRly
FJAubVRZet751QLwN5ht2PByWjSL/4OnTd2xDmlcCWHlF5x/bnZ1MZi736tpnABX
WMrM6frQTFH97oQctmGrrpRturcQ2a4FZI0qGT4v97gCFXVez1TUXl+2vqZShJ0J
DDmZq8lq7Ny9OcyZE8oREQwwiV5RNHUFYwtRer7OBoag+aO643QOTf0K1WZAikKa
eaRNQj1kYgm3nBP1gnqrCSaWQhBMszg7cG2hAOeXG+tcThnbaVsEaqwzgZuwPVVQ
8MWXoFKsJE5s44DzTuD3ZA93A/JCMiPUt+49EVhcnZdoENg0VzIPfwq/KCsbH+9X
lfg/NVyMmZQrhnXf+eZapV6xdTTQruucRYHeZV06UjeTPL1u+Snx7UGl9xJ0SnNj
BdmIxxdlRzLHGWj5q66+QCT7f4z04/CZmKU9X19fIzEfx3rz9JNk6dTCHlIo2uPQ
DyX/UeArOAu0WEMHkvH84kD1J060h+nFn2QdREoBsdX/Drcn0hLuLPASfLfZqkVN
qXfnZJ86Yi3HqG09US6fRDkKhuKpIHbD61CVViY5yX5OqerAFHpKLmBOjrz/RgX6
T9Q+8qWXPAwrrn/eQnzSvXZLUULHYrQ4waIlE7CqA7SocslBfiz/GRB4bBfh8+cr
oLCimDINrWjxJ1tMN7DZzJYvwBNulB9PnhqDKZ6kRZq8BXJ3y6ipkR5s8FfB3uz/
IXJMytDbw81eRwu1CHMV3Iim7vGaMtLn4B+OEUyMgDjrnUDS7HbTZROItezjOxGo
Qry4Dnq6t7SYwtfA0+HHD4sTwAspASuO0hXttcqW5TqhhuCaGF8Y34FXYxoUfJeL
X8lvArwyRZcFR8d2iOTpCzCGXUj8c2HeRa0wiXfhFX4IMdYP9WHC3Q/01xjGLImY
Zo/naZ+u2JJFN47yfrNEO6NMAGe2Q3BtMpr+MNRNESe5opqw9P8fYx6T/krX/EXL
doyXt+O/Chxe8i0al/V/uyFlD7eFKVw31D0Fwc6bUorK8aEvJ3G6jYf0MnukCBeJ
B/714pXlk2dAH4bDq4ztT7hos/mtzr4iollIUTNDjBQB+AiTNStROwJFa26omNSC
keSZ/kNAO/W9mrp37xet/9NXZ6cPDOkXa9bOYYjSUS5Z0mwPBnwVj4cR/IwhtNsF
u8Ab6td0UK/YPHWIymRn0FrsR4kCjoGx3rziNGA4RC9e5KUjs1j602UkE7O0mD8r
U8CTYP62az8FYHM2Elt7SaJuIlJxh43Nx+Hl6TXk/usF2NSvCZl8EJaIrO0X3r7J
eTlKqfu3INOje8VvoTMo2QLWYB0z7SQb2RuydmTREeV9s5oXbXwtYEDH/DagvhcA
A4Fp2JhYAMcdQxxrV1uoGbxdnPAwPeZbS3Wu/iLfU/2Yn6upGZ9zITouzqQ6LFZ0
uEBpVJ0CAZ64jQosZimNEYwjSSWg7wlREDy4mzWY5VJfyWm+fT2tvGtopaqXU0gt
71s0qnIZxoeUvBuJvTmm+YAafHcgms19i/Euq8DmFDN3nUS1KWPDn8VHsahFQA1T
hHkQRJDa3AUnOTLoGAgiSfkQaXZXqSzU0wZVljJ6QgYfUYH711nkZTEW62t/jOvl
eGQCCugy+P6f7pCMojBF7Mzas+nWoh7Hu/1S6BaM0Snvif+QNKGrP5CAbAP8s5ar
nfoZP2wDTbay+04i9wXO5ItPFkEoTSMWrVskii48sTrDp93txb6xiD/LBqBVwhH+
BiL/9BqKBtbKluWOmoje/iZN6rSKFZ7FGMIS9oCpx4PrypXk8FlXRptm80QfYSN4
6vWcuR0Kdy3E6eQZBzCfTq/4SBjCnVuEDJP0HPuVK2Xj+Dxi3g1KM4PBrw6zCpT4
lP8ZbJWHhsQ8xKV0g00ltYsbsgUARPol5YZ8ESPnJKxy8V1eGZrriAwKzSkgcRzt
+DTuNfdbmqJbPDM4SQNRfxWMyZ9K0DbXoXJ20KLvVqLcukcb2W1hCYPxotjMWlOd
tBGFzrR2cHHifmmShw00+oTvfgKq3vwk9zhBxlz5B2CcOwDETKgtxPWPMtZksQE8
MoTTsBV4kX4w+DQIvv8V2qtHfTRBQyE+79O6SyGFJ6nrO78fyt0lL5aqDf9diTy9
E2kITSDfZ98lzGNQMqt59v+Aj43EJkCnvWIDXImZ++UZsFAx/TRROcBn0RAJjABW
Ba7NLmnduf4/MQiVGTWjRqXaHT65b648MopHEvEZy114sfR+UTXoUZHooDQ8F+bQ
QK+y2m4i7+O1kxacrZpBE0fBd71o/RhhzQUBN8gkpu6lGXk6j39i8wF+TixuItxj
QzkhRpD2UndCfy3wS/hvvvQBO7Zs19B/izXJ02aJ230AkXShBgK/Gv3HP86q1nZ+
LPbQF2MmxF4Ny9rb73279vmDn6YhZQAY1SIu47sY3ARJ20qO611IzQElTAq/w/jo
vVgCZuH32cCPlY6L+JdX3Et3iLSNybg5uWc3RWebgC7cvLfYvZmhfCH9bSas9C9u
b0sFNh5H6tjogHMSNM9EIRYXWLNxoZgRrZOrRHlza7L/nX66vWF2dADonEUpYqWi
kEOAPlupLwQAAaUmxO3Dg0jKLINQLzq2f+8eTJyInMHQbSoCeAWnxqAVS5g+EljQ
IpMzzfCivVW508Troy24RfiwNWF2GXlpElr0V30qAMe80n7f+/hiUJqaM8jmLvph
IA5+aHgy69JnJUAJwXOiwUgIWN3Nb6npUkGSWNKFfBxGPiJeK3t0zTaY25L1gDBf
cMNaIAK2OnZ+r7WFk3eQ9XM1drZFWxltUK6dHSI0nr/hr16wxpKnXy5U5vbkCKql
wreONeSJDDyD2TaxdVT38n9EDCeMp8AHxhBtg/J0VHhrt6t99PEl7lYxvkO/LoL1
ws2t3aX/SdcE7Ww+k9acVHrNiHonOhrisqs1pPx3XDSUysAPEUoi7G3pTo+enSA3
MswBQSaUUJkfrTv8oxLgtuoAQ7wIvzDpw/CUBWbzd7clTyDqf8sAq7SEXE4/L5fE
XNWTUKeIz7Fx0SQzq+BUZLTAOk0AeWhgWFkPFa9b+C7olXfG7g11pLKTEaIxQpuT
AdYEkSGe0e9xG0z0NJ5XqqkiTsvpAlpfKofrIGh6YFmkUpT6E3bMnATdlmAt5LHn
GhYDPFBYZAX4MlS1QRhwsZRonXn9yJzYAPlR93BQWz3Y3iyfRp3y6cTWgpt+icyR
oJRNZ9IkV7os7rMy88eNYydhxj7k7vc2VhrImZTOlhpwLLq+TT7Ffmsb291qbmeD
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X0vvNgtqDeNylxXxrN7pI61D2zor5bgOVGjSV0RDpDHCoUMkl4sGT27xBz218nBP
e46n1/DHG8bXDZGNHP00+KyFzSCfzwVeQUFKSnrfuyNR/GcAfNeBAS2cd3s7lhPw
/f7jDMSeUDan7pp2N5To6GxgXy5icPzMty6KDZT/ljQCwJ31YCFK3PsSIK+GsjS4
E+gWS+fr6HsmnuF0TcANHTaJ8KnPFz9b5aFunec3WplkaXr6EItn5FZx4LS19o1y
NnwytfH93NLMGRVbYRR0VaUNAz5vw79HiW7cDtew280zLZSvVuiyvRce6zd+6Pcz
/9eXKRNWCL5bilf4LWx9oix42sqkj6CpHvl546aneKFY9vj/07NBTVnrHMDDo6kX
Uq5y+1sYIXeLBrY+pY2HyY2/2+C7rJ9zzEDJ6Ji8PaqM4xwRHxozd5OHiNtVYBlx
F+RZin1HKl77ySmhPBCRNkVQXvztL1pBrKbIB0bsE/axqBeQlW6N97GqgE5JZziX
9iQ2GwOZbwdPm6ThLNdARdN2GiPeF/5NzNXZJvgQH7py282peLjlOaN4Tw9h3SC/
+qhfySFEIIdIInZn0P44XnYdQ8KTtRaAkYy82501zb5fE8xrgcsj55ixLilzsvrB
fF8Tevtr8RZEagHxEUcinPnBX7oKqZ+kkAPIJgf8Vg3t3HxuaOOBLZV/W2ZbFene
83+w+gsulj4JDpVAJfdRL9rF2jX1c0vKRvXDMgOAvz4rX0LBbW4Uw9Nna8D/lK2c
7UJ6lP6VeE9IVI79nQFpth2mOIKp6yXxlv/b0T1r8HMWvHYcdTW6CloIlSHmqXqf
qDxlxUY0xzx/vsd6PM/ciQ==
`protect END_PROTECTED

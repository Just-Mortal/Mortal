`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RoeOKuig9aMbQ7AkCYhppqt/AtV62pDg5+OjnzijX3tvVBb3A0V6IF/JZ2DzYz/i
/Fcr5o5aUHf+OUE5C+7W27TBoaSH15/dFZrOEdYAVD3NNMU5coZXe6xzZbgacpYm
P2FQDAIL53jSX7xuu5NifV0qkjdwJoNMFVH1HSZK791Znkm/uYIGAaDdveY/YTBn
LmEcjLma6ppjoo1v48oPesdytz6/du+k4cZuzNEZ38EZT2t1aL3L41jZtyQ6qk5D
EnAVS3nmzLl5Mm4/wKyjOf1ixIxSyVFF4HhxNicPaXEavW9fLf6sVFdxyyWMtIYD
EU9sNOq+oMbxlVb6s0B1UO/IXpJBau2RFka9Ru/mbacRldQ6+fVxLnMo4ipRQf7n
arvTdczH25n8d/Zo0cxNg4rRTfvAIThIECLC0S+x12E=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Jo0lvosrjhNhEUduNSLuFjvctQKF+A68AdmuIhYmR96B75mpszuqRBgN82Q5tcp
LNNNoyJ5Ibk9hn0s1RuIC4QWeR2pWsFD7bf6uc6i8JXxyCRb65E0Ruql9hJ5RXvz
jRg2XJYclDQVyjbcutYqqQkxiOG2pYI27bS5/T19Zh8LqkJxHVumE4ttUi7Rscgu
7lMcbSJ6RYG2RoSbB7q8zEibDPmH1HUCGTs3JpMbYkmeWQNT4jbx7gCMW77o8Y3i
fKGYc9JYG2jp3NpvVNByvAFl2utph/4m1EbdkVgOQjFELxfZ/V+RMRLqCSgbGGZo
Z7cJndu1qTCE6Oq/eQ4W05YV50JLqDltJRswiPK83FI22bOp3gx9EntVE+hFLbwT
7/JpaOsFJjvy76ziHCNwW2p1dEm6CM5+wDviB+SFxZwXhdo0WxzUiAAodzVssdpu
SKg0o4ODeergHqdS91S3TonGPbOqbObzaTCmYJFGZiJm5vct7DPpp9hIwNr5SlPO
XWSJ669A4Jvbl73HzOS726nAUoVLRcSZu+B8Qj9N47wXHySGDfGetF69qxz29MhU
8vA6QGggSHECbJuIxTVb1z5N6oHxAWR4RdgeSjIqUR/tlt+vJOLdBk1Q0V/g5KH2
goMk3Wu8rzxvoIJc880fpH0Gc7EZBtIDWnYN1BioMrxnuAqvSqtg2znIFngXT69L
XHQLe3cyzclRSZeX6yI+1stMZPv30usbhU5hZC0Lsp+2tvjsrmLOniuucGXXyKw/
abJpR/KMjFzukm9MbRO2/p8mK9wpNWP12haw8Dc3LaL8C1vcLWxNqixFMoB15L/4
8l7hCj6s/aMVZ2GQJZNv1yTBedZdhOlaLrxngQUbySdY/yeMwvxtX1V2cWdfiQ3Z
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKZKzufHKb5MlOXJJJPFYnErWsSMrIxDR8Y0dp1my2FL8uVKAIghyc8iCVVbTjHC
MH0Y0zQpgIWRMAJU2fUS0Es2ooMfmb/OqurdN22Wpoti09b5vM8DHKGly2f9vXqo
Nk7sDprklH6Ltr/MNos4ETZoM+v9Fa/Ou3PB6z+UBsxVDE4GAbNlGn6Y9UujWnxa
sXbsJZB8MMVoAgAXPmZRz9UpUXdyHWeHCiv1TttFHLDV8YmhGPzZU5jerADtJFbD
OqgeSOC38QhF3XYdSCtj0oNY1mobg556CmhMfezHznc6GjwKzashnuoABNGdiqfo
Hza3k6Sgtx4T41KC83CTGJKcYrn/ME5ClM4EI7HKHh6MwlEY+Godgh3vN5pVoNtB
5iW/EW6R5HFzjDuKs/JiPHBNvs5MiXKfUMeGG/rROHM2CGqnFqQDdxz5urjkvqLz
AUQZWLks0ltERlI83qvPteZwGUE8F01zgxavg8VxNjt/nEchaYQ9bJXTG8da5v9b
q89ZtG6gqiiVmr9m3Q4feZdnbh82FxpTZyO+9f5r1imqFWyhD0HKmJT3z3vL7O3d
7W6bGEixNGamUoHldhZWxZ8FZ3dL/KZsT0mV8dC7+vnxmYNucg8A8owDcu40wkzc
ywUiHDlKv39h1lIp7WrLaIOJe6cBQuH3/gb4J9nG9DHfHEKGHCjMhrUkkj7sywVr
NG+T/3pgIT3iWm+72m2YkJk3E6hhqbIfSyioQC3MVDgHDk2zL2k/OMv17omcYcV1
sr6i6BXe1sO5bs9w/+/s7NYucdoozOsHl0ZVmvg2u8E6eWpZuLJb6H9w0naSNv2E
AoOAosWahfliIk7q7dnqGkC7ITOFAr3qaOWqXv5qGxgXovZkM14q2KV+hnGANdia
cp8JryxW+MqyRKAuFOcSgiI1KCjhx1xvS5b14z9OBMS18kObBSnIHmQqIip9/8Ub
SOeHFAmSir3fxXOiNNF2ERkPx9eWhKpdGeso8R6l1sRWbBUpLmOcNOqehrsgLIDv
qDBxHPo3K215Z3YudjgU1Mi7Uk+YzSHpkoOU/qHvnXx7ATpAiDCxtdm+ylT1fPbn
MEDIUsWDt+hy+73iao3kfR+J2IXBr2uEHZJYXme4VHuCqdEoJ+P7v+E6fAnOAipj
JUwoTa783kVojXrOyAZkrfhXOY+v1ai0PAmlpWHel+o4XHI60EQN157b7VF6x0tJ
EHV5BMN7Ejcz/VhWImXXrdeeCfzSxTeSCie7ZKqetmoXHjRyawp87dXT1H0wTLRn
QmlCqywvAle6tbCi7fVD7UYhaagUlrGDhgK9IDWEoGaZdUZAfuJtbPd7Egzh4ole
pga4uwFCms8di7q0XJ/CFuP4UhJA/zhl/tLSfm6+qTb28OYayLvRHAu0YVdaxVbP
YpUeSNOF3C3Dvfr/0BKCh8hYCyivE7D0cCNgR9SOnuQ0Nvd0C/c13OaZp1wN/690
BXKGYJDmz6Gvif8VCsBEan3IFDemivZMAgW45c461KGsj/+JEW/zy4DXZFrya3AP
tmNgS7u6beg5yb1xYQuu1ZlI97pFuIah5JJCcB1++QxJEtxs1glDg4sPgO0rd/nT
MI4eRjyxUnZ4qM5Xf7ze/ng4wedDulSVvL0fVIiZwzGl7xlj7ddY599nzH02cdnC
oLs2wqxkDf9KvhPMcfUo1H0gbVQ3a7HcCOXlJPukU7GX5rXN0zXFtZ2sUacVptCS
qSjQVImDIp8dqOy2D1C+0t4/5XtVyP8DsnD+JjQI9loFEBjqcg2ESwQfjQkf/zAk
ZG942hCYTsOKTZ53g41T2+LMt10jcYXDBgyCHtdGiDpCguJKN8XkS3RbwcUXyLH3
CZxxVpyjjYRfr2JbCR0QqZ+gv7BOFLESelX/QYVE5jFbXoSnEmG5oF+G4IkcLKdz
tKrQz1EbF2mGqUWxbaYLoJgQ4RLMBYzwPZVUbIbHcJF1R2bD74Aqtn//rXn07URf
nGDcmB1zvT9oDakxBhjCiZFavCu8qpfuBati75wxVoyYjF5bGnSKow4L8EdC4TM3
JCwBhlazM5IyILV1o6eAWUdjUTf6BTzwtJdXcBB4Px0TSS4X3bcjG5OCOVXi7WBR
RYBOHdxaNOC0pgHi7njgepMPdQ9ryI+W1zedsPsVjULTo/ITgA4HDsjGxPZufR8p
icn8ZPiY4fEyzebpb8FaxSAhj+NIH/jOtCY4iCih0TrpIewN9XVZI4K2sy9CYs6m
QiORamVYaJ1FXtoO/tUJADr+6aDIjYcvV7td7ClzPgtVVXo0ljqS0lSNcy61tFiX
g4zTX5mI7dFNDe11GJJKrubMbGidGF4SeRLkbOLETMgWOv7IA5+OsZ4lu7JofAic
y1pGqZwt3Z/mk3iIksg2DQwdFUHL6ie+lc6OQhSQn/VbD6QB0547vJV5V1WYcW2t
i4JCCtqTu6Xx/AeXNYYKFTxfN4b0rz1h/mIHq2U6WsE8Gcz8EC/w6QryVkU7Jjzl
chKm6OMEmqGMp5yJfzve0ho3f65an3pz0YNK4QodgEpCtPsmihww0Sy4nCuSRNNU
QImKzWE/HuDdxVZfNZR3ZshUxDbwMsbYxe24NEC1VqrRiNRdfwko5WijrJ0YqPfb
29phkUl3PKQC0dc3lYXV37fm8GcpU129GuNaWpjeVmt73NNQKwqw3fOdG8TI8PO5
9tY9i8UEBId8MZAocHdNT/bvgZauLbaur2UewbsKbSh8uYufRhjixqe0ZgUqkmh6
zpEInpFgYC6htf2DViTCAK3SIQSvrdku41bDwZgDzFZms+noZIQpoxbVfHl5c4TM
gIIJROgWTFhjd0RHKvm+cUyNFmJF/VLRFdXYuJl4BIfZBPLycsqO53DhOSqHLEES
gkeTIK7L5/rKLcNMDEemLrMSWv0PSL3F0OMGhvD1s9Q4KZNjuzNxKMJ6WhgBgXQ/
YOaT5fr7UBE6IAWIlLvykDpRBx4cKHh7rz621tITn1Dc7KjBL5sjoxtqvtc5tXhx
/sIV81KAVepfnFDQe5nGdYN0Qg7DUKNsZW9/2pGRVX5JpN76k3P9idd7wqfWoBTH
AppmwKe8Y5sSyR+Tj9TQ+qyzs2ZTeWkT90G/vNu9VnqBcmUJuuUbFmBBIO3WhTPM
dqDfbymC4haIujQ/dYIfh4fgxDRpVsyywmDv46qTB0HJMf4no6j0cCa1VS/Qkyhi
1G3mkcLbYQ3NkgLunudhsKdJ7AX/TYOb9dRuDkLwS0PUmkBOqL4q+93RBGkb6VPU
u4NRyCALPyT0ANCgSDKC3uOcbgK+9NTcm22pUAlw8WTfV0+KpdUVPBtKxRKaq4zS
OGWY3fYxJm3JokidLyW6D00EkCO7SFlrfOqDcf+q0156LGO4c6hTlmfb/tt0mXQ5
f+gzTfWZJNd0woktHs2PHdDHMhod/J/JzBTot4eNHSmSaUO98eiN/BstPMHEvo1L
nwRrXECngrntAWe5CL5mafzErs3tlDLNcI+EQ0+el2aqh5OHJw57YP0CG6J01hkO
tI1AdT7zi+wWsEVVqbC0YPXCGYQeIAOqXOWZvpVl0yyG0EXmFCo0LKDDcnYD+oe5
SjWA+TMCs+JEtMjHF4eEKcvb38BByg+D+pqoc1AUhTQFd1mZTqU90810KYsc8MEN
2SqDqFR8RKBiIU66Emw9IrXRoizSREWM99pMQ+ZtTprv+TIKn5svLFuu04CUfPzP
pJt5n4XhkG9UbqvcB/x4kmwVvq4zVniP4Q7+FtJkgMKyyy7xlIgOa1ytXGq2JJNj
46N0LbKL0JI0AnHh8vLnyTLBnANTDGjv/Var+Sq6Aa6Mwywdg+7tZaFNFxy9nnJ8
LCpe2E3QBW70jD+CIWWjx5I4CedlVY5L2nbZjxiGkEg8+hFBTFuyp0bgvzZ57uxQ
g7dwNCLMb6+OzaaOJ+FyNVlcOtggP9FW7QYeJ+xMsZqqBOLNwrBmB4BbI9gdguXV
OHTrs9mQG1kuO8WfCzykgLfY3apARcfJYS+F4Gln+idwXUxPZUBvLArH0Oos0lXq
9tvazNOegXU67MF8IXqQhOju9NZ7OFfMN9++dskNQmjwdklUftFvpMBzdOa74fzr
n0+sIRsIzvFN0+MDpCboD4cXuxlbmMLwrUCZanNYJ1vlSChYzb1wIEvG8RLCO6zb
dT5Myl20n4n2rzzsoZRPYAwkwguY8luaCH+2mUgnjuA2JyA5q+ai3fue6WNK2wDn
ZXmXER4iPw1gCu06xE1Qx7aJQ3pzbDIw874YVfm+k2yhxsZ2jw36VCigtJYmLZeh
HCx+Bbi1mRG39IIxPwiSNLyoPRDqytZWgFdcVqiQu1Psn5MFtTOzQvNBYUqkLP7u
OrP2Atf/PS/9g/bWQTbfSSrO10D2Sz2b4keBQLcN4YWrLiYfIs+LU3OEsAMxIKHt
kadAPGk4OiHbg2LrMJkkmic9eqTFtXJP2zIgHslpQZJWWAnxaR9OieV+TRxvmAP1
Tkqmno+EnS1t50wCzsDKsupMvuH9M+UlxXk1GGo7HM5EbDlZ6qDaAAEpB4WZog9n
4JMxMa237xbzwJwk9uOsL+fbaIiVSkT2Y/DsPJZyG3SpwN5oo3S9+rfeDAUSsQzm
BrGdAbPARuibuGLx4hB0kkRxEYl2MgZeFESGHmvxiHYTPE1+N21FMK03iLh1NQeV
oB5DKs9Z5DRZibz53RRIE8kjy6/URMiL+yRuYqC5ZyJLgXc1cR+SmK4i8ndXw3Be
og+RppneKkc+GbUTfPtTIzKGE+u6PjbFD1emBwfey2N9LVvBYFcvnDGESQaaGcae
JcsvCnIhw7bRmqMGrCC5csBNqBtm5ijGuuUfrpbcPA1XMsOg9MdMG4C1yDJuUZpU
BcHPIiWtAtFqqwzRsPCwMhe68RDPa9GA5pWTxkMOsC0qI4Lve/B680XjzVgNCwyV
9kexdUSAnj2UhFi1mkHGkKrnzTr5drFB4eAANWLTDF1nj6LgbF8TKjI2SizoYpdH
+EnvnAmE4QYCFc7t51iNkN8g7YKVFDt7vLvS8rgvLsqumyEdegwt5ay19TPugkFH
2EnEje8XDlYmOqZbxKPTJ3Md0AeUiNXakyBmmwAEWgcubYmKiDrwx3xPl6BOrJRg
o38Bgkh3tP5F7cTUPdR20qwcd9/N1k6DAPBraw4XE/+je2uaLRXdT0OfBOjz7Fiv
sDVp8oifxJcEHpa2y2ww8fHYGGTmHzDQI2W1PFNICR8LfG1bx8erWgEbcojf+jBl
14fqJmLsxDcJO7P0UfF+EF+FxUHXUN+gw65ViaHZ82GLRYk5h4jCp/P3xBYLSDhY
QQ45EuBoyNUwfMpBliY2EJjbQoN6HpFUBVQWH6gGHPLNgMF7j9C/nW6+lftAGbnL
3pPxgmncn6n09C+/Ae4CxYQdDZGHsDcRaAONwUvFQlecOWy53x8raz/HVg/w7T3u
8WMTwTIthHszCpGWaiFB3xipxLHLA2a5oxut808264g5GiLCmy7xMGm7b+1IBfKV
vAZ4eDC37FpeJz/UjYbi2qhiBbNEUTw8AFUS+dDKlnoEg6n5ApjKC0Sko6QIfK3E
y6rrq+4UgiVV62XFATuvJ617VPp3h8W8BzWIBZXhkY1NYOP3XOl8gnIp1Lq/Vjwz
Mfx584rAAdy/9gOInzMGjv1ZiIVvDrSZVhy0/AAPaJHOzZs5CSK9tphz9dy15lGb
9Hwc2d1uTdt0feWVv+ljHk/Lw/RVsnRxJmTjOypmRl+TAtJjZCHlb7IwJE5MRf+9
yUM4Ux2eJfpyVZr2JMc2mtfqUUsH5nqgg6ywS9+gsDm1bSe7S38PjceydYfy+VZd
xDWU9JyKm5sdVhoWCk/BfG85EGu5vueio4Brs0gSgjS4pOc2U3ywDOC3pzInx1Af
H/Zp/Deqb4DzM9bzbklQ/DyRfx6dW/Py4bv/xFrmTBldq6jrBnlDPlaO0/vjQpZt
/FcwO8Ycgne1ukykCIygpPAkQWYaBZIrV6f4MAICq+yNUmqqmw1FIJB7Jizk7pDn
ECj0TNDOdeIgT20c4Ytl9c5UvL5a9cHm0DdIspxqATKkJ2RJ2s8N67437TE3ojlK
yMFeY8lw51M6MfNeXblsGWZHhwjkeAXq0MLnmmJ8qb7/9cRT1EGiiwg4UIAEfKFY
kFkJgQcYJf3cvaPXFmfEF7bEnvzjNJKxR4aIUjPSFdyeP1CSBQJsybRgE8xsZGp+
2VeuvsPNFowmpD/sVnfuIDwCFludwqvVovTkzLEzRYR3umHc+EO6ROxcyqB+WQf3
iwzitkcQSmlcyUBIBZtv39/8PdvHqOcquHEQqSB0/xVON0//2+LKwmB0UrcBa4Gb
WYiE4p2FNHY7Sqjhfdqnvd2obCj+NsxZijodhdyBEMbIcz45x+hJqg3Ew1AXlOZs
5liKvfdKX4FVhkj3OEljFN6HaE9bbPmFRbjkoC5YV+8g2pedD8YgWmhF164TF1+D
WQyxr9IgfsEwpzf7F+U+UTgwP0MB8da4fOEZbp8PwZa7EGSzBFdabB+PLEjHSi1e
Zel6Pwsnt0echAqrYD9pq9KHRGhkGtp4bctQ3OZk0a2Cscur3OsWXrhGTyyVMphb
b76EfTLy+unAdaOxC1IYa5LVL4tZMruD3EdeQx9yP01Q3ofLSzK2lBHaDavlWB/X
Knkh2WoBc0RjIf6dbgRM12sKbnwGn6nyURNdGvaqkpwv3jwS3p4L/YlZw9Amq85Q
1VsFt5olUCy8ILqhMM/LOE+zHzhc39Vc/1KbojAyKprMsirEp/VwO2IjI/dmooc4
+5+5z1J0iKvbEvOX6CVrBbkBT2TflrYn8Oz+tAaXMYRKcHHOp8wZIjbs3NtlXFNw
TXUY6djJveRO5eHP1epylguhs5C9Z0KAZtZSC+0e9S64+eeublR/d+Et+TARmnCF
5erjMTQqO4ygsXSQmaMXvpHqESUgDGc/mK0HUq+dE8NDVQL5zWmJNFGHEUqj4Dtd
3YQ2gVhLc25KrHFaNg87gIuBQb1stvFtpFrpYIKPK5WErb2PQ2tKOhsCZbmYor8j
x4Sg+RRyfG37My+ooPGQMxrr8zhIm92wUIRDdhLK5WLPEFEsd/JnVFdZ9uBzTu/D
QJvj9+310NrDwGg5dYsd2LU+exVQENzUUt3CDaiy+4RZUYmnOM51vtzVSHOcOpBW
X/DOzsZDNbtCnhjaUDV5Qe6ftqCmf5mg65bKA11DXSF9TlV0JyCKN8BJfay4Cfg6
jDvZAMJWKpyW5egg/p/10FX5aLPp0ht/4TfexY7sfp2RVlWKemEgb2XdhwiLH+9N
zwD75/drKhR4xK+kKjCoxgysd+3123O9bmDLuhPWqjIotUNa1WiBtnGi6pXlbYUV
wRUQ8G+/SzR7BDeyeigj70KKcTeArMv86XCpc3RvulMfQQQMtPEObd9YCEbKZ85B
X8Hz6SS4LrhCy3BpYM/O6/znB9Lmh2wva0Q/P5YhLSCY7l7i8/vGfVTauITlcvl8
fJxrEHKNGfUZ0bgSllJdH6A2Jst3TMU1SHOrQnyFcBje+WzVk4g/4febM++v/TOo
benMWmD4V+OSUyD+zuMkEWRhPb0J8dvDbTiBAYD0BTtnEzZU1wE7+gjSmavkjKYe
T4PZgykQFqs6jZq6T1fUjfmfIEMIbE445jiu6vo2aS0bSUM7nf7CIXvTsrSkF568
2fHjqKGxxCOt9M9SkRFK87JlOltMYar+pHgegJ/lAcY8MxsXtUMvXpsF/8u920uB
rPs6Iy4YBfN7mduEHFhFL51/Gaiuzxl7X/Ce9fOscEUY8V/o568KuOcNTvFRb53e
/NkAbxW7SoSa0SNhJtrqaLF/zPvkGELkzVenvdwd5byRrYkrSuzt9QrZTiqgvtjg
9yN15wCytjo1F1Q41PLm1lSHGSMY1do4jxykTm0jOEhehud20ut4rG8VBwA5x+le
1ZIs+2Xp7watQHN+OsHhTm0MZl+EgwRfdrC6J3dL9prodf6BbmenF4rPxk0kDbRJ
Baqlfohw5JM/xjr5M5/zXURJnwXgTGsL5j3bryz0OlWiTgIFh0LBpD4TqRRiCQq0
7xqv/4+s0utYuZ2uNByriZvkOEKPhnlgRoBYUjd5leePqkmk4nqpE7LjK/YcdC+p
obnyDA/ouS0R8U1tFGOVpk7iWt8gsXD6ug6kiMMSeY1/uOO3+NlTZ/H/SNWS+X4U
6GyytJSEeFWvznQbsSUMazjzrzuG1fYULkbwg9a/+2cZITmx+b1o8dsKopUz25eA
Ikj2FVagA5vc//K0XCIU07b6azNptzcKbONFT/wWCp/Lpj7dsrdfl1xvLjhQTmVw
jIbNA8vbwBU9RITI4QR+mT54UlxQwkmxAzx2lX9mQQfyUY1WIDhw/PevVCODiQ6b
lUI/JuyXMuzs0QS6WSvFJmuUoTTUjrQ0ZKeGW774zxrHoh56Q1taLkohnW6TloQc
4r2lwP7wQ0OXtgOAkAMSjANgnrPiISAd0i/aEPxDsMZgxa6862XiqSbrHbVBtcEZ
gMM+CLQ4wh/CNunIBMbj5ADIi+/ZOvAPs04ZGElZQC4IBFb+SeN4pU1YDesfFRq8
2HdUvKGsOIuD05IZPV2FxzZKOMdpll2sFhG8KIvzzbXCYxtofDiplRw59/pwl3cM
TUBUZsLSn8ZSm9Bia7loLFKvPIThJ6LwyqHESbAc2iqSMBhKvPApk/lvXit/J51Q
9BIO2fINKYuq0MwOHSlK0Qmn8PthqPc/1bTQXt21wJnUs8BDDHVrac363WeyKx0H
7kZHHh+aTX6Oidhi75ncEW30v2IQyWZPBCPRdvrAIX8WEMrWxJdpmF4oVknPc0ao
35eRIh4FKeq15XNWBKpfUUDnFa+PAKEMbWtz2zkHbmI98t17LMJ6sGA2V/OrhAHz
0MVhFfRX+QNnLOtqtatDvT0qjWCxxDmuPpG7+UP2TCQG/bsaMKDmR4gq96cPgMyR
4DqY66YmI5rqhXEl97GU4vBnpBsPGRzgWjMj9A1V53/d8eFqCSdWT2ONjkAFCOHt
XDp8IrQBYGyh5pHWjFUG76dcYjUiA3VY5z1g1F11DBR4HBAQVIgakP96x1jNguL0
v8kZtrnqta4Hm4YXwOSBycJJJzdAFUXyHlueCgALlctJ6SYv3PrFDQwGyvx3aDOO
vcARI+BX4SgJK8Q9LPx5+67NuKZIKyuw1QeEy+Td/3pS0eZqX+nFYOxvo0dSKcif
AprGYSVtZrwtncIMu/6PilD9HTmgAIwqXl6LxaDR1waj6k4oarn/6HrLSrhBJ1nm
KE2tH3rPjf3Pc+lsZv6RmO/I/X+HnSdCqPPhvHwQGQtPXIW0G/qZepkwTDhNTdT1
R8w79Bn7kM+iYVOOsW6FwdBjuce6KkHsQlMThJ04u0V/B3gZFiu0FyC6j3gqBKDm
7/B+9i4l0ycgGsQJtcqq+0EU4wty8VsNPnIsIbzMTEvaH2fYA6n6B/9ctR0GHPe6
2sYlNbkVtGIixkGBoGoTlqd2W6DpzkP8MysjZCvNfRfX4AheolX1wS19/rWvQR0k
GF0SIRQHAUmysEjgs0IyIxOH0/QQvdH5AnBsWFKWQCENwIOc+gO4+d/GvaTacSfx
1/whXvRRkePFaTW8bKZ5xnk1VvZRWvg0DLzSUiZVrTW1YCxRtmJMIIpMPz22+ijh
RqaOlu4+y7dWWx2rk8CNYG7Zg8MHvf80sPtIJPRi/oA1wLYyzWGldrIa21f2zLPx
HrTJba4crFtlE5Qr3elPwPt2wuTbLHdUjR7q01nem5+m6OjXd3AJYAKyXhhbenQW
sfl/VtWepYy/zh5YHAMORuR2GUi64iqOxVBgYgLtGjEM64kD6Bm8v69kzND3WnqZ
qkGdPX2PsvIYTgzJO3pJ5FdLuiOXNyGQxd9hcgxD6Kva3o2Sv8Xk/jvnnGrCWHRx
yYkoFkY8tk697etTz+jn4wWj1iCPdKYJxfQNVy7oR4I8ddCSgjvlrAT2hxfsUnon
vqB/vn3Lp0JDPVaTrlDg+glJN9hYeS3BorPGKy6iNWNLMNbupa+hylF4J55uKauT
v10unSQcmMMaNsr5sUDonI18iMvhDT4DXnKO/u4SGpaONk+8AGCbQDidyoq+Rka5
eTMFFJlKZD5/aRsxayHRsBmWBojP3bAwQIS/ztRNvKNcYclBLuu5gjcEXBv57D2r
oWcLgEhbec0bZzEkEPVOA/Yia8HsjGhI+pF/Vbw4ihllRcMgM0EJTjwByPmeZDtJ
gZVGJrsEn7vEKJT/W4v7SWc9ciVTteUI7HNvAf7BSlI4uv1bS1Bi85bZ0M6pbq2P
drs4dnUklajQ3/mwxLyCKAPHGnaFDxJrGOB2Oyjf6Jlwbg5VFpXFgbylqJN6EFXw
pX7lTr/HRUn3YVaEYKmiYYcll6O8DGzJv0rNGGkG0j05r3lPEDPfdecgkOPigFP4
bnZ7MbMFr6xBq55fO6SCwXDDjPDdkorI+6NlCf+SIRkuIk2+wZ1PLy1aKX9PoV+z
AN+hqrFDYH72fmrKxxkA5vYRAynpfnLpolRJUpItSPKm/87TuoS5ZysvH6aoJMWX
M5072U2EGYBwJtHQX/sujmc+mbMOI5UoUGP6ItASN+YwcIQHRjEzF1JgM7ETIxw9
PWrkpb4ZCfe3N0+zWBSnsnEAwOjKXTPO09hggvyqhI7nGUYAjqYWK7nHN5lCN80a
T+zMulQxJonl/qPXDg/+eeTgccbw2G/jGjKV0nUZWjQkpTt0+TwK4Uw24QzXNl5H
sBXk+SuFzxKOHwWnc72P64raqixhrTG5KcJOgH4UtIfxNEE7fuFC2vVCjj4Cia9d
7ZSCMzWpfkW6N1EzmJJ5xO1p5yV/57joBAnus+LMaBq0woyFvNaqBUZiBR+hhzB8
IjIdkGcCLtyCE4p683yHFLxOOyarEVgzn/H1gwPxJ+TgYSrr5nKPIekEzuowMaDH
Po3DdzTpL81i7F3AgHMhcgkWt3ySuBg2wJHhOiqtQaIa6rCTswbcc4Y5ewh405Fi
3mW4WOqQkZJwseCUnr/GlgFgnNiCTgZcOOJGLTNksak5pSZ/3MxI/x0tFv6shYrZ
HCZ1cKGVE7VRpY5iPfFKzV+Q4GLIjC4WTUFRVeSvmWx0CkchhuKtKsoTzmhOCriK
L2bpa3LcRh7J61hiva/+lN41G/F3vGNLCRuDZXX1Jmu5wE/5BdoDwZGFyA2PrkRS
7qRlrzLiBGYFI15wAs7U+zYMY4jOV0PKSwBNX5XjVUyi0cvvAUU49JTJLykOBkJG
HjOGBzb8o3S8hhGTm5VZesO6j2EbMUSBTOUHXWllcYN4K4A3nB2//kHiB1PN0hsv
mjv00X1nOBXlJlIq9r2pMIcaahaoWlURNBy8V3r0olGIzk9NTpGGhV5SDyjrQ3TF
fBOoZ4YrOuJioF/9Zw22zwgH2ml31IwlUw5msddpgw1OqvDYL9RqR7JOn2lqip94
xPJdN4TmXljnMOxN5KyWMgClraEFgn8pc+/lWk+tZpFmdgnJ5/r13kfefsf6toTX
ITB0l9NENNynk7SNDxVj0mgC4hnWDaTY6GX3qWLF3fmmWVSLR82g+0eGVGtuh1yg
HoohY6kPYebmjV0Oo+XGk86OcucxDRdrdfSmA2ZSnljf6nkRXIyLrRiPR3v6a5O3
R75+Kr3SOlBoMwIfb6BcOWG34Y9c5OScyeQjSjHvVakafNERfbuWxHV47QjCf483
4906srjmiqNxBFFUZEW8pEAZ1yscP1swfYiSXsdUvTm3oSm0AonjWgddK2GuwRJN
WeIjoNy9oC4afo0tQs4LjI4x6zJBISLFe/6j86Uz2yIjlG/pXFC3Qad8Q0vZ69bh
HQ5yT5McSSO5I6bfJj9ryQi/LwLo3BVkSuEAOrghuYxdq5V0wGzBy6+CotjNLp7z
e9SWCh3QLbioX0YqNRNjjj+AmhKYDw9xJrwVZ7aNZQoOsCd3EOEOeo5kyg1V+++5
1y3AgqCqtKMuB/8N5tj523g0Mq7sagFA7ZWiX+7ewfAVhqez3xubC8j2OXF+hyt9
x8BFUYhCT4kdUzzZgFFoKALHilm0zOxwMS862Zs+prATXxtd10P4jbD2GAyeBM4W
LAnt8w6dsRFMiWpAgx5TnOG/SWxPPfeyaZP8z7fzoLkSNNY1FIzg+9d3BPzj9I3Z
EelSITkna/lYr2VUrJd7ifkqDk94dQO7EdBweu86l+GHFUih3Zop/D7zOvKBK8Z9
LUSofaF6NpO8S3Vp3OMV3lUHRxtNnoWBK9xEwRF7QBlgWFy2Gy+CwDISwpwbXMDr
/dPUopjddl6K39FhJuUe+K5/agN3jSSHk9MRvYLbIOEQ0QMiyDazEHnSKuSddvzl
cSzJuOiYmA68scLwv2qPtE9CsbM2nZaRnzNoDWgZyCtTvXlGFft3FrEptMMUaDrq
l675Zed3ArgUZY0/uGRoTI/AbqgpRpOytknSKIp7SKh16R3mW/h0oKFujZAwzbLR
WqlvvNgiPmRutUvyRBSbm3ApOSYp/SueYEeI+ATyeSKGTlNF31OnjCaE4cVNpBfU
d9cI4IPLtbFjA3ENBCMcX4UnCtpL+los8YDVPMlhXd6c21Mk3hfbClhrprlHQLTm
kTncnszxzjYEQ52E9pkOQhSi7JenDnLopH6r+4mWS7Ezz+0X980J0yyk95/M0TX0
FvOmO8mVnY1eHrWicoZOgQ==
`protect END_PROTECTED

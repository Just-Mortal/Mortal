`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DRkdV0zedc35GEICq281lUmCOyO62NtGrd6XscffJsz83r5W/qnqdo/Zbe0tW1uD
xtuTUhqKnBynkZa5oYpw6Xr2wLB+pVCxW0fClgCBdKVzIs91vGugQ6UYcS3fvv7x
YjzXhvSKEXtsg4tEivbtt7t4vUm4VjlpJ/yunYssIf3mV8fd3seMJvv3cyU0qFkF
YuuC4e3rU/WL9Pf7B5eZGwdPSl84ZoIa2y9fv/Olgk0bRWf93Za40nyzuZg5gals
vMWkfEAOJsJhgi9O7kOHzQyNwG+lFlJJh7N42IkXxU38V+ieOkDo1r8hyamdqjKm
v8bijkKIFB3e/OiZ4VKrG/dhhUF/cZEtTolNd5MOOMAAUx5iameRGjJtMUR1hRy8
IvqYXtTUeLEnFynyygwBz2KfdQbKLH8uOGDjsPl4u3vAHr3MO61S0ShS4M1Uupsr
gqJ6/IKzLltgTFhLYBV3uUbac7MdMkqqSx0XIA5mChruDIrWkROrCr8aewoiWywa
EVz8xlwh+jgNCp8y6klAdGEHfrox3yzgJEuFDTleLGQYq0h7vnVJRgCc4Oq6J2YW
M0TbrXG0sNHWaLx1s6RpSaQtTgXH8903hOf/6Y25K+LbLsvOPU9lI8tEe/rKAh5Y
GokEBieeA/Wqe8WRbXZgkRbCeXpS+Pa7ue4LNCSU3qB0giIXl9VBIntM8FBFVrgK
Q0CqJbVLTgOFHYlNxkNK+AdLAul1DF3vlw+NiV1JhAuUuPP615q5i6Ip4iDD3da5
GiFeEPP/iGwENPK24p1AChrezPnqPDmkqs7d7hRycCXDGsrkQt/J7OS4Fh04yCMg
on30Hzzec6pS8/dQ9Q7wgyzEJGuNaxeg214VI68sg8gXOnKQbuVHISiMyBgfraOS
78FlW/OkXc8oBMzxMir4yoy9rZvRRzXA5Ci6GDNlQJtOa3cCzihSUs0k3QkH5gPR
BVPkdI/p0at9EBrxkNLKCxMSZzLkzGffXycSbMRDfiz+aPz0mduBLJ/6+/WEWkOu
JClzd4dsZvUNSN2Q2Uf5/Y7BgkfZ3jk3sOwQvOrc5NxdO+FVqK1OVusmnHAel7s+
6rpzWufwYHHTDl8qBq0/riE5GlDgwJfg89zcQntm6+QgTUl76zzlh8wOAWe7L2YD
bJQorH2eRUmxzhhhCoIFu11bpUd4WsJroeKI+YGriG41p6QpeYBbwJqG8oX/JJW+
KxK+5Y8k5R4lGRHb7t3qvuQ5M4mX2UDhOMrMH5qTVNvVRVcr81zwooVyzgPnfpaY
lL0gDca7kbzE1slHxJ+LfM9nnjn0XBQBzfKzwdMPk2dA70eD7esmbna9VQdSShTf
`protect END_PROTECTED

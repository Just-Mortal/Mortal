`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gqHY0uH12vgb56L2ZtsJasSB8u46VBUmc+SfCP7ws67ZGr9OAJnNvSqcV4Z8Mg3
huBaL4aOdKqoaAJ9hdX3oZyIuOEvCBhVGqlfzrqPc8WE/PsOG4AsKtpxaPyIpmsl
IK3ZQkYdJ0QrthymzvYGGw7Dax+S8ExDO019ogBKDQSouTEKPbdU60TVsHjEeo4j
rnvaorF+ZQ2FdCPEc8HTXbK9LJmMGlVABoYOGqWBV8fx4WEz8gL4jAXCYpFQ0XDO
rSRZbbuNZjEIsfq9mJNpKuc9R4T9biGPL2Krrregzx1Q2OABHmP88RnHPFXB30x2
z0Mkzu7Bgp5islMvsjHMkg==
`protect END_PROTECTED

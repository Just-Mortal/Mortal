`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R8LJwnpcqkrKjngqI+nMH9BVU8b5mOyr0NE4/MrPvOVRbWq0YhZF1LAIPCdoXogH
/Gusv8WVjiOHSRF/b8+ZlRV0dc3q4/NTCmwhME98DDZAQGM/SsAjgFaSDaSj5SwP
qnNKdXknd+uA6Nk9wgxQaQYXpcL1QbWdcEp6dvh6je5FGxEGGQShYipyr3u3WTH4
XSa3tkfqKi0PISULOo6WF7PUzny3GrIIQOniUYwANBaSoAtbV92WjhgTZXmsfujM
3HudC2ipyldhB4nDt4G2Zcf1ZSca2xZDGuhHbTBvxUZ2Ay0rEvswj5FdUF3TE8XC
6WPpiom2rycCZ9sDzergH4noJBJhbtGflo3bBIBuEllwC2h24y6k3MweQ2+qE1D/
IKRcSQ4Rmo9oLO2LOoDhAzRfP9y4nWk3FJzlBy4yrXjODLIYdE1Pykz/1xYxPbx5
w+X4NlvdqCorz8L+mqdzIsZ5rYK/aWWohcuZjPD/FZu82lCoNVco4RvVJJNuqa4z
tP6UfP5Y8VzBoINtpzVVuMMF3767wDY1iPAYbzd7/wVNUdWePohLIIP7eSHiDOgS
9zEcnCwuCudA09AOMGtHUECTXzLXqHq3EtJLzIZoqc0vh7A/bimF6imKXz3cjWxh
U9KjoX2bkhCDGPttS04cF04xAQlQQIlJ2baUZgZ8dEhzBaeTSB4twAq96CUqLh6J
iOTI0u88Epk3SpGc8iVdWcuMCi0GHXn6rIswuFbcD8/s23q4bX7OT9OvPOJ0n3Gl
NpYHuNnfzorLPWtuj2DRnZDmxVl0nGAcaXdThxK+BgTmnMNxeFUAueAR24wrUvqG
W183I1VYvxdyUSAwqpGJbKJcMj+eh0F5dauFAJ2c2GMsSHu1rz/dk+dSg7nfC0Xq
jtqrCFczrQ5ftQG+644IYGyZ6tQmgaZI4BU9KVTkefVtzaktSL+3IWdq1AGCtpPB
QVq+FA4XbUsIDugIMVSz0DcXrMqfe5obIDGKCBONyla3W3yshcuDu2Tykp0MJq4g
F60Gy2KjNvn1ICjTqFxh80T7k1DAQiQxtp5rBZcGWcc23VGAl2PTQE/6LrZH+/vB
JrbVdsBvLSGjqZt2M82RYinYYvbpPSgEQuHsYoOJhGWiCISwpZAyD+gZJx1o3oni
zMStyj+3imht4uRgJpso69j5ZfW1EVIq5jV8rJfvkrexrEzVeDseSEfojW6Jgw00
uck+btWcPYQyUH1gc5YQkaZinIrSdWIP+8MHMH7KGTHXsCO2AxhGuXjIgGNV+Mb0
4WhpYbSJ9p67dpGC8q7DMHnH5fr/HEAxytZ0hvxdyLjkcBD7C7RIi4Ft+6M/AFRw
/9BLEDrFRzAyZe9q+f87C76iCC4Li6m9oS5PyIcU4tir7UWtGY6+ncsqnkcbWeMU
mu7uYTRZfSBDq3mbJ2QI4yQc3XE8f8D56C8aEeKnWub/6elefeuoPGg/Axo8coGl
/+OCA3fX6oZarR/cGm+ob97SRHNlAcC0Nerg3TJS+v7JbuMRdobkw7J+OdgwoAe8
PBbi8rlTpNAnjLa7pWzR4iz4Opm4G1fjGAl5Y0WI+MdxMAr6lJanp0a9YmO2Lv4r
t1Kl4LlALLtjoHBmDnrnFMcqjbgReyCxyrPVoXpePZriwmjhuN6dlHP2snxRDZFv
RshX3xOR9oq5lLb/6PI75DU6NGPf0NHrFNj0LEWAYs3O3K9xUXJwzIEEkCgxNpbJ
0LFNq0OjRyeXGsdM4ikcRFzxQRDIU/zjAgwo4vs3qhiwbBiRDMZGmP85jZMO62td
ec8LOg74fCeGO45+hvCNHTUmSaD8x+hS2ZD6q0xYs0KCq2hQ/Pub5QhIvXrbonuk
BHeuKAgjIa4tjOTWcPNyQRC8vXxuNWBxH/FYXRsi4IMm/7RtlYWcrZQWBJKuvNjZ
BMuIM+lRc0BUETmegBXL6ki64YPJ42LcEobU8Ht9taUsXSqlvnvOV9VpfNqjr1G/
MlxXBlTw/og9HQ0alOClTGl7CbVd9zIIRYfXph4dl+yUNdQ1kmlwIeaouK4Hu6Rh
s2ymHEUR4nzOnkzMqjPny/fFgMWxiQ9E3D8ftcCQmFoCp28vag7CZpTuuHiy/b+w
jzLFty6otW15o7PBwD1b/RBfEwaQwnG3WtoeWMT4c9owXYu2GYvH2vq0/2y9qEmD
llefPBxFqdtDWDyWHaqG/fH+zkwM6I4gLSbliXW1EqQmSofw7HJrOFpttYwf375t
6yGyRVeE++fOSBB+Ipc0HKZi8QHwtyWT9gTtetD1IX3shxeUnqjcKitlMnprnWuw
2Phqs12BVwOzuJp5UYQSQafgd/TfB35itNG8VNXTGhoma9vFI0eSF9BwvHxHIcwR
jEJCH8L6H8TojQQt0THfd3pGfxhBfrNqS3jLvSb29CU35PXxsjd2/EEoo/vSgJV8
dCOVUkLmf5dLZ2/NiQyINNcoFNX/sdITE94IgLiz4QCE9AegVjcbE1XaMFboWiVJ
P8tdrb3EXGLrQk0GjvLVVXsZVko5qWC8MitU/wIQEkl0iCOpOl0BKKRP/Dmc1BUd
EoQPnMeO3foCBFPiv2KwTYAW+c/7nXJ4iMDpL7F8NyAy1A/8IZmzvS2a13RYxRMn
k8tRi2AB/v9bGUqNataHaFX2hDblVzZVd4Ihbio3b8L4Mnb3dx59PlfKVB2pT+hP
3IL3C+PKaJL/H/LyFODtAfIcaN4XnhJY2jFrTJaHdEUdSxWMnwVcAMbgnlB1AQ60
NoB/kvQimReO2kuQOAb5msbH9qt1Tq6p5W9nV9AnoroD1xkNn24sVQ0OEBWmVHAy
wB1cX9Opf1DZHXAZBXsbfcuI/Ll6yYN+5eJmskx3DsjMm2h54IVBWCW83kSZxDAs
uWj/vBSzJrV+RgHQ0ZoipphXrAvcu5ykPPu9qBmy4c+xm592qt2VR3ES+ZvUq5tf
cqGKyI1Mrxq1Pwz2aakuOkqV0hbJOniRBapkBXXfXmFrDmCI1iFMsq5jhQGKSQCo
+ARm0UThZLvSjmNyBF1F+2mmKcRXdHF4ORLaCNSYWbw/H3BkJial+bImz7m6W3nT
EIRveojc9r7CPn4Hub5Ni0iLx2cXq5dGqC33jBzxIw5isKvTLZTDnubauFgF7Ke0
pXedrDCSJS/ltt3XdO92cZfzBer1N+QwgveETmUaLJQo1yaOYrw1/+nJHcUmrgsg
v0ReoE0+27eztc0cfaQvHAt9+O9wywCcdNioKtvccf+N9AzdZPAddDBvCXJffxBX
JIqJUefAAP2SeXcLFZ6Wn1aN1dELDoBRhejK6dWETuC3bMElSkorCefiw+wIg9/D
/zV3Mvaw4nSHCZ4fTMYhu8iS/PEQRa45aHzd+vEXpW05b4+7Z4oDfSkulufiHXd4
1aIeqLmpuePSkheRCZ1f3fiiNRDM1MVsumrKkjsYiETOsvKi/OIc30Cu5SY4WaSX
aEF0T6bbkK+2dt9MDyRDox8qVKO1v4uTcd8TzOMlwSU37+KU0E24S+cR9Q6y0AAq
vplfFY9JPNlKI5POgCWRrIAmtEPRemID1KFJ+eJeLUa5RVV9QKc7edlFyf7Co/Am
FOGiibkL4QSK2NAQoy6lBNqYf4Ar/Exu+1Mq/VsiKY17RpNaqep64PKulvzt56l3
G/3e7bC3Lk/16xnWbVoVeOiRUjy2jUtHHfZJOGn3E8vFtpf+IiMocvSNEVDuVXbX
64vKz4UKvIMKMOXmVgOW+bPBsRKHTovpE67iHunU8ghvs8b/1lvSnJ0wGwgz7WbT
YYpqOzMIoRCM/fLp4TIYx/eL845DQUFPRaNol0Y3rsdRggM5fGePK4VnHG4fmRcw
7dWXpnlu0zy9Y8+c3I6n31TuVL+Vp5G4yVRT0R7544S0jw44l4mwjC2NDcWUKm3y
y2VJXsUSH1Nbvlf4oTF7inoaKqOkx0IOa81LQNTkkhPFLBdmPdOvUgSwyHXAnKRw
SIk8NI9NRZPZNreSVtcXGVp5JTghAT407MGagN3yNsccfJtIHQiQplU7iMg+FbaN
IMYyMNpWEqyyIVb4ulrnewf20U8UrpXiGxL9u+vET2xTkDR1eoHI1LjPuFl6nbiJ
lIEplOU/aQQ8Hp9S5v1t2U6jxXXKl2cUF8ddAU0t2Tz5nPfGY3CkLjQ6AfH6bNVX
4OETyDA6up9nNuHFCMTPVAIglB9fKt339KRnWm8xu4yyuJ09r/AGIiuz3XnP9Z3b
A3+SMXvfqeFdYcT44Lj3dN7RZPy/iBuZmreYUogcKyFMcBu4G0D3+wGWLMLXMxgN
OYcQax8sdD8wTYg8Rij1lIqFnElMenKtk/yHf25p9Z7mX14WribFdS4EzF6JwgEq
ZHhnoK/sQdtsYvcQ71bdr6lfoCHnBxvmlU85uCI7EhcW2J0Xi7hTm5eLKDaH1umo
AOuGWrjmwIyf75p8G4HlhKGLbeRbDO9zHWcZXgXuIsMMD30xW4GhJTq0nuekC1AQ
R2e6/yQsJVrTGkFG91YL3eUQNaYAbRaVl4hto6mwyNJt/CEKonfr9dbUlW2LOp5I
vUP1hXra+vM+6oCfSvlVSjRIjIMt746Jki6G0x5qtXGcMTUsps3YfSS+WuJ9O1Gh
NtQBaG5AQmdauVcsnRg0iwDpoWucHI1fGzFsU/Nh+i/H7htorOsNHJHxEpqlIKrp
tr5lCWs81dDW35B0x35TQc5ea6Z20EcLBcAxVxru1c0eG9vqdry8H+AllMggIt6R
6PpkId8UtVvjsTuvRwFfAoItQAUvCn+u7+AgUZPLI5PQkr8R6xInRFHu06jeP+kp
tv77CVhO7+fG0V9HeKUNIfkfbNiC/o5IwmRg050dM6DB8w4EPtgS94nLR+3LFjJ+
UbezZRCM5bh9Yud9ZsLuY0U/pXZXS7khv47+bJTz11midWHi7/XDR2SIkx1c5uBh
ZzItwYWuw+TdVzaFYUOwrWgd997xtF0tGJGIM/5qq0UnhTE52ihi6aJ+YppzERr1
22Dgz05LrdsJWT7FCKmFzLdMDKHsAKLiOzBUTGxNeAcqCTjKHV2LGDcHBaccduQK
wqZWLzXXXtugSLHs/iCL/SM98Ex/JyAG6u2e9AkqhXYht3TtjzrXPsA6WgZW919p
2dnxxGTgtOZp56hdSgGFj7l5hGvizo0t598Rr+2lG8oa0azj2UVtYTBM/uHP7nZh
NLSeq3yosl5BfUokFXXk5kgShMlWhu54jhjHjLCEsnHEqreNamHAEV3V++dasupR
2mgkW/od8oCSH3JMzlxDuDhpLZjaS9IB98lsFKXTw4Pwg5cPlobJ18LKXB0I60TA
ebgT3aycxE9tVTHqGJZCyCXtEv+/NiepP3kjnEle/nI2B+69dtdK6BI1F5+a2MXx
+qDc8XJ2GKvnr2u5YkwbP5EU/FJiOEsTU37KLKIXa9bwZBtowKTyXHoUBboDgvud
erRXYWl9XL2QCXTwb1b6yYzcYKspmCtALrKF24ffOH3P9J9aAt+/C+rrclQM7pn/
Ml7rBoPvZwag7CZJGWB3KMtrdHS/CibSjp73PoEhAYf1rhCZu0i/rWZ86nxtnK9j
q3GDCN+0e6Z3lT7/gQlY2srZIA0XccIgQpAgZTrfbmp4jygN2ctjvNIQ5EiqRYuP
PliyKc4LTNa/Ky679y/pK4u6YP4kX66suYNyY+xWC5K8QRS8oe/7ts3PJAPyT0kI
72nvD0GNvBVCWQA+OuGwWhbRb+zRCSH6JnycQZlNVItjZamcFxUkhZOtRErNJ0lY
3ClHp9Pks9M70rbALfTQ5AKfNQfRglbQQdhkkdNG1FCsQbvPWlzrri78JicITYaf
UsybV0u674NIl+ND8dJ5Ed+cIZwqMJuCOHg821dozSTV8ZQxq5D69Hr2bH9+TO8B
EtIWrR/xoAVRq1oLiPY3nDgfKlAv/dewVTVOS521LfA8nzGjZ8QetEAg4CCmGQtA
8rRB6DMu+2JLMO45NwS2HeQB1UrSdKpRYSxoKrZFB31d/n//luw8ilXMyLJS0CWv
mW/VAc2PG47AIrc5L6HAXLsV1gJ2YQw9Xbn0uMpq9I5WPhxC80LHnMortRgssG73
qS2fLM+vfvP/drywxoSvqZi/HqEmExEzoZzwU6+Bk3oOaUUvvtcPl7RGGsS1ujXs
gdH/2Diy/b7Lo/kQqgmEfU3ZCP0Y8m7ZFP1d4L63CTEVChElgOYKWz/v3gTS6t2C
Pv7y/b+Tark2gZrzUeG9U25ikbeWAUNCoP5HK5YoB8cqI3vUF18b/mgTVO6ckCuh
mAovWe6+NcwjJk1PcA7RDBZUH6qxCQuaVtfYZtWMgnxaPV4gKtV311C4IxDLcqXw
F169zMIOK+nlN0htWkFwt2C0iCohNNz8PmqRIENVT5mY+SAAC1ig/URPBBVQXGwK
g7xHR1OWBfj08OAIzBiwPe7xF6W3WcGtdTdT0zsxb9IW9vvGY3Vom/bowaFXWZhz
thZv2XQmXdnxJM24jn2JW3AiAP659mC3DopaqEODtAwcuE87NOoBXcKJwX9Re3YG
WkgOQqJ2WOhAy31c97Lz28qo94af3NSRhtz25fgSwz2qPoKUzRDXPAQS4N6Y0BHc
Bh+ZUW1unMZStB9kmgdvdJIk4+zYCuxPuPlo3VEN9TcZBXWhplINrnNULRNd9D5k
pnb+ZgFK2Ijhe1TbMia85jlyI476da2+dZwGs1cHN0hg4A1uQ/oIX5Jb+Fe7oXqW
VTe9walVarHhhSU3IxfFHrKdFcn8njIetHGLHx2G5j/L9eelwunpUp47aKjLIVfE
KCmaDULwQjLO2k+IYhFTTggMkgTFIrOISRswe11+0zwEs1LBJtJGs+J6KzpQjodG
`protect END_PROTECTED

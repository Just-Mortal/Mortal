`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TW0hg1xfD3JI3l6As21lA92GgHD808cOtR/iRdI3lwZAgiKxhpGHrKzXlQH4DXy0
H7H2eEjRWhAs7qkzgliD6flR2B3MxYkdEEqZUNDZhNK1KqGNfdk/xnQ4LX+Bg7Vw
KE9HGIxx22ZIiojBqEDF9poGmZPSsKZrdXH63RKrDyJCQSSR8ssRH+JT8M11p3Zg
/uQySuuWTTy+8FnMPdZM5Fl9Icrr6lm8fT8F9dMpu9bzANeaSijXm3J73wwEEIlM
05hIiisYV834kO05tX8hBNlP7H5OGoDa06RXPqmqMRPC72xaLirj8TEYKiOgYzq6
rAK8L+n6GP3ZcZ3dvRFrCzNlk+zgtgyvFs+fMoNctlNGO4fPNcPcv9W6kSKYMHuK
UQ4rxnaV+t2UvWKAmrwqQmDghq+7o33R0Out/wvDCM9F/i0+Jwoma6OqCglj/ACV
TPFZHNp+Ba1ifFk27xBVEfrW6Hjy3uwpIFg6S415+dZqM1gEO0JyQAPg8NI2JO2L
nyEBgaR3e1u6miKKkj7VHctkP7u0buvo4Dut9S9sDA55jz+h6AT4/O7Ousa0yMoT
QdFFxfl+i5Nl92Wx1o2h5EIKWK9ebuuYQKjx35LCTomAo/rHpdQTFyHqx+ww8C5m
qAyM7wXHJx3zoDCoOUkOX8GifgLt6dxuB1CuUMW5CxB5YQm9RnySW6E7ftdUr23S
`protect END_PROTECTED

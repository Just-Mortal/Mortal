`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwLo+aOjqtJKiCS0ulME0DQ8Bzw5zdFYw6Q86C3oMZ8ZiAsZ99XEuFRMD8eZxcDe
TZ98NpdRuqsfpFvVSvQoF43Fw2K8cQiJwVtvaiy0ic8srf2oZqEZ/tBEle3yg7bn
GB5mtvMVt6aP9duv8HqlcJO2jhmLDTj70y5SNGHrY46LyMO9vQzcrU2L63xyyIR6
dBJbcRx7djDaMwmSG5sq8CkJUuUFVacBdPrh1WEmtcEe8PLyvr55z0449tLSqZ+Z
7Xc1oouoyNr28CaZsUUppXcYchB4YczUzEKW9LuJgncx8A6yI7wN9CPCvkXyM3VU
vmourS1JEM4T/+gem4s07NSItIRtrsOKhdoI0rxUrL6YVw6jMoxLy7P0QFC3n8zZ
rfeZEQZuT/RhY6GjzwHlig7Vml+TbXesW/I7WUTZCXvasct0AhdDKMPRkpLt6e58
0ju0KS6R0xFO+UQDRf3IqH7EW6ROJXqg0yn/3YkPYMHzgw7AmRQN7rj6gweeHOY4
Ahb5Xf61OIXGyla2/5iQ46E2fkSnO3TPdi+A7383RjibKJV/gq1mX/EnlH3ySq+0
qJ02ZVX56f2fICDdGT2sKYcsXd9aH9OtaYtFpWwkhMd2oWlKqj60lcbNF6z0S2J4
eIkzwR6Lrveqe5G35KAH6OmZ8Bfv55XRdidtSa19aGymJo354Ny5njUlZbFcx/3D
QYyUkAiAslPUQIEdFCB5mYDtCKUPngdzE0cW+C37asTjJO9Rg+0xldUf+G9/CihU
/Lh98fI7Ei1ii9tciMqT/9INtCQYH/6FJ+l268SE0DCp91L163gvfzVctNxsSqDt
cqHusXha5JXgBOI8lu54dFi+8WJGP+u9QIF3pPKCEVUTNRkMKhfZFfL4SXYdf99c
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0OKPxZj2g8e9Ban6E+jro16rjR9VFWx3lPT2pJbEnXZ7YdvjL8WOhCAul2LWxHu
F++Afh1qopCQlJfuFPEhT/9i5bS8AqMrx5QYpsE+VG50bWYqwjsoV1jxHyig7TnU
5ay+lLtpYiFrkWKgXMbJLomLIbemS7yHRmryYZAQE+qKmYOGxECc/dNMooOFdqfc
mPCN1sDdaEKbwlKduVKjgVLeN+saGwLcJYNdoUzG+zhD/OfY8T2dQdFjEffEt/Qr
pymEBByAA7f0jrZcvPDmQ0tIfzBmmRWU3L6CW3mfg0NdnV8r0V2MHxDk1THZNwwK
HeN6yiWvuyn/ef6Qb9Dd++/1/lNcBOOJH3WYz47ft5I7J8t/FyQ6OmHt+phQ1T9j
y/crQPpSJ3lQZH7f3erSWahn3wKTSiWKDcVhxsknYyh+XAi8Ai2tCTWgs+AQ8sT+
BVj+4zW9CW9ZyNnMcdSUNRKqR5wHnSp5GORx0ztfGA4pZf2UwkqwneCvxApe7RZ8
tpY8tk3e0DsrJjK2xPmjVQasSutj4cvsvhWIjvZa0bjb8u3Ktpa+VCoQLj76Qyit
NJVG8po1bJtdmg+mevanLNJxk6ZKIMW/CTbBa/I/jRvDAda/v1dVWFj7lucn3VK7
PzquPvWl4ovrAdN5g4QwCxCzvBNExxSSx4Vu8gOyuj5cl1F7JBqQu+ahNyj5LK8x
oDL/wBy3VH1Nhn9RZRXlcQLjAQMFQes/9STWAUoD4pZgZhjWdRINXlwfD6/X1AJ9
y48ezEjeBtv9uQJ2UBr391iWth2N0g+I6JBlGNbyemhzNWIl91NlwfObnGozvoQ8
dsFbdcDEInTgaQ2NCgO51A==
`protect END_PROTECTED

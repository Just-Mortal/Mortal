`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68IKDFjuI0okHhdDdfsXH5WSrnBawAuYXgXedEoQsoamZlVBIy5PACvFA6f70WKv
l8MXMa/HdOL5ARFFmyHwD8FlQF3uD46ChqrNPwTJCrml0adQT6HLjijmACPM2Q4H
0TjIfwb4XwWpVkH/hEH1dCz1w2WEpI6Pg2deKI/Ws6AFYjhq7IvXV1kzwzgbC2Oy
xwTwi11ksKnzTmJ9wIXGPzTroI4aX95JgGuIN16h3899TDtIAP8BTmyqDlzuMC0E
3LtPBjqQPpRQ8AKtUBwmxUBHO7T3dXOZRpGQuWJrqBHrq4ZrpDAvTnDb5bjCL8qO
Rv11DLW0j3Db5TS1ikneGkgxXqFQbMQhxDrhm2kyZPv7Rlpk4plT6uvoqNKPH1SO
SSpPBtWOdDpPw0ZQQKlzlIExfl2N6YENX4rT8sUsTaXDRM5AkrV6RoqtvRD4L1h7
Iy1aoURw+F/vfQovG09Q3nQsa1dGHOYQ5p1e3oGX9VCDa9Or2mxajfSer4yZrmys
qx33vFMuX1Mf38guGDj+1ZbmVlQFjNAboTrharteCPQyIIu6uaTfFDuIVEu0Ioek
PvA9SsmCj3/S4k+x/PqmWoZbedzP8qzTBPe+cFms2u5O69eoVtrCndHFLZYxVcdJ
fI+SME0FC87iEaHca6mDE3L/GQebSX35utoUyGxOo14rE+28848AMrlUOQMbwXhH
YGKnb5lzE5uGtgTOrSmxfkYzToJukTbk8EceMQJPY0NjJ8X25FytX8JZJKCqJ5C0
e2KBZeXx+UiegXRoSOJJZHnOqkLjaZxTMa167RqaEqKWSxcd5HT355az4xSvqOfE
ZE0a6PQC3UFDfi/u+ApTawHueJN92IXNedjCIRJd4PAVAG105Qz5T1qk8gc7tFSQ
AXnN5GyeUQP1DV71AZDOi5kkuRxq3v+9NfJfokQ5YHX/HQsrhGGck/maGA4Fym1I
aba3zW0++cFwhIVzeq9KlemqvThY9mwFUlWYTn+7+nfdlJueY0yqxXCjiQSp9O2V
RujjEhijGDFg9rC1uhZxCGpEUz2d+59EHnp48AkR2DZCtuaChgPvu3Gk/Q/UHNsC
FTR1flx6lzz74ERY0HK12Iieci0STc8jYC3qZ9eT3whdjd8LfRvOhweD+GDSWxlH
MSG46KsQz53eCTcRtuBN0JE4l4D732lGhXMG0hiXG9JBzH+0KPgEcz436Dt6sY49
+AHj9qQOa3Lko1mSHpOX2lBNA+V65jYkp1FpzHrH4Hgc8+JI2VMFPwmIvsEp/3FD
xU1Cw3BMGM99bn+KncZDIj6/hjyHmDROe3n6XSKOtGgx9J/3AvetWFD5UBZusGrj
srhRqb0bpU4YRtYWmjD/BJWLvYrEioWmzKEgAEyk3fva8gs5aZ85dvlxEwje7CZf
0NUa8Ow9GZR1GQG/nSk5h2t5i9wvE3sJMN8q9WH0jO8EPPLoFXXk6dLdI5cRgzKQ
tzBUS6fKpQNgX8lypei+I8oiajQiwOiln5TWScSHr0CK9rEQVtfe/rOyXQgiyKAo
q6hw38hCoyhcpDQen8ZF9vJBGdtA/dqbr3d+GRfPXk9DFWUDdSYESwJ7jPIEc9b6
I6LQUFZomuzoL/cJWiCg1jOW+Cy9P5c6YHSvREvkWAaJHRuLuth7XfTJOgoCKLWE
2nmO/f71k+6o6N6zhroynRzB3QSOBSwGOu2DUv3/PGMhFie7vQpM7/a1uJQosuPT
5jPkCeowgUODjSBdWyHvW7ZxqU9QG44vdDWR/PY5SuSkCkuR7sLcEb+q1D1I2X0i
ABaW/c9TBCr8qu6o54eW30to0QwBv2odS+e4uf9ycBfc2s7PMN+NGbfPoU+jQUmb
Lj96bd+YuOalxo49cnqem+du0ZwHVA2LOmwcJLmcZK8c21BUmRUQzzzvKX0wMQjp
gjLu2U1/KVMpY6F6ZqAxr/M7RzTvjUdjC3VYiTqwrfpkXX01eqHBXBjIcVXQ93eK
m2crdoA2/O1C2EGoBxTxODCmj04kWwsD7vZQ/CLNvoWOIjvSfVrD5QYS/cKlxNK7
G5QpOtqka1LyuqehUUPNKrB28TT2lRTp2zmQuJgCKMeA81vxs6mfN2gW2lnYkmUX
5jLCV8gX5z/EW8zvLCcHuK7svgKx/MCbyOYZhu9kprOjpxNKNjoZABKYgKrltH97
fwGqL3DbmmIXBwlStWmGddgYDIbbSZNt+4twm6ayo5KAfBAbKXbi8WcgqxxWekGC
jqWuect69l2dcXzgh8/3EKB8E/G2jOCIKgGFGUaxAMwnWMuIs46qwM2txhkVeTrZ
I09VYfRDhPZWEjZJVdbQW+fPmWRqW74khkYTjfy+nCSujv1snrc3LaVy4NAoS8Ox
Pk4I4cyoTnDel8VuJwpd7RcauuZzBGKr+M+pR75eC0mJxx3UH0eKfh9aYmZp+Qp1
fEtSWp37a2mufLZ0PhanBc0hs3Ytj/xJAKpePpdrv0wGv9j/ayvHh8eGSsLD8xKe
5nV8tJZVdcIu9TqKbh1OQQo6Zmwq/u29H7+nCHLTjXOFUZm+qUrvaaiRvJN9Ok42
w7AkkYY2TifZCxJP5V/GPegLl4P+AiTKnqN26vWlxSzdez+gAkfwOyxlWaAq1MgQ
oX9D9rFlOPkNwkmTMFiRT45FHQOf0a7QOGFWdJa1WVLqSKeCGrtKmEOUPvj39arv
RB0HXYeKFwHwKPDU3Tl2pO6xN3Y4IjB7fj8g4BOdUALh7G3vWEIcc5v/TCd3z7tH
NvpwLNuUeiq533t/o0mTzlC1gZ0LMl9iBrcVjXmRs7sjj+oMELcdupFBNqzl6GVj
EcQ7IRqBU6eOqCvAF4UKU0SS0DrTgf0ht9Vn95WdX/wfROJgJcYovL3JaTJQ5VRl
uYWbp4wzoWkpzjw3UslWtpHASNjPn0u007ggirS/xf2Xq+ghwX9vBoc6mdOphx8s
fDl4rznTJ/IJ/zrRMHCYQeDRiHWxEtkYGCeW6H9ycOGSxYePWQndFoWS8/YY+c/1
WHDflY0O8SsMm4WWiGR4emLLv+k7LBDT31Rj1Sxvt6rAztCGbyzq0qFAnJcyR2Sb
2aN2DU3g9ydhtBojtkHK4e5/z6UFXNUYn8oTtD5ZsTfgPevr7LzsLpnLnCYI0yJE
nsP+dne56/Yk7PY9bmBjyZnSh4Qm/vhIcP1mFOpwsa4KoINgcHmnt2jkgWP9a6iW
6Yeibvv5Hz8GuEz2QbrtOYixKKOFw0eH1FCYXxNCiXs6q8x7OIRYAtJHssgn7rhg
Ywmui1ofnNNgCFboUoiP8NIJhgKOB0FvEG1UOzBDYazGnuDmBC0YIXmzAKh5b5vR
wJvTnVcz0S5ClOAMDIuy8lzC31QEXtxTcRh2++SEi6CSLYMeay4a3gGaqhazGUQY
AN/vTXNH8gq3Vb3PA/2DhOkNljof8G9JzHvt4j0PeA3C4yeUCryPI1upzyfyDFD/
suFuqXi2HHuy79MOmVx/+7vD9SlfEkTZJjLu1tGzAfYcIxRb3LOK6zM4ApzSN/1x
EuqAF+m1lEk74QnN7/DoY4EtoYqN6B9iY9xgpB3OwoQsaWCtqa7Go8TJZYWsqABa
0E5OS107ylNaRrOq1xWlzO8MZ8nA0FlGOCWnDvxOCODVxSwCNCjkhVROkLpl9/XJ
8+wJAALcRb/rvaGoSUDrIlhDROkwcNKFrJenMN/wos/20Jq4oMox2EhfrKbYHICB
I5hYLDFeFHLUCY0EoEdp6vkZsXz7fGNzveKMRsTm/BG9IjsufE8vNQYdtWZmPzDg
cnb6pt2P0xM6M9v5IXMU/YPyC54Fnd1b+EX+8SvN7CHEX+IlxdDGbFGV9o1DLYH9
SBCZubjtI9KnpeYeWFhqsztV9sSiWlOg5CEQ/d9l/9aHXK3p3zPnBJsCnVtGBtj0
mH7SCExcX6qkDQxVldFSKMIbkyL5HrPoqAvO8pFprESktbwsUbN0FZWWWkmGNamA
JajS/fYfq+FcbCYK1BBRsPtfxBcxmpOIa8Rvtja4L8qYLSCcc0pQFg1TanUeOzB4
sbj38vozRhUwBUO7gyg4zTPBNFNoARBe1hyA1tNRZBxj0+5LcwxC8ukyjunG2m7z
eJ0rDIaXm4neL3NqJMLN5S/bSddEZ3fITQA5678ozhxsEeZcLDe4/zWGhubOMSj8
2CPTOkduFJK9I0QZLJghre85ELsbbeXjom83MqJXz+sbFMUmN3FRPbs7ehFLCFrL
UBy8rD9BzWwadko2OZmzh8dKwqfye5mGWhR/Zi0l9vNTrPPJAl8WUxH6YBtHgFzv
Ms7pcu9TeWDaqbJkJv26ys0Qc0E95sCib/57BtJa+tsifAhkxZdARX1dMMSUmTsT
7INJCvPqXbnvzU0GuoDg10mvaO/eHgqfNq0JsEajKAkW314Vhtvbce8q1sye8ybV
gt0f/R2FOqhU7x+wz+XeO9gQ4BygI6Jtoy4vjjUNO5wP7KOeq8i7HhCcIamT/vnN
vQv+Q1SB8m3TA9l/lXTIJNiePep+8NcKglzeSja+3VkvT4C0+uO5qJ9G8WOHyCGG
07ZhPFONtJgYt3ktR84htm+Ca34cS25ogScrSLJgCuUSgXXfpuPb+69Jm2q1jFKr
GRsbVZlIlUDmNke2hUE0hwVwB9cB3li2Zwqf0B/2qFv6yq9suasrqDwFr04sKIRl
ZCHHXn91kTL8mX+GiH8fH0S4zWI5AfDssUHNxaLtb/zxI+lm4oMZzT58XjnVv0t/
4NPFecvGjpbF+e6CXVe7/NrkbaZnTMrerieRC/TD/0iswOuw9WlFjJiDWcacfjuJ
n8rTmaNpPG0vhZjvy38D6tgO1v7VGWPnmmpRGT/NdEaPggcKtNaeT1uIWv1IOcju
WyUc7GHR6I1N1Npn1jWStGAEzyUlG4OQjS1x68F8P2CTZsSlgfL3zZng7pDIbrKo
eeVwS6uowiN6GXJaQ4a7+mmWM5He2Vauo7hNTyBnzAL4vqi2YaXl34nJnZh4790P
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GgZbZr6OefRVC3ViQYMbUXXuVc44ybE9VbJ2khHjjEsR2U1uCtLAcrwqHEZ0sFnO
72ADVg5kteEzq05Yl47DT5TR1+tz1VTd6MsaU3g8CQnaIGWB9QqzOu51wG4yUfzR
ejeda9M8Pnday9PnsMnliOoc0k47IuW7UJ655to/0nirMlFMc+rnQWuQesBd19/M
GyPtD6OFQ9kTwUEz7sSt4Wp4WKbmvNapyx18vtbDO5FzxvnJKNNUjlAbagi50hLr
I+re2Xp5q28PCBvgIPBLwqswvf7YxBInHeXzPCljmG3yLqlvagioN92/qWk96FIi
ogCCCYjDHc9ktWoG6OxEvQn11SYYbxf5BmiqURUVWP3UlOCm9BYrfqNsfjih8mD5
Nm8nn044tmztPp9kCst/SxJsjkVoP4XzaJ3y0fyvWUrToK9JGSMZt0bsjYj7qw/J
QbWWuUOBzed68lsgzeAb74tt5rIMMbxc3zqlNdv1zKxrGhDxCvKvEuYyL7793kpw
EM9/QXQ1u+/VA3oCu0HtVMvSksrFFReVb/rrQHxEB+sQTmYu5OgxCtjObb6CKzMw
W8A5q99PqavMun+JuZs/ukKhk2pHu92z2rXZYSMJC2bI9NbFjct3+27FELX3KmYf
1qmlmJAiviowcQdKzzSJV+SaInDb7G9s3+GH+uIW/CzFAMMMzmpk0s309WYLwC34
s6Ogm7KLTCFdLJSCNX486hsy4fMoUl8WSDrVSyJFL7bDT13M4bChUqd6yFRBM2lo
0KBXgaNQiuvE+uq5iKnjFAT1AEyx7hLs5jHWnXAcRt69E3EqXtCCK/peMhAKWmaj
wOSrCL+tGdFvbDvzI4n44JG9i+QhJ6bbbxW2WixMusw8Z9F7voKQlVaZCzjqTQWM
3+BDiCBexdgUzcrq+s85F1Y6tuWs15+tAE/tR3r9/AyGvuVlb+CCewsX7d/25mLq
lnog3zSt8pQUbdAdU8MVhAoB1IZ3ufNGEzSgb4okUvZu2zp3mVXGirbo1wEvT8NI
WSE8vamLxkd8AJFRYWX/oLo0E4fG5F6adaFoLnEvfCGg4P+mbzbPvdW+VNsSRbK8
8mLM0B+E5hyBLeZRBTkwHX/aW2Bj4CrL94An2pUNeiQ/6BuEUlByNGhsBaL7wrFq
vsQkwrbwZerrgmL57dd4bli8cNIW8HXLcQ38y6dOQW4f8Q3hHweuDrklJI8k4PYD
X+MnmsBvHotpjBAao2K03M+NcrpLGJheKVzcwxw1h5PkiUS+Z2n36VnRN1hTaO5q
WRWMXvgw3pCdEaErVwRzwV8dXyir7WPVpKj6+crRMwA3VZzZ9ooXh8K0FFu/5BAj
a4u+1lKmewf6MWlKxbspD2aVfaSEDxZ/49WgV3lzrEMUG/GruWhSHm5fqJXXDlZA
PiuyUEmckJBgjEWWSExejr3wrbvYubw2qAheaaVYlQCmyY++3Nzndod8995r4pLd
DdyUyXNBXt49SmWGGGQSWqCgvyOn2jDjpwp0TDwZoHbPQr5yQrCnCNovjpV5azWv
5hr7IZP3chi2fioRV9+/VHz+uD/BCKKPT2Oi2I+/0IhqRzRgdZenkkN21QTg98J6
`protect END_PROTECTED

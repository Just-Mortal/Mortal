`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+uUx2bvBhX97CWMa1wUFZMC8V1wYN+VtiM28Z2zF/GQl/4ITVRTNpgOrN7BvbwO
0aju09NDDcRQqGCKPHGWu7qhF4/5pVNKrKsXWRKgqiRFs8FJ7VsZDq09XpVGRZGV
VEaDJzpJwAXMqx1jpBd0l6w/J0MUP+FyEW1LqXYk939AxRatns6zGbDmlSrs3f4A
aYSZNUaIaow41fbIB8kL8iWcpaOLr4O78KtreJywZEFEFf8Eg6LjmmmrXYGQiJmt
UV3ytDRMBvebDh6Q1CG878GSxFcn4kKkVUydT+oSvfhaq7TtPlds3kfh17l/MDSt
C+2u1V3va6vvAyuhw7xFast4FpJysZX5gGLMsmBfpmf+C8IXEZI5A5mNw+LjuXkc
h8tQJ8YExnMbO63RRi4xkfGn3xsBLUM8qW2p+A01yT04gfz9zBD9lyBYnPGQcLap
0GDGFVCLP3Vv0uQYw5ddxAV8A3cqS2W0ifdK0IcSOH4T6G6WYXpD9TMz/jITsuWQ
lQLZBeomNhXq42aFQTRurCCAptH+w3K7rp+Wl3ZRkiz8lynefFkCITuT+QvxiBUC
N6iQ0s+Z1Pn4z3gqi/SpIjCs8AOapbACJ7DqeDknyenxyLNtA/DxGUyBOEinGi0w
1fuNUmnqI8cdPFjDdsp6A9/rYtKNwPsZwtI57NWGAZ6gVuFaEnpU+Xrb3Q2xEAPG
yK6uaHGIofQ8mWM+U1wW4swkZnSnB6LTufj3Q8FFkKPYgq0d8DWUYH7hCSNLIMtZ
137m8QPzj68BgTF9XsS60WSrp8p0OlfwXXbBSFu8yDix40bOTGZnDSTIXZPjGZdw
yGA7Ffx0GJimCzKZLQlqwqJQPVE5k6xaVieCzo2csXQm6DqcHOFAmKEZKcahfvcG
pie7mIrdZlUvSKtEnlHKK1tWqUspIqZdF/Te8xJPyUXCohFw4dOMwlrjbVxi1Wy1
sc56q/QS2ZHi3MU8P2bv0HpI+61alCCmRSIL4bBj/zM5lCM7nsype6XY6PMjBPqM
A354unQlVrNTB6gUnpm6x6xX+zD4S/esXAi+O9dPx0HbJl8EkpW8OyhjDGmv9bGV
/7rc7Y5bs/kIyVP2vAReDTEqDSoQvP+YTGBZVRwyRd8Fb8/brmYGxmcI4cRF83G2
K+624dHSegmPALgeHyMPG25f+rekr80vZswj/Oldl1l4A1ApA+796gCR5GnUo+/b
x7nMN7xIMQnhhqVUS3QsfHB0a6nIErQeWGS9jWi7k+APhRfEhQ9XEyNDPA5PR0UY
AJ8pbZZeNQ+dNXAf7NQHZF0vWzDW28EenZq4lwhXCy3y9dCpamK4hoVAcYmYsw71
JVpkhP+J7fKjNJTr4AtZ/zZ1qRdc9rYH93DNJ4AVCn3WS9ETiLA44f+f2oLid1GU
K+JgpG3ii93JMNOG1/pwFjDtZlGUrTWoPT/RIHUqWsLSNq2VoICGeQqxCXTPwliY
mKh9h2UKBuNE3G06anVxaEO9Z+R4lpB5IhwWS3r0EgtyGlCThWxZO4OGCnzeFoQ9
+tdVtsDr6kPEgyyZcBA/xUG1Nqeh9tnrGfjyQJ3F24LkDCA8Kcfst6RT7RkBzHly
KEoYxL49skZgUxamW9PBG3WWXuudpAvTfo4YLK/j8mM4DNkD1qbTkZHekUn2Kp5Z
FTKYr7K33aoju2D8MrbwvzlVKbqALxDMt5D5nJdH7VqsWdUxffoCYCxXU0lmyfpM
LCO79cScC1BjfjvoDt8XauuyouQ2Adj0Dxvf2Kg1GlmWvvR7gU9FLrDL94+9hQ9D
Xp4GRS00HTfrpxuVbC2L6WpGqRsXHKDt55UbqHI6w5pQUURcTkrfEJLZIdY/Izyc
pRcgYnoUBG967pM+QZFCk8SDRwpQgSJJwovKODqvONFe+N8yjVwVwTz4xDdNtwkD
VIsH6aENP9plhooz20JabfiHPgyEhCWgTwBi4H/dVgUGMrT3FaH/fncUfj0MxLdS
d3L0Uwnb0RtciOwuXBD8nFgfr0ClU7IgQBfs5K8paw/BUQHyWFgWn8gzO7hYuQFa
vQJIpAxUmbSOAl0YwATc7VGziOESIphj6yiqOy616vX/HzvZWJVpHuZ6rPbBJaO2
uimFxi56sO+tevnlwzd+bzuVJMecEP77kIbrfefKPZiWjOU309EqKVKWizPb+Xze
UefJwP3JFFMeY7JeVWWYtohrX+CILZDgFse4aEvGM8HavGz+cs82m8g7Eueg8XbS
Qo22//H+wMENNIKfpsuXzDiFQViFL+k+Sxk1UeqO5+HhqzEyyUpbTSmRFRg9z0rE
8gycGoFEGgbvTEzwBiLMrSyojO6kVnsMW/E/Anx2a8JDUlpS3lVVCWff2F89QnfP
SdMcUcsAWO4mpov8fcBtdt0sN6Ls/ydBEeDbqq562CusaIjB4S3heIosGY7w5Kme
APDvHrcXbScrszJM3VKAsZszYyPe6v2O90FBzZf+jtKXf1omLLM+UQfFc89ocRiK
8GX5/uNhaxLo07fsdYXFeYJj3Gpb1m8i8gEwY1pzJFH6z/W7yKuNUtnfi1/3Z4C7
RG6rU5e+VApse/rJBlK46wHq+QMo8JPeNLNofSXgPk0rDFX6PMbl8Nxms40vrrV4
ngZsmNrjdcsKRO502o8v9ruEu/BA8i9DBHH7It+/mGewQ0yYQgtCPqnlFjc15rJ8
Wb5hStyFL2HCkU7TX8yqyIQNFxtz+mzamAV9s3GM72qj1TC/+65Jw7n3xt17lJ/f
907zXa6t+XKTalnMdWsoPaMj+7GhAKQ8oEog04dq4167Iz70e8CBZaaK5cvoGzhO
pKkbxgC9k5NXaC9HJWWUDdn7nFGaHgzuwm8vB3TC8RI3DhGBKidRgLuSso5ql832
TZgD14El8tgKrrLQhCMkTkRyadwrfUwcrd7TugAq1ynxCSa5DoevpG8Xt8/Rm9+B
V9o44+ZhHaqCZVrXhSJFFivr+QMTg3LDSU636aMqGIR7sxDsWfh8sGm11M7d0IKW
wcszA0q5/bp78IGKL6ExRe5Q91kdgK/wW+mKCAJaz8oewQkUR6C6hBepPRQiG1IK
8/cDxoAUxP5ZrjvJj+iKhPHvO/ichBOxbXrlnlMms7w4iFCNlb+4rjFGcDCpxDlW
aPkPng85Wf3QyW1XItdrHkAqvNSiSEGpPNLe4C/DZzFAvOSxVQioPFwgkNXob7bM
j56TLT8N8gq/F2QM3owGUOaIwBJcJAOSOiTXlcMgNUB5BD0lqPlktsPgg6mIcGDS
IJVXE3uulvGXkglQTUIUZl00hI0GiCYcz8HsMzuDiLGh9/GSxXBeNMFzs9Yu0DM5
jbVyewHckER/gQwu0zZ7xuQCQYxgTGa2eO56Qe6WNr6ugpeZj+jCf2LZ2VN9Uh5h
/5Sq05TvlBwcSEHGTMeZSGgVR8S5hFf8bZnwwKM7CCdb6814EFm5trA2zl7A0Uqm
tIpJ7VIUxXzPTfEGJ1jYQvyKOC0bBp4GYpAc85t/UwDQVSPhRnTPPnDHQfgYB8Hl
AWt+0MYQgsCqn/COxiM8c+mXrdQapkqFhGkhLUI3UYf0xTScicyZCPHeLEqpPH7v
NWbfi53so+8PhaLP1tHodixTH/aQHLd6NtpeXQn161zYLtZJF07kLUalxuBjS17h
ovrQKVi4YQl9jsuM2K5efgxA3zUrKA5FYfxAfi6jyMb6TxgKkUHt910bxVoHmosR
IaTvEWd/Civg7vBSJAdfzHmKPjlN5anGwiwXYZ4YGx+G3/LLJitVKSfCNrCea/m7
GSXYBZgxSNTZ81+dmlVt1OhQqgv5Z7L7i9WPPZHOeF608b3zfQIa3XQFowOyWlW2
9O8B0bBYZ/foelwNCHbXPXGfou52px5Cd6Jb/Fi45DoW0CYwx7/gel2Ehp5UHdUO
84fAPNhMvvbTYHcEPApNZuFu9Vv5dz6PF/V9ei0ahgTNBI07V+prVdxEfKvioMfv
/r783K5n/i48GXHRVfH8VS2jJgo4+fdERwydeNheLF2QXrOWCUuXGV8pDJAiTaLp
YZncNWR/36oYQYaSiy0oU/hT2Afx2rIS+7yTfQkv6mM8YpqavArevhA/4rQpJ11X
+BxUWXpzTRuSZjEQg4kjXltIHxmSyJECRLK/bb+jTDKGCGOoNiNIEoTjHJJleGcm
`protect END_PROTECTED

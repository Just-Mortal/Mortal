`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdRD5vP/0Gk6aYsMxn1uPkxxSVUOC9i38nnkJoYPosXxe8KZSd0VduGpCgJxiL9b
capwROCjR9FelkrbSud9V3LFxEosJOzS5R5fpiRVobdysw4mawDkdSsamzCT6Mz5
/DkC/IQqh4jSSP9POsh0p/RPAg304JBSQiKMLYnpdrbpODWwmA3GmC12VbSSTwi/
cbKqpX8tQnruKjjSzlqmxvWvowSMy2Dy0MeB3AxLnjTXkD0J7e+WBuGrqdRDIlsv
aX5BwZzme+8UC7x+wO4Z/Ztf9lpLbaAI9vGX7bUnwh4/ssSaMzD6uXSTEraG2ynm
f6taKHFjZxlqX+A4gVjQm3UbyjU0Vb6u4yc8+dkLmxBIh7wg3nvcH6ueYsxTcwPx
KaERTDMqQqrmu7l6j5lA3IxLQQHbzqy+tgcBotf3WbIqj1KO2WUjZrzEVtIKzuXK
PPpl5UFXzXVUb6YKm49qsjFmbd8uz1U2C4Pql2I17mHIEHACiTS1ryutnf9bqP9q
CuXFVYTxz/SQAggQv460fbIPU8j9X2/ixwNuJp+5X0paT1CKCAj0eQj6Xc6wHjFa
rfnyDfhkweNG/Bhv/jsF7YXX07utLzs1UiXtLhKNVLj+n8/yqSHDdGtXcR9KktDP
j8BESPTaIdqkcigR3Chp/mHvsk3XHNDdwGt5fbDtRXNf8vJFqaISI4jsCzUqO1md
DIAwcnVUtEBjnUE1fNOmYn7tcHx9JL2pJYQJ1W6LypBLfDBmkfjm4rkqvZZbsvYP
7xesCNbf6FDldKwlIlU+c1/R6mit5xHITCyXZyyTHUMe7cGqtrSOpW4aNhn6sODp
SPNf1dj60CLXcmlyfQjbEr6l870b8uPF+0SZ50FnH+iexjPqBmDErNFAGvtS8x7p
MYENSMd09QmI489J41QrxD2tcI+Vs/vYrXKRAvC0ML62TtfJADQFibc33xv6JD1H
CqIfjMxpyUBCWQSC1/j6cmF5degswQW2BOKhW5oGzf46L5kNII9C2ZiGavO3oySj
zzE6HaMbWExPtCi6Te3Pc03vPmxBoV4YU535jTMH6RI=
`protect END_PROTECTED

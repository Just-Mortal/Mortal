`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GU6Passs0YFnYYlPjZpv79/NgSC6Eog2xpYOkmGuEQHqMgp1nAmuMS2tqSJ1OYAD
zKVLhxMaDTxAhKbVkE5mhorC2WYr1vBqZTpBChZGr2tRWZTHDCNRd1U7azVWlwLs
uu7Dh57PXCgEajWVG7dLYrkijUvmppjXgYRtwLQ5vWMuuZ+4MIsnKRPcm/qsfBAz
gqN9lPF9f0TG2rrkm9vGCTMCYV0pNwae4LNh1A7YIL8nOikr4FV62kQCtiFtyBvU
l6k66Bwp19saDmAgsgqI7HWd4RwvI6h30JNTBTtGYe1CADTkM0Br1foRrc21wQzZ
8Y7Kzz5LDuumRO0wyj3SAqdZru05otlnGEacnC0fJGwVusm2+xOaTBuOQU3ruYDy
+2KirEbtVH3wtLYAjwUuf7zn/jSSGEg9C+zVEbc+wcuvtWHMfv10loiCOG6zrfXu
AQZJ1e8ih+HPm36t3XjNSDcRpl0TcixR+7siXjHZ/BRqJo+7dV9V0RZDl4euhT+Y
GLbguf7wcrOM117Jge2DtjaOhuZGaV5Kx4oEpKGE9/EOl+4FojK/SZ6qvq2E7wMX
WXYpxgvBD1P1SCLhcV3/rnVqTKCFhi7ly004gC3bTMfWCd9kJi/risgWq4jt9Ajr
CIhaZvNdoZpGsWGmfqXYeQWrfsDmY3HNoi5UK8h0iIUxfjhvI6nfeNBOxo75CrBe
NfMe21SsWb8R9B4gzBOPWl0QgtM4wNzE9cF7JF6sTym+m7qdqr2V4xHDQ65/5e+C
ByQWIrVaF7ggmxx4PoUOzneKDwOXw1Wb6ZW91sX4q9Z8oTwnuh9oP7eaMg0qqLdi
6eljATbdrHAqPeIFyteigjyq1VipWD54Oh6Vrw1n7+ewTm4+6fQzrDxp24aOEJIO
AgR7ZJHOzgmuDXntRVSqc/1Kj+vviU4Aldzt+M1Dr3TQUobjt9ZjqEJpCalP4WcE
wbEyH9NcfpwNn2kjqXP+Fc6HngALKQcAYo03oDhcm61W3sIwpHrl5mXC/TW+5SJ/
hQxDP/Vi89bhQBQSiedhym3KO7tg1EjUa0KDMcgUMhOKhT8ETxvd36I2kBUa6bKZ
kMWylGXdGMAaCdQiwHGYyhnQZgFsE4YEoy+XY8FJpM7AN71FFApbVlPMpVf23Gmj
0SIahqDYcc8BGzLB33hP31CV0xF7a6hzE4U/Wujw6/MYazh5S3yeKpCj3h+ntugM
8B9YV+ETc0NCZFcVNzF82ibbbTMeYfHBngARX/L93+3lcVNRb/YUX1eQOi9Npjns
LhyId0BVNEERt07eOcDxlCh/dD70iDnu2cNH+UchrRt1yLGJUFeBa+UpnT2PGGdh
LzK31I2kI19ciow1S9wKcQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cy+HJZNkURh/I8p2Md5VvfDDXwWS3LW43EdPZv9il8djeM3FwbZAZ/hk2erGyFdC
aWnzJzoPM0Nwe/QIGGHLJVOmsURFWi+wkJG5y1wjm2vM7kX5GIXLLuDYxYXCDpfR
/JhOSqEikszW/LH6aU6AtRFD+zOXxGlBYdd4Ng//WH5YvXB4h2NCPe2Ahfrjv1qL
Jti1aFg9sS7e7PUWKhPO5gXVgIk8Ricg246IMWPXtu4nqZarmAdBa7R/Fwv+E/Z+
n5MtnnJpY41H9yeya6rleHxbs/fS94DV6eKPm8bcyAow6V6szwj8OHXnlfBPwx6Y
lzvgFsY6j5ddfYyebj6a3duG59mvS+6VtXAHk9EEIOKCcC7ziMq0tYbjI2550H+4
N3S1w5WZTB148nsEQC3aYZtBYgp5zEeCCsK6+uapu2JpgNw/gSNtuuH6dINH/dZX
5ETZo4ECqQnWBrEOhSDyuOu4et35hwjdomVh8k+AyLW2dX1Q6DM1MgHkCwWLKqxC
X9wLVON6Q87yhzSr0hSkb4NtUk6x/z+LGOexhOKuRFISeyTHeILvmzFa9ylSlFBj
3w+iBeJROYOxaVEqqgWtNPX7DpkkxfLDrQnaV3sWu82gzRoodg33K0y1O8aoLt01
ejsPLNaoLRGNdaW15PgVluQVaqwZWGAy6KQaoRlp/fpBt72O79TbOnQ9DOKY65lh
a1sG0TKmdfuIjBodW1Ml6flvSyIz4S4KCLREWguqjpdv0QWjXIYoDdE7IqVidahl
n524GnvtrtV2CuLxekZ5W0PCtZ9vVrs7vv1KYqcNJT+1haNIkVKAMQ/oRXgRufS3
M3czkMrMG+lMg38HBz1RciDiIJr7jmJpTCcDk4LbJgrXSJLtjjseLeDnupx3af5W
3OJg+t324sWjLUYlsWcp4wHtZExoSkTFPnuElGufac0GOBynqvxk3hqH62MXD6zm
18CimmrlYd4e+soof9KKj+bt48COBMhf8fOaAfhymcaz4PmUJde2cU3wEEqNWZbB
VM7wtlQ8L2hnLnrtoe53U42SznFdAkCTt9Pl0jAHCoHBHySDEkc9b5/1tBbGa0uH
F8y2Ob1ER4M/EFawzr5j3Z8yOdGk/wJWsUSDNJEY/1mXW813CToiAc2HRU1AwuIk
QPW74Jb6RPy9oN7LlXO9Qy9mX9McyHMOWIHh0BSgNvi1ozfpqHnH1i1RDgSg8NsJ
F9Efg9NHUuYk8/Ml3wIa6TfhoeMzTjglDqTvzaoI7UC3qc2wA5jQ9Dt+y6VEub9h
+aRVzdO7ropZSL4QhSJh6kG8XO45Dbj135vTGyryqqTm3VVqBqrcJ90wVQpaKY8X
aup3OFwWUGHsWfIahXb8hhHd4ohFqVfO5bLsMNmqI6j6rKrBWOJe8qTrdC0XeGvA
81e5+4BFcVvXnnQabQs3JEm66R7pdfsLZo+ZU5digydZ8UGUH6ck1p+V0qMxHQUA
TPjSuyTCwunaKhaXABrCnjS5hcyozdiBJ8e3CN/Doos=
`protect END_PROTECTED

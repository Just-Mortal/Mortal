`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7LQMfRRxtE3PV27SlkLQMiEWa41hYZh1F72fcDa4lCYiMlSr6MPVRZfVxh8YSw3
JxJlLoj6d5Lz8OZr2jouGuZqyUM9hn2ekW5B9T1xsZ7H8j6SfmXtF9vpZubMJbLI
pIRlOgAtluULA4ReOWmwbnNjrf37xlSubPmIryUez44xHBF3BUgjJmyFp0JEQoU5
+4uU3CE5ZUy4Xe6FcRjRgfqs9Ts3qQRkgmvG3FylyK1SYSrVyEODsktvzrdgSf8F
e4jkz+NtoC8B1PfmGtTm2sJX9szo6apjkdpVnPFFYo8qc5UHEOmTcvarENfti0GM
AKl6E/hxek++dt5hSGOQYDcuxAzQ7YephQ0KWZtjgIoJLawy19PrG3i3SJk1iqeR
xivnRJC3CUlENajvrKUkApLlKkYE6tSAeD1y8KXhoP6uplUFNxOwZNxP4MuTS3MD
VnrgoTZBmZI9VoRSql8LWbhC/MJfErPdGU6d88woM9I=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djvInFnbNM2OH043TiohXP23/nuHhgfQILvwJ7gC1e0dfVAPJVbJHJex1/U7742x
TsX+N1P3UsTqwlLms38oAnMRPHiSAOlo16bp7mYgZG3pY7Zz5DN20NCAlo0pQqw6
d30LXAAzJFBAK3PxmX5wMcOEJN1TPqyRaWlSPosHGXrVOtVUh7QrGIjfosyBnTGJ
1rQgB3nwsa5nGaMz1hZXWarJVRMAaYwB2H7juLpOw0BufGIb4O+dm7J6pqN5ff5B
xmEXEKouPZDISwmTSHLTS5h4ylZEQvUv50U01hBKUE6xm81M1cLseMVOcp0QD7te
zYTCN+nPgr53jvFuosacoEaGbQE4/lRyh/eCs4f3EYt8vV1llm0RiMQeFgxi0wG0
8sI+gvvuBEULhJpCXBL0+I/L6prhb6yZX6ea+XYxv5CTyh/+Z/4A4JP+hwpP9scr
EKrfeiaxLy/ADpS/z15xCP2ZlstEuMiam+wAnO9jNZEAkVmCiCHoSHVgYyP5RUcJ
10KluHAdR5xVjk4ERGU+O3/CpYrKqN292Wg5M4y8bh9yS0D1ZpOlL8199jcPeU1X
o7EqAsOX0B72EBla1xQEcVU3tq5eiU4Ao4Iy2yJcstbhagU+1SyYNE+OALk3jcbi
lS7N2T75xZhX3kYQChpKQBo7ZljRpjMe+ET1oeBFYaKzAL9RXsQdFLj/mGSrkdEQ
KKQkrtsIirBhEhr4Z1tVop8YWVF1QgGlBdcbk9zHpk+MIieGyWG2KU/wZcX90Q9e
ulw0k8BHC0GEhsJEkAIIgzCB58PNBGoBR6Q1RDtrh0HljSbLPKmXSYjxGGQ/4vwf
LMHxoqKGhdVJBpt1fmSYWPI+iCdu7hrAJp95jliccf8BNxaTTyNmF9qsYkeXFZY8
X8/VoCsYCYwsKCgERphpQU8j77xjJjq473uVFuH2jd2cU2nitJmZCnvrQe1izCZ7
3p3Qs4gHiuUZSQCbUnsmk/bu08Pw3eIh+qK7K7ECKYpuQw3u23fjO4eE07GRxPLA
cOVARLJmqYpM4wUWWZhEFTuJD49MzB/u6Xi9/rhEIr3N977Op3Dbbn7WZUKPWq7R
DFWIEtJ0f4zuNKStmBLy4pdLm6uu3/gLhiCZirYD3kt8tHln4YLn/DJy5jlQ2NU+
54oidbW9VcyjhJVuljtMfIOP2Vs8ut8gmOLZKgzRHhXn/on0s6qZWSq2Xdy+hHmR
A1JPa6dxDbFhBnW0X1Shu9dORPcvn8hUYrDpqj18ZZ2xonE8s57AxipuJWgpDt6o
TKyAcSxRnQwxPf9XLj8BI4Se6iQI/VYe3wULm7a+8/lN/IYyae4XQ7/4vq++Z6Cy
u0IFVF1fHg0gdYN67hRU+RywDHdr3jE6G2LzOJisbGZrt4cbcl24T1joi6QBbqt5
ZVS5r5Y1nE7S12EfOogQINjMr7JkXRecUsAMaXdBxCTN7wKB//i8TKF0MkthdvwG
FBRhb2tkhf+OedH+W1FyHjY86Pq96Ji7+0+usV1um6pUpZiW8WJLir6uMtnRzSBc
ABnBaxnxDuTQyH6gsRteh0KNS4YM8wQrSRZkKeM0WLuOyKvuz28NmjB7j+n7CK1p
4wMa7l9jaEWVBeStZ8Grz4OXfLsa3hHBla3WbXjoO3CcHG3L/ioHLWAjnSR3agTn
qu/jwI5H++DA2oCWAbazS+IKbFDf3trU01nJYb+yca7iasXdIz4TeKtC2VIDUQA9
RG5suArzYYz+2BPD1X04zGiEpekcyOGSJ8eTlgCaV0wJpUU2F8CL4xjgMcj1fv7c
mpDvkPFxZyV8hn3DzUiq1K1DlYwl1igPqJlmz1aHvZDjQ0LeTs30IUIlFIncSGxF
/FYyNkZhyOPRdNMS9/EcUyk6SYsQ2Q6huqtNw3sVJQakqPFtToyxq7qMDJjJ/BLd
8nrjeJJgc550TFQP/u5jXokwXLRUbjwaLknOlueKpeGTmNYQ/cWUx2hHoR47UijM
k4KpHpGumwPinQ2P1ej2Qy5hLmgbYt+UIPot/g2ykESu+6KNvqEpYZfmvd+TUmNx
wCapqHUUmxIcfQ+Yrq/lF2IUGx6KSbI/uLqhddKaKVAFbjD2FJXYo8gbuTExCz1F
siDA9dCdbkSD9ZkpscCM+X7SjbI0ODtGpQV39QBieiXyE5+Stn2y70bzIZwNry4X
7XX3PUH6JNd9rPKjcOfSNMZXcOR05E19McMJVFrs1ieNNXJFmgXtHisVeIgamgiP
Okbqj95zJQ94edAakWzPqJqQJ8LCC5XC8wIVZ7kScfexNy364w7aAWsQ5hzENEYF
otsj00JXbxetqtjGIv9z6fLSuFf9f31t7sAZAAqp2i6x8l4ZvODEYaopb6fcT6/A
4rZ0Z5aCcS52Y+6EjpVq3tl3jN9z8T2pf6iHIKSJ1gQXdNEhm6ff/ZKbi7bDsQq/
l3hznMnE8oiErkywOCOVDvKDWPbwGrVfj2PnbLOCoFF4gOjdcf6FjsW2vRSFXy7j
Rlvuog58Rj17QElZJPJcIQ==
`protect END_PROTECTED

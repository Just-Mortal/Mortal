`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vcfj51bPitxQTJqtwFPtLZjQOGjm76oLC/K/W0t8UfZhExEHyIxzU3MrJZxAA0uQ
BW/gx/vf3ja0WgZ7HS69BRo5L1p6DF39ATFu84PoqiomwBgICd2SD7eXSzMXbXIE
qHI0fDtBkniOxzBxQXTkKB3xmiHoMMSUbkMoC8ltJR5TidE9HHPH2qBWRtFPUTJ7
aGJV9tjw0m39gHjDFbaeTv4lkVZiQd3AdjhhDs7p3c3f2TIJ5cf7ng01ykPkrDm7
Hp+fOavDKEovVKwqMwzNRVB8fSh3jLHcy6xT4iCoQTiY3xk9uV3yBzVNXG9XYgVX
avJeS0wXHDku8L946WCH34tf1cUrofaKrmCtNbcyXi8AEouIJ5D+I6W6OF/0jTQl
TO7l3Q3uh8Ps3HYvAjSM+fqRYR+p2LPOnGEQpeM9swe9HAYswAyL2qv8i4fZRhyZ
qN8mR72lRiYrTgaLEYEA4PO8tYb1EjyjDaJm68Uy5KjATLFQBjkUfbai8iH+HVgT
4dCtLO0wbNF2LHAt5FlgePk/pKwn+femB/0qVriTPDyyLEqmpBTAu9yHBiB6GS1h
u/yHarnXKTxckZP14k2fM01iSk/AO/f52vNKf13Bf97tGqo5TwA01sBrq7XbJt+a
K03GKz4wHDetkZeiVrvvDSI+Buc08pf8sGgkwo/iSRVCv7j4RHIXkAp8AvYSyKtc
IMaIpMurZ27WZPPJddRUMI/TKwXkeu0PePDrot81AjfKwyva7HXmyCsh7aE3F+ij
+jkTPpPtM1vWMGdntIuASjQdW+4Lf2CqBe/uUkRLKW2NIV+RhKmLOPieiOCNYgz5
PYlYi+RbzByewFtbcRrp4WXVhobPXeehLdukNgHi9ICebzxZnDv1vwqx5cBn/8NV
fW+LrWA2LVQXLMR1elQRNrQ02uyPHCErNpD9hisV5No9jj7SgbyLCZxiBB/FbJAg
i2APYWgqHhXBHQZ7Zkv1vb4Ht9tZ2XUG3Vrt0CN+xw4yubASYasLFFlbS0FdSd5n
dSK8u5l7G/0RPFULali5TlKZNt+3bxcyfrY1A90VmR9ingO3pLmu7WD3rD8MiiPs
iedqIHANwQINs+qF6KU3C6ppltLYDnZxIf1hm9PFwxp4fLO5SmTgbV+oqz5jWYNS
ghtOcbRGsm0Eq00v/VL8YnwBNPW/B+LLSrsaozlGyAxkfnCmg/AGW+K6R4jn77i8
B6ApODRZTKpVSnHUYW5mHy+AVkNKFWd6ERLupIPkKhdk1lspU7k1KxtnttHIC2ka
n4qdajDa6UzsfwdMFz0DiA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B7lTzRXVHqOk0lTxbQ/8Bn/mL6gA44WVaLJef3xhgz0YNdF15PQheFU3V0fRwN6l
nIDS0F8RTAub1ZnGa1bXaq2DZD0vSa17sRuQCkBUK/+alX+xbHXHIjb2tmJ6uKbs
yh7irUcJxUkWJwc9ttY7ilGOCT12jxpBS2SnsakyDuJ0xZQahr/peT4HRE3uAjrD
F74FBWl4FhSbXbvOR7A/CrRhbB5hGh3ZjQmWmDd176h5U1bi57hrsxwRajVg3r/I
kx8tZ/skc1axxZe0eAMhrfta+6gXgc44Qcvzs7aO9ua6wVhsZL/IxY3pNb9OZjEu
ip0veOXYCuw1sa5l/PakM14DB+88krdQ0b8VwoTuOUa9zq3y6lNIR8cTHWTJqIvP
FNyVm4C1aRH2XINLLjTngKSGPbmd7egmZhEtFURPCkHKvl4FvbjDcjs5P/PiS8qE
dtqn50nYMwSNcspzw63BBh5ku+DiCqAFIHX7Sj9tHWL68ohTtxnf8usdrV9xy59B
Ti7xY+DvbrYfK3ZqQi8KZBxcnhmuSd4RxF9LQykL9KIGyZD5osfqfIsNSaTap3kl
IrYU0zRQ3A3nDchQ2lO/xwJU0VT8zW9I4+gmAgGLO9JcfPiJt+rN6Hx/Q2Id9IAM
/s8EB7Qr5qoeJ9cXeR+5AYYTRorHqOOIiA2oq9vJqJ+LO/d2BeN2ViymL8XVbG8d
Xb1365iDdR0rrFGfMzAvgWqlX1QreRLeyU1GPX0M+YnVeFF0xP8iSSUxMp2opt5H
KNElczP0FYvpuuXg7i9MMNC5DaJty+CMhFX/udrzDhl9tvQtYQqGxcGeKIhEsC1E
Qakqe+/TnNkI6HQYgPZzx8vYbjqoZAL6n6/2a43Td9GPZtSlqBGGcC2oRgm1vks7
kerhvwV1s8ubyvFbHU+Ot/vsZ2ivgXzHaZbjiFktkCGuBfLW/mjI5sMIIvALpnSk
DUfueolxo0/idhJDjO6wykM0MRCKGVd3SgpTGMz6fNfEj9rrTy9zY4JdbGx1Z8TJ
CQd3F/5XlB9QYXcVZ5EkjrhvpIyuzNdOVbd3tgXSzNfTxeWc1CmSmafmNdmjO8oO
JTTg7P0bgxN6iBBgr6vIDyN9YNTUSFQUHFIHiGeeVaPhBbOXKEJGfu1NmpIoJ7TF
EN2qMFshcsDeei3mp5D5yu1qgdSrpD95jGN0wQuGLQT3KKcqmyytDw7zLOQ4+19+
E7Y8nARdu46KZKQDNwZWZ29NInTEecw7zpTCkMkk4ftUBF2ZnUUsTFtjhHSDl/wM
TrSb0RQJQrpeEdR1d6kh8Xe5k8cYYwLN2pxZydxL4bl6Ls4JkVjAxZ+/wkXI7yK4
BOqGa881h5YT0BDJ1bCbnUyGyUZPmm1SiUO5gor1JGUY6O4Y3W6Zuh9BjWnDP8H0
Be77LQ/VAm9K4zAtpZW5amq9ZXsL+Khknvf9pAu5bT2N2iqu2+ebegppe7KM+nzV
/wDTAWKw1cxsVZcgivmx74ek6bxNbtk5+CderGH4p2DxWXb4j7iRJMq2+HvG7Gd5
+461ednI2FJtcZbnMjYOiv580U6mGyM5Wld6g+CUZ/9WzTYHsd6vKyc1HhxP4F8c
IOTuq1lxD+UdBUA0nl+uHowPif+7EdaoDb0MdeCUDNvUC79bC50domM7Z60T9vpR
BQMK/NCr07wZ0+Qg2DnavFCY3J7OmeXPQGnC6zVKLxlF5yg7E/WniTTq1tjum/41
O8o2nziSsI3g7DJbJU8ljofsleuDas8z3dXLFwPAJ+bT9WFlNrnKwOa98un3cFFl
IcvskKBtu13xS8/hdudvWsN6Jd8QzGL9gb1AOVB7rsT5wHTjCq0IPlQ7lLJ3HFpD
p8jYcQRTyxVpMxmfhAKKm5Neb/Q28X+y+vGgDtJR4BPvjN4tdrxsCmHiQoMlgyZl
hbUgfTFn29RFj9wkEfyqInFq9mfC2iVfqYqPhA3gV77Q2ZxSJQ5QMV4mmuiRSa7k
z4GCItTMrZqK6/d/42faYhHaqnO9DVocpzqur9b+eMz7IsYl0Lu6M/cCnlavLwog
0dy6xQBYCGe1v5iz881LKU22eOVy9KjpotjXZK/PtgnIMqs14r4LcMDdBO1CrSpR
mSFNoCvu+thfX4c5f9osJp6U6hmOLanWcHqIWLvQMF09Dtr2Sn7l8PlrnNfukyxE
/TF2iZs4dvOTuxce+gnkSDCKGV4ZllsPxomS05Q/Ib1t8PKpGZOxCNu6Tn8+zMye
qHc+shf+wZmjQ9PyhKfn/1r37poqK8VKN7E9wNQtfmNJ+gDfFulJ9/8HHJJAVAYQ
JuOSV24AONkCcYumXdl7FoQlpPQa7DcaebetcnmYosTqk1sQw59uaE0idFVk3Ht7
MIr0AcCwIeOjGRae6qkhpiUXUNm94iEWiY8XWRy6KUo5UxT9qNNbnyZjsJ8s6Ne1
a08vcDVNJZwN45CWO9bTbcdO/mOujdmIF/KN41U+QxGPT09r8DJ46k4MCTocdCz5
wtkjXifY5nvFcn0tvHYTaDpyYoLk2+Tb/uXKxbDPvGvbFbY19Gpc5L9LVcbYsiji
52JMhVpRWAIAFdJuvc8cwygkW/nWFzCYu4osNpiJIFrFlvKiwwuxzdUPEMKLcm9H
MELbBYGi50rBAs3QYhMWH4NY5/nODllgci1J0NpDPu1rgPwfiXp3GMU6YMD8o/vD
gYRbywtOXpluttTdhm7kxNPU6/Fmhm2hreK7GVKfSsHJievM0zjkAstnY4OF3eDS
lDoA9pHE0Abce1VaakmxoU2bL5+ivu9ZPuaBfBSpBFLIjf89iXxtrR5VFL93uMTs
rK8wq2WU7p/9j4tQKcK8RBAJLx1CqNHE85uWI3uqW/vr6ve9Qg/8fBlBuRAh0wO7
zarwd6Fr2aWn0rSrnkb/s1IIr4e3YviC3YdyYLXd4zoNLHRHgFJmfcpXDVYDwaA6
Ch4jmgwUCZWCiRAhPUPf6JqTPq/8QuY2FH3OP+adz+RUROiIEQP9hFCkUIBahMP1
0s4Mo3uQKJ2i7s+lrmn28YdCosrb4p65dcRghMTNp9iN9sdWQ57MWtbdwqMBViyc
oNivD1plmgMwy7Ap7lRNsFedE2AVp8j1N5D68bPiEQX+lj0sspGbObobu9cphrpp
r+fq148pmVXmZ4tYi3p2zIdv/AvEkKqpsEYTEsb/pXlLPw46VI4RpMeox/HWt0RS
WxLQykmpm5ekeltT6+zqpJGZZrfRbZXKjE1tH9QS3QN9d5lR/vV64j+EyDobYObu
VhmiL6ztt6J2v89gHzAt88+7GaaDHjmjD2bIqA2trNN3TOUyoUFdduyP1ERH6Uzp
vXmKWysvoj2rw8viMzKdlfqdwygpe91tbIwL+am5UMsS+3msssOuFYOE9Rzb90hJ
2DJVTi3meAXDTVVXXl5DOFX71inn6q3VzOOr0ePHE4bxipI3v3k8ytmbgNzRMyMh
lZ3D887ZgIBFz7W8O4y3Yq5UVUamlGSk8qrgzwEA2X/jRV0wyX/yr9qfamOwxXvR
0IFB34fVhdPBa7mj5YFdtYHwe4XZj6/dCPI+t62IOc8XUmanP+I9qJC7J7tUeDu/
wUFkgA+iktQTS8ZHBkvGWajwLhIlFKMaEjLrTYnMOnmkatw7JzPStoZYgZqDhpNq
bGdthfqjNLAIy6Z7bp0uShOgdoVADH9/hEA4n0z9/GIAIRLn0aLqY1S95JwYAZXT
1h7GT/LhOemFRFJKW8+rnAQ/iYwtLxduGgdFQNXW0CuL9VDUe9400qkckHUu7Uy8
egmSS5FxeJoH+agg+b93GVcyEaEUNp69pZJ98RxTIXDRgnvN2Ej+S97TrayzMcEz
SWiBRekTKnZwhMMjPZMf4tc76wqrn9w6w3nFr3XkTjsTs3fjy3ZSYRexBG5H5yMD
n5djZpKW5WGTZs/JrunxU3gMKCV9OZniXhK1ijcruwkPzbKW7+wJ4q5qatCpIYRi
4xPF3Z+jo8h8O9oRzfpeJAYA1L/ZkUK9sdDbgMwX3aAuynfIRVcs1oyNZWG+7CUL
TVSQyp25GSLS3FMJ2cTMaRAug8IVnYEMCTrvwF5Moi0DnQlR1VgmTPxen6xn7BCl
5RC3v4yUUNePPV6eZBd5b1ZeyDWth+/BrlMPnBNAl3XeGHnZqvavneqonF6EWoZw
DWmk6JuTEYpjNI1od43bWmjC0Ja3m6lwT7HLZY4Rv6fzxfB0uWkDkmAVWkQ7NiHq
9VPcA51KMjwFcj1vun6enuEoQSAJ7MPVh+9vZZdQh5/K7WAcEGKx1xu10t+wr9jK
hvwEwn81lRQnPf1/2ayRBWraNcAtC96ELu0Bfw436x6jy6GR5c+o8jY5A2okdz3W
JTtOvupLw6SLSi/JN60uFcqljqnuzPXIaWT6s8yq+8fQt5MTlflxgks//jJnSa+N
tqTcYuuPPwE0RiYEo6fJOM052+RtCubpgc0Arur+VGD7HMFdDzUpsF3Pdnkz9eWB
WXe3iacHQua7Je3WWHC8NzIcBCUWArE2qMp11j9V8XCtKUKKd008ScOfLU625Fgj
bK5vNPIzY6/PXT5YWcmXJ/1pB/OhSOnPbsNn6qU+0uTabJILK/4DN1o253hypBL6
R9uiu9F9C1R0yF7nlNPI6jGsheEx6MG9EX7Klkf2+tGUvWlikv0ToTWjXCiVzXzh
gNmeXe7vcCkhpiMk0CVIUaZF5dMkxuq5RJ9YXjrBXCUGootLkKe2to2xzamORr8u
RcVJgaNF+eWazuBJCKbe3MhyVUsBLdX0GHXLr4YH1Jry58C1XQXHkdRmK89oEux+
YDWooLLyiafb5BCnRCOuNJNAJkVlShExDxBtrRR6E9FD/5tp5Q93tkzMmOl84YP8
jTFGyk2+PNK9lQ7egFwz+1gs636duGY8oSDiM0kFvE+7NbISuWwuVJxSV0tXnUHq
AfganHi4v+RqFb3hWCnteMjCyYYfZ8ppDvsywTuxqXn11QANrAp85BieiuUAvhYw
wFs/0E4BMQwfE322C/TsLEfkpoBj8YivGq8aGkSpJjIcn1RH8vSExEfmGiUzmAQl
oaq/UqXZOq9jYap39r1YSLxRd7o6PSMA++5zlT6YxybKiiw6A0dJUD6xr2Kq2Elw
cHwl1LPzggDfTmMzFpuclYPPs53U+9bKuGqtmkHSEwgd1PwwHj+WbKa8KNpJez6d
SojEq+u9IiB3yL+cuBJk3dMdTVu6n3p09MIhFF4s+g9wDT+XqFx3MTkhkAIeusIt
55oklkhwIB/ImnKtsAl/S/0rUyVRd9ae+JD/UF68lXWbAx9nvTTefTcQ74A58MRM
/l23FvlQ9080+uqw7xm+sddvJLdX+4iyH0W+SBuTI8kwnI5+u2pS9VCkzgCLOXCM
5ffSSEboRiG8zxyBB5kSBRMwHAB0+HfSrDBbh1i2prbVT3iFt+3Y3mbUXDwvsUly
2VfgwD9/RVydw/tmzAvnLd25cyT8uXowqdaDGKt7VAoBfqqOII3gmJJ0T2rMzpWe
H9tPmB+vF7x+YCZTJOSdVDmT9vsg8cFBon5XUm9my0IROQe+8RhAHS98skVdlksO
HB4/80PTEx3MWxZSiydSV0WGaWNzxfsiqwAJwJ+ve7mRK3NpGPA17BfhBIa0Q/ji
iFRcir8rV0prxs8D9WSxufW6X3MVprFOfLN8yG6X+al8qLjGwZ73lGK8qq3/y0Mr
fo0UcHyPvkkbvqXsAtrYXXcnWzLRROtB9j5iPM5VbyIcDPWiZb1jwF597HZ8P+FZ
P2GECwN2lHZvgI5pJM4rq/J92KY4dS0PSf/AR8eOAXaEhXHsyHYBybRkOGHTTQXT
h/U+DMmvyeo64y7KuK3qJfp3v8Dzyn6oWR9NfbYHRpUVccUZZsCbXyNS16XGoPxi
IA3YLBRiOmredkMomY0MMORN1NhAJfpM2m/Cdh/b6TXJQ43mKq7kg4aqlW7qvUSf
2Or0+8b4PmlOLuba04qDHlh6/XbTxo2HsA55VcfS9mI7L4778cKhKBuIq9LkGC67
awUAWh7S7sCnxWQF7dBDC2GSC2eMqEv33r3gKlOCVQsajRHYVbOLBoRl5Zl7zom4
RwbGTFUWYCAK7eVf92tdYMoMeYXmSb6P2byBDKWE0Hx8YxoYmtPvd9V9/1XQU+sM
0IYHhgADz9+PCBkIF4yREbASiIyBk7vtpBKn63sILbY//UekXSesmcHgRt+EfaWD
D8KQg7qXd77Gp/DfgfWMi1/gJUngIsJggm5pgohGNS8btZ3pS4YgS7uNRJpF4u5Y
w3LFqA5G/SXiP5KdEm+yHZc9NuXFxsuOrY6nHbbGaEri2yGKQ/zp9+Jn2Hlob4/J
7qAvVXytEWUMAOjq8iwoTi7i9iJ6iQ2VPzrWXmDd6SOQxoTzwGpgsC9H7YX/XaqT
9KRdY6UI1GFEcbCSXvp1WQ==
`protect END_PROTECTED

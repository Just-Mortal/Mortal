`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8PRss/CVZvHY71GXkXfvAHU4z76oPVVuizsvCqUQX/6iWR09A9R7YL7p/t03IoR1
FDHddI5AjG49miyZinrxTPm00OcJDQF27L5BtLn8lTri1ayrRSrkFnu3Fokuel0b
HJEfa+wwCM/5G+kXXrSD/6oGhgNJRFFOC68pePuBzhRR9GWJwsz0Ok8qLgWcZEN0
4X3iRFpjz2eeioSBotvZe7kX+xINvnTZXjpnRma7a7TcZIYtmk6LBRWxq6gTiatF
g5MkZb+l9NG6AmA8jl0gjbU3JyoG1n0yzwt3JLgg05oGl1b7KtRd32Z8lgaMR5OF
fh8ff+fjxwVgjoJgFVF8lqvcf9xzK8E0X2FA1Aen4ZpC+1IkP43sp01E/CtwFpBT
X4CLWnBInBcaY05qorgmiiXRuKTLqge5i2PRSbKDdZELKyOyRX00mtbMuyvwj+qW
1/tTLxfYfTPxfuAuH0pNRB1cjebnLzE1wNm87poe1MjKopD5xXq+K4zQdKE0QrcI
CujC8QNiAV0jNSg3GA2Dgu+IhF3N/4FhgnSPltd5XjxNp1OkqcXSjYud3T+f/SFo
nh9HeS/7dMZ6mTNuj3lZAM91OSlGjn7+IdOMeT+ufGAj+7tjHD/Dc0ECJIeMXQgX
qay5MxyVo9bxxF8A8qWbveJBLeAfs0dsH/Jr6d0bnbfTlzlONES9VjAx2Ot6+gaz
+xqyRvN7xi1qK1mWTJwb389z71FRGHXIYasWEXFyb/LD1vGyLlG5Avqd9B+oGtpR
l8dzqKRl8g031621Ci+JLlf7gNA6Jx5ozSN0eOQyCGENqCF0tFnRZZXG2wjjf3aL
OdN3YWFF2QCNSEjYGbl1PL3Po5RUrbln+6IKuk8S5rlKvfUujiFSyIPh+Hv3xNpa
NHv3sIPbBfo3sEDtf0UaXC9rxTaVf38kQqXDwBfpfw0FuZuU2JwCmgTA45PrwBor
F4sh1eE47kRuB26ZNAhrOQxuwpZ9VyyspqPKH62yNwZvMWpW2uxrC4cRvCb+l010
r7Z8Gz25tai7KteJLaLtWOvk/Vok4kbMwQxAGd/m3uausMJIWLVq/69hPfEwjq7c
TMa8zBBfVBpghkT+Goy26vfVwn0EdLHMJe35TQQS62t4zxwr/T3fFiGw4NiP6kah
7jyxHJGAEYlc+dwtUiqJVdkv3JaKKIhQYorpW8t7un7MLMeJmgBW//EivIcS/0Iz
0pur3GpNsPou96eGRyiz+CY/f1Q9qlYfT4R5bAzoz+EsQCy9O88AMmtKQMOlmKds
4Ph0Czfih11S+XFn+gnbudeRBQM5QVpSkPdaNrS2tgEKW2y/WDgR5tWlKqB4Mnh2
vn6z2FagSedZrog8Ct8NqJW2f0zSahNpBMmA0RCm2bHSgHGb/y42y3np6PyzmZTx
qGv0gl/0j2VAChy98gGjR89okkZM9FqXt0ZVbjbzbXMwOEdJRHl4NpncpY6beiyl
S29vm+gy6KyBDrroAEUQYHe/CCTr1KeN0hH4pFSe4O4RW9F9EmEExZPnuj67mJTP
xi63jftl6VUYP3vcbvRJ7iU5442ZfqADVmEYjhbuUDckE2VweuGcjezB0bqysmyf
qGpTEXiH6zFxawyLZRN9vVB7fTE7TMgq0mI6gIkNwuOMuyNepQz1zxWhozXFqFIr
gNhRtLxnbzrrq+jtkkoaDnHc37KyapkoXLOgbgwBjjJo0ci+xUUjL65K1+iCdiLz
kEz1+mhuM0T6OqGbjYSxmmU+cxX6sQfQiJ1QmwXOAOjTI8RUx6dMIIz6tSfQkyt3
HTQCX1WTV8FKP34fHCS4ZTJ1b3m5XhE6uAozzyNVDyeTAUwKJ2L6YRZB9WT67saU
xRgPikYg9lQwyk4895k38Od8u9bq3+2Q6LBlMf/FvI3bFAYmpN9UUTXxFABJl65O
LQ2fFsV40DBay2re0aucb8hiQ+2tzWwVPvlNZQB4duBfKQ4TSR3HM+ZqbCZrVgB6
VD+BSYM3BKKtVGd5SX8mThdbD8lt0n9uIIuQdKnExG6HS5QgzNxHBJo4yPeKmEfA
s3Gdut9SpaRJ6gRhhICRryZMyx4wQBoLyy9EuT5tpKGDBeVFvSmkauZHEkogX63Q
i4v+hIdEPBRDbha9b7dH1eRl6ltfV3Hz0mmmBxz2OuZJM/A62Iu7d1uch2tpcyZv
Zox+vg1T52NvcBNsTNI5cMYtfWnFQOI0vwNjt3AB7V2pjt/drkvpTsJBDJATsZo+
FTDzXuGxV4hviKl8LF1ecCLiax1zb8XMgbI8GNEeJGSKEkPtyLBEWxEjCXI1XJkf
VRbBFVhOOWf8myyuhebfFGB4ScwQtRnDkKfWxM/RFgwt3pOkqHu0vSyClBU/6m52
j2OE0I8R9UEvzC9jSo+lC0e9nvewrP3UhsmJTpgSkmf0yJY9Aff/XRRG0BdjC+FX
re0hmsHKDVUL1Ud/DsMUJXoT2E6ajEJWf4E6GtpEH7vqNqf8mF1uaLX7XXoaDlNW
3jTa2QjIWmqTMduk5Qzwk2aGJoSd6LzGtzEE6zoeQ2J1pbk8iegAnI7tuYDeljiU
p5hVSJiSEg+kZV0TR4X2SzxqqetBtUsWv0NEUdHIKR1414qQhtg/JoVdMoTWg8Ir
ur4SWUwCRsRWzVt+zK7oSuUvyamGMYq4Yrd2Jeh0fCHel5exjp4dWQs3zLopp4NU
5kT2C8mXM03ft3WFeDU9kBYLs5kAv2zXwTBofj1Ad3WzGy5HGDRD5d5HxnHSlGcL
kKn6D2utaqpeta7UgOqfYvwShZfKmr4aMY0mHfl0qzqczPqNd1wxx7EV5tKVWYDF
SmbgkCo+IATsUU8zJau0Rgm4SkbU5GN4VOIo0iSF6cHGKsGDkbg2qsXM2KkAVAkv
szqm4hbSI2ztWZHfgw2eQub+9piAOk5PRxbuRdZQQ1shZcwjg7dq4gnyvWlngEh0
MPR3ZkcfY7gMmqh0LrSFjnzVfAomYoC5+ev1L2QiwktAJn5X4W0xM3c+PuEhhaJm
aaLzOPkVW5za8dVZdlNTNAVbOeXqKbNY3PveA8FFsKMWmZ4nEtsDAavX+8pVWRGG
G4jZuHSIe2sD1mUoPh1GBXO12wloLsr83mJxn9p2rBiRkqj53du/dDufRpY1MzSZ
2UDphpasz9oBSVlPK9gbhDgmg0eeGrn4nJ08XesIfNyturwlDlOMvsVdHCZm5Bfw
OnrZpkL3keuxc80I731T8Vns1LMod2Ma6GRniBpqQ1SWYdrB7fB2lGtxrrHWBIGd
lJB4XIMXih8ygu3O/CfecyVadj9MUMWXO7onZK64Zr3bmKzBR+bfSchEJ1zDnO1x
YzkccdSBaqH/N3Pzp/C+XbgSA5Gr21aUamipA24kjJOtlT4+Mj+3WwkFxSbOqdGQ
8MuxBvkGgeKGcJCH0usF01iH8vXQ6tBnuPrgBzy8k1KIoQImcAtDta8lrJ8JU6uW
dzlZmWdDSGCvCny/lRMVVFiah0DR9BTxRXLSbydZHdIF2w2MTcNh/rW/71Z/dfpd
ggwGzF+wvYyLrcv1jsKbFXZHO3kBmOugKC1l3sQ8HFvbOPZ3d4DliSDilUzGlVky
aqVbPXTxIDiWIldHFkDir7DHd2zkGvydbLL124E4PpwisFf09HDIugNgkIUzDLIP
8B9FpfoZA+6rrMSS9pmmAodxJHCpBV0ZZ49sqG2ATWjK4KPpgsqXBWogTauP3LZW
oxdYkTU7cRPdXo3TdnJ8zHdgYt5BVHBujKeeV8ls3FlVuUGrQa2hU6dINRb/7qRs
DeqFq/o5taENx+VGQgyCJWJYxa1KjFddV89vg0omqNWPWGdy898Nm8jwBfHERr+I
EK/D8Wg8ELmFQq2EDI+du7kFaxOr7Zk4iyp4fHQqc3tQnfrTUpVD12vH3Q4xbIlg
tthFpJdQfyJir+3UejnUZCH+rSkoIUOT5mcWoAOyoW3DMHg9jx7F64QGfIKIoeAB
uLspcAfPHvvYuGAa3bLl2sxh0fHHkfLDMXx6VeE1FtodsZ8uLcHsG+riqlA5TSNG
LUpZNxKki6PIxcoLBtczBIbRzXNUNxHeAidjh+UzctVh4lgDuHrAV5RPbIj2kN/C
RhdZUkSB7/zmTiGdSA6nR9v5Kx5WkVIUshLu00BGJ9O/n6uk7oaelB3Upph7txys
VFmIL3VMLsHhNC5ftU100PyV8e1Zj+zRfiTaLShYujXi0V501IR4vI20Ibkbeu+R
qELw4Qm0auNnjS8q/LbcgTKuLvQ1gRoeGx6HdNMIqmhvt85RwBMvDBqvF9qUoW+l
YduNSahhMzSadujXja3UT8erF5jNmVH80sJY4JlSPKo1oSMwcGVHomrdZrtn2pAq
27+2sfkJ1cf6+uuXkYCJPJiUBWwVkWoGgs/+h7GuyWnOSbwvBEd9CH6lnmYfZXBb
ss/SxsjE57Ft9fdXYWmW7rhBU2PWbybpuGqJCfd5rlmAq51BOyMR/S/UzLvc63mk
e/F2hsl9gV6QHYbP9uScOY+p42FriU89ePJO5h9kd1AzVfEwi/RrvHM8/M3kNiHf
silwRhS9+F4ermJkpbZqkQlemQSkw+N6R419O4uLbqveP00P/TGAs9QiLt+hr2Qd
w11ygwRVZdj/eAt6URQ29UYjyTnMuiUhZJKmPC4k3gRIAqUjoAXprbu2u4JNxJFo
3OGHN4IDntx3JmSkhIpQ5bqIpCRHmv7842EPkFEwHmvTabAtB5yPvscppUwFueTT
r15TYIivy0glDnRpX0sTfTbowG+/jgam9IxRZ+idKT8WIfc8J7OYjkUQkuE918ws
02pqTtWyblVIwas9GQvmZgv6IiISxwIUog+KETSxAU+o614Vaaap+j+x/Ag5NZun
2DaQfkmV0m7E7IAwuCrSCwOt0ZVvE1Z9RJFDAbP3QkVq5wn5qWk013eKXhiboi2T
xfqcKGBt80BUUV8ALmAfOoXkKCjCtWRKujD1p7/PAs2U5gJjOx1Ot+Lw6PxOzNtI
+K7dHjJpxa/FWdlarotQMxS0DCf4k9QZ5SoSVSg/fCkqgDVDU/vQ59rJzXtK7fMv
lT0aZoElIAnf1Ip1SKc53tRKbeff9SoshvJZIM11NYFkijVsEQUO9cdds/Ixse/y
7lvoN5tKGDlSfKpRK1BwbLs6spCuZQSkS9/D7ZhT20baiSzUqOBFx9zAgZdaxZGq
J5FHKrSG6or5mlbw7mc9sfFvMQASC8f9ugMbVjmk8YhvYPUgmDRblErOmFMWfRGf
caeuvXf7NSs7kS/XlCMvGUMDmBkJBVJrg4g7dCN1jX02lASSUbMwcU9L16657qM1
KtixKsXuHzyhlGM3fJaERG7t760Ik/pHcmB/2m+XZr4LFW/YTwx3v2avSax0t2bX
8wPSLzbUOjdkwNiXpVQT8uR+DvyDBHUmXdZrXWRrPp/R1VEB157c6pF44bG9D4v0
isu1vDz2ErquIkrgg4IA/OugnDwtgmHdBQS4EwA8kWW+UOEg/U8ul7df5DogpgVT
BzzGK//abQ1MmGSH9ru76YMjEtoV0KDBO5xfHgkVwpQPOCQl3oNG28rURWJQ8TGb
+MTjrtDERHdOxncpK7vg1ohHa6SZtocjnITJ5VSHMayDg5K7h+hRDjPj8TFJgg61
1T544bpsw3S6Ih2COkGdBD9nQeYnlzgJvUDodEqn/5vNHt5R3Xe6zRRoXfyU1Zu6
L9Bb+0/RcCrhFHBoE8dXWUuqTIppGICqZW2e3wktDI7ek+oFmJAuySj1hazp7ez/
Ivk2WetJ+3uH50HrAtFQ5XQh4QEVLOvCwk873j/TcekOjH72pVk8T3T2AHxfoOZq
pczifIEsYPheZeiRSd9Yip/0Zq7e8pVeqWtAGEnTyJxLlIiOnFaUELBrTdtZxkYq
KF8Il0UIZml3tnB3ZEaODYiUxjbvYHMIQZH+BBku2Knh2JzcNX3r7l5wy2lYt9Xz
hIbK/qDEGa055lwLj7Z8Io3b0U0PuODm64QgWiELlVwnePEAQgHsRFogU8L52qCN
PXIP+45RerNPGklQcLNucnWYcPDSDcXtFRsDZHaQxZ8OxmRM0reKj39boTNS7pA6
oumylNEGmS0gJo87jGbpG287itq2W+vRbyq6XJ67s2aVYHOjyb+BMs1sStUKXR1e
V8aE+74Op2OxcdxzqxC3C6XEP/2PayFbReordRI+4m0tBw2kxR9UHZ63xQKWprr+
K/I17cMANksKY7wcId9lWY9tA67dXPTm7RFJ5OluksS48xTEpe8VQGLwZ+ZwghFH
NBM6TwoqkaXjpFVicKFWkXRTvXVOYb2W44JIAkxhyfsbYAzY4475D2x/ej9C/4wM
C2qCmTwEVbYT9IULGgQCn5TkhfzR2XJ7HmF6sj4AtKOuN1X8LeYzF/Nf+mrXsZHY
j/Nz2MIy+DN9QtKXtQUuTnIsHeWoF6hI6wvryVzL72OwMfQVCKesAG4l5gS2K70r
pW4PUPlVJdxU713ldjsXSKWbu/F18HDVm2VdRzIBYGbV0btxqH8NrLxXwwaULU/q
q8u960wRuLn1UrrZK5R8KrjPgDpPqhtINr5M75bo4K7CLuHSOgHwhqQz42RAiPwZ
QUIrS4FCN2+ybL6WPfXlT+igY8N8dpYsQnvAZPvTG350aRa5y04Q8rKmmJEA6/8J
nO1UxF3br9Yve5Uj0Hh6AEV3sbuhszSs04cjy7YAAN2r4SgywGWa9fV1QTdIOhTL
e860Uq0iefll8jP+xDL4pHxsFp2Z4lm/81UDecZKSBo/kMwIYA7XY7PnzKYPcvUn
dlgHf5UjWt2vpiszn6k3ob84iEyrpt3V0RC2jTwteIlIpHZvPIX38VWN7gqbmaDh
4THq5xnC3uYXBQTmwNVSDkMFOeLMMV+hJIUjpe2LXF/WWNmMRUMlcKFsdTQCISTz
k+rxPAvXqZNTgLcKmaRqQBOkouIYW6L+1jmte9G1xvED/Wx+62WsXtCgQCwhXhXo
vltd+kDcVOK4JZXStSzuMGAsQp/mSjOmVMe4HfZ8L48zVfIm2MX1stZjqvt1Ba3G
N4OqW6i1eIfFOD+yR9V5cePShylMLsPMnZfk0eeQ11F1Q9uVL+hFw0mO7DomdApf
QLH770m8YHJpP1iDYTukQq9WyXUGfQr4wxm5GEHZ9xJWPqFvX+lrx5RU4XlR/mYk
FQ/o1XswNBitI2f1Eghc/fb42xqcJrsPwpbkTRZRTeC7H8HCBajeFcYpHTxhjS0Z
SUC1UB+YiP9WCdhpFsTa3wFEQnF+WWEB9L5Fntvkj3xzoFYie5Rgywdxz7FYqWjn
HB2bVdW8LctvGbG8FQsWND44Fxc+0BLILlgODLYJeuV7GnObyd/7baZD++OF6mzx
+yxjMrkFGQu9mWTj3A35YAjVFQetHx7to7W5W8zw6U/n3Tfa983jaeaa5mBoEcSe
YG7okAieWgxgWZtcUBykLr6Ef1/qZ622DQMHb+Y8nAVvhkwaAMMW9wQch0mheMRW
FPFi1D2o77Jfqh74Rio4HW6QiWnWB2/dK6eZbpSp0WUFNaLKp0GudIuaSf4368Ta
9ICM/+2sVoNDpUiAckjYNJQb8cnAHHqFufVaIQ4ZdKsIcdambab/jLPaLTQsCv2x
muhNgFfh0SSYpYt5vUSLdxh1uf5HvOWpQjtACwm0QetURx4bPJ9dcZEST/fDqTPb
z9kHVJYX1Cm5K+NqXjEL0G58uoKEYPjVkslRMRFIRPX0sAiIKs2jYMzldf32VG1+
h4Q1hMwm3b+eN1DQYygsBkbpmrIUB3nuxe2XAxFnNBn9iSVxwjKXkRd3/F40fh8Z
2MYdcaKU7FmdasNdB3mMsMXJckgkEggbA74aVdTJJzj91d9aOYDSfMZF9AWlJJV7
GsQIFNzlXFaByzaejmO1eGBuWRuJ0UoQv0IY74V5zbQmpUlYviB/vCGFApdSrWj0
T0Vc6ihme26sFlIxPYOxQRCyEA1VG4nisRjTAl0OGwydDEeA1Th/Bmf6TVAMQPfz
dICnG+4tqGh0sGRSIo3y0lv5g4qjSMh3DM0Pg2ZaMV+KW+Ahre89SET5uBVy7LGa
HQXkeLwhDTyTSGE0v2Qz+KmsVfil8KeGaxAso18tfQccqzCICM3Hgf9LVJeSizS+
x+BksfY0p8bZ8FYTf8layu5SdrC/T3QkA+Tpam9VT8A7MThaCVJSCJ5ye/ydXKy7
cssRxMo/JCqbTboc/9z1wXaYYQxHd6YCBwTihbB0qW2cavpMyzqBUCYkyBWOgffB
kjVzFqn2yW0Ys7ESFD3ZOhgfmv9FroTuUHC41YJ0Oa8qRvjU3d1VQFMQ9SeOk3dG
MqN1VUAzs+2y7bHoPlIp1uk1/bPrLyDUdVXijHsONva9HQ2MZz4rEXXmElDZd4Nn
XyLDSsm4/4GwnXxwa5R9VYsctE2LqYHhZ3md60P90TduPQsMY//nQJwt2/HuPoev
j+mVSnWPK5kDp35kV4JdyLg9Lfj/ZuQubfqoDjpDlD7QKFUpURnPQlCV4pFCtOHo
m58nr1LHGouLdcA0NDrMuy1AtTbhTqJcrV4f8OYrF+71Y6TzCd90vJWy0T5S78mb
fYf3dMGHZG1Uvk4Cu2HEKjYNVz50+ZTkIq4+fmV5Da5GH/7ztCCVbvhrczvxBK2D
7VSB6f6b+TLm89MVIvMRiFgc3V0G+clWlhqyL5z+M6wsjt/mEYTSxZBseAMBVPiw
jKiH6MK2P/+a/4lbBwWaPRjxyNg/ekLyYZ7oN9wIwen8rECbl01vKfRuXM0DWtF4
gUr1kOaikU861mDhDbvR52DnFFGRK+Xs/hkYHnQeBsmtIFjn+mckqbBI8x/MW3oW
qliFYV7bNxNGks0PgNJglHvg6RogcZ05IQsLdaq+ckHy5XHhgAS+yA9TdRL+M92r
h8uUCZ13VZbHzpTDc1fAQSB0oqE5H7p63h017nQsBvPtA6qY+l4xRD4K+zkXWqtj
r6l8Tb3yBhlbDVZbW3g0ZiWLNuTDR9M6IWYoNnUdVWA7LiWxP6F7cgBMVJjwfYpI
e4KhYFkEkeZjbf5Pp7iQm3tVLpl2v9Ef4x+rUm9nq5FlANWb0qoVc2/GaNsJgNGw
JPWaA6zb16jmq32CsPY2ZUQF04k1Pa2tqtsnLVdDpYVvcDqVDsWRrzCCpDXDeCcc
utCaUT0avCwp/fnSa+6vOvjRw/+s2T/AEAob5sUTaDNV7DQYj7rflBPswZrCskQW
9a7bjIxe5w5zUE6T+MtgtDZ4FSnBxA2kwpRLljYA1uWpnXMONgO/jnDlg7gLe0E0
Q1G7C5Zq92jBcTXUSRtmvBR2xhySbyopwy9htc6f7Hh9bb+OgsUCKRfw4c+L7oVJ
l/u1POSkI2A4ROb9+B5L9+uyi46oDOaGFsx5oMAKNVjVA4KrD2ujJh8NjATzB3lF
N3w70J8QNbQhkiWDNLTNKGDGJvWqkCRwRnvtzvX+05ZKologG1dyJh7W6GyBorck
I2U7mVQzUNQ3hrLKxWyuROh8/O4BiMYVtufKKoKLUAI0MTGKvW15SXkO+AZSvi82
i2LA0bp95cetNqRjQZ89I0B5YZYQJiyHyPSfRtJcivANKiYCyDXgmlIOMtS1PVNx
Req6Dr0izfPvl4/Klg0ozydeY2qkm610lIJrxv5WVGP7IxqidalJhP4HSSOZJJrA
GQToowDO2uV4p/Y8KKH2eW/99MY0frurUo3dBLMvU4xBmajGIFd7XxeMXn8f8DnL
6MwOh7+rJbSpzM75L4UjqK6gKVt9i8TjLI/EzRsr4pmz4nhc4QNReTCKuPXurzvJ
IN0JSGRUWHDIRdR+dqXUn65Y9xwVLssmg+cnwXu3hT0niB4KGuRqikN5xX7BMXGP
CABFaSgKxORQ7R6/ipgoCrzPBau0vJQMWMoXsur7u0NwjVe3n5Rh/TGUqs3s35ch
yFf9TEvuFbkjNt/YeT67Rpg0yYyJRkQ18pcHvI7fd4wNvznw57PiVc0xYreMR9xW
feHRBbqphfi22moCBTctNKQyZ4t8I9bZnV5/xOLLD3ytcNN5pAgA3HA781/Ed9nv
YXI+N2aLW3R1Fzqw9X+V/Z6fZdUC3tuOgZ/85cX+hx/bwJLQNm0IvjL8QYScGzTJ
6E6kIRE5cldHyZ4Sxoip0P6JZ5PYX35yZSWq2S76Dw/Qz1/8Ye8qVfJEhy0Yh5Uc
uwYhl6ijRKUPU51OGQ9OEz8M7WyI5kDt4ujy82ggh4aLQDbcrGoQ4Xvt11bFxgFY
y+415wfTEaikJ0HW/pM+77qjzy2KrwJcedq9J8yaUb7RuajzJ4yzlcJ/K1blVC7+
N9QZy7p8VubhauLA+YLS1ncsNKzifo1G0GCHfNrhsa+GwCg4ASu20+oDODGXLQl+
d/SBgkGw1Kx97Copo+DT23pg+4ssCmo/McR0QLYe+bo6AbOjI00Ub9Mejxax8LYJ
z/OVCVDvYAxc6LgPuXPHdG40kNixtNticidHc0f0TSICmpU0BksvqDRC9YXqmFuG
Pn4u2m+xOn42BwJdl2K56X+NOMQhsSimTcMtyFkoG1d30bSNvT4RK44HJkfhBCKv
qUwChNSNri42UtS2GgDuWoMhcbl+CdGI/fo+/8Yet8yPp9xwbBkolhSa5RkopuXq
NUv5gKnHxNm+WWU3rWIGqKdt6Z1aUo0UFkpheQFTISTKYpmgicVtk1jznrMfoLPh
KFmUxeMxB9IOL5M/LrsE3a4dFryt7fmAvBopbHiONBTPQrdAeml+zAC5bjjN3nYP
ambC8dRZ15eUwdcPJaNA6NY5+XlL+e1eVLFa55kKwLDYUce9l0lgiVpwS692We0O
Op9lw0KqfL49E7TGQ5XvLA4xI647rHQ0i9pB5L+Wfq/Et2D2gVAeH9MN1H5CLCSc
s5+AajrmXUHhYh5hmpTepzVs4U5ZKd3+moSKWh38vnHuJBL1Hrm0KYQCGJfYdb99
JLjgaXTW6RUZ4+bitv1i1dKyEqngoiqUYEznwTtLtDeYB+qR5FXVTjqp6frYf88w
3u4ZnNB9+8YeFE6GwXC/KE2VHGn8HgP1zyENUVlo9VgihbEj1BZqaauw8wn6skJX
OKQ58meGggWTPym2iZ+SGwuIRzIiE61Lr76V5THMX96cbsbJ6MALOJrs6l1XY6CQ
Y64wW38ACkZZgu4OZ3MjlpgUfuEaXh0JgPZ70hqzsvflX/wjg/krqZnvZoJtIwq7
Q9khsi2iQyHkRdikOIay8aXog9bdKYUOhWLj9Qs9KIxnZlFRiyV4HRGJcUNUpwGF
TYlGdjJf8vPb4A+lj0+FOwQ6OO8TFJDdaoHaN8b5dXmLRFqTezjI8RmPTBLhIH1y
DLIQp1qFGGk3oBwYT5mlBwLNN0HG3dh6oSAiF5vgzsrHVQ99fFm2Sd/9QkTvLH3L
5TyrwxHHBF6Zz3noZ4t8QvlugGjCOjgRprj0DHGIYG630/35tOQ8cBi0tVOhY4KE
ECqvX7SFIdBGQBd43Dti/x8wjYdy5FpWuq+5H1hvDRreRXw2+T3vI9vwhyjK4m/O
dgeUnT+Q0jUt/aH5QyH2kmnl5UY12jghHP4QZBkHxHUSNbRxSj+ALLVwRtfL8sMz
Lg9bRqmAuSytDbADRJ1/wqMUMrbRKnLz/FkX6xEytQ0M7pk1Wh8bisdggTWzWsp8
RwRgVka0+bK28Vqo2iXxn0Z6LZK867OU3+4m37Tlep6sRvlPT2tmhQe5kf0CztD1
aly/wZAiCBae5RmsB5wAkcqBK86K30BQlzckpz+11SpgbNcBE57rxHPLrwg0pBhK
8FGXgUT/4fsqMXiaKEeLnbLQt8NoM9F0WZ6G73/OK9wMry4kkVoFt2Bv0ikkCgoq
+du2b8tVNcwi3KHcq1+NXDGFAfc7pmv6FJcgVXb8bIUJpGPqrK9I7JXe5kLkTwA+
wqExH8lhIu2qysv0cxkwveUD79LspJkygk2vlYIvFlwE/Lw3n1OHAD78HyA5B35X
15SkzsLY+vfU0o+JWm/ZFD65c+CWwGcTbR0jYBUJ+MdtprKxzsDNtYCnypX4kZgY
+hByZ1rgD9UwKBlyL/Ka5BzuSTa+SoMBgupI4bNf7UyHSJHjslXAGftX1cLPGPw3
bnV08jCbwCCd85K7l0V/1aeffFXft4nKqC6UHuGrLHZzz35HF7bonDoeB9PiPatm
c1s1mlpwl5TxUrC2uw36MWLt87ntdAInB1skZXHJQcZ40x8Sy1DOWh1fdVLFgx5/
6X2+nv5vIXF8Am9N7S0SG6jqzS5we3VGOO/m+jQn5j62W7okXhYb73H+YELrjcnM
HfheNwCQ/l6XlxhMFTD4UUzmemiTkOGENLRO00X4WQ4XDhHN5FjTJTybvgdXyMPv
fGjx6FukMJyTWCxvvvsQjciXKmqeRYT8rM2ti+sEW6BzUqr3fo44yKMe5Lv9SZSc
JWEYRDSrZiQOLftCWWHjCzpVTkv9xQOK+XepCWaiPWyO0RMj8MKjJbHeyWGeFzxm
n2yFZ1WF6pv4I92xhE46Mb4Bx5YJ5rQ2Fl0EQlWU+cHGaDaHHN194t7uVf+Xq8U7
txAlG0yACUtrHFUWFvlH5sZiE1x8vNBerBiAj6hVJD+R41zylDcEemvuPTfXVH9V
Gc0CFlAh5HXMZPkswMFsxRUtJ2E3woldjHO2O6sAXHWDqlxmg4hqq1Ba5qiZtlym
8wbVS9uxkQy1v36//y8v5i5JbOY+/mVcnXHBKz+nDnQWcRcFrrJzClOTHvRoqnJI
AvYaVIcpEiakLbORe6c72l+dKN21WTqDmMLkR55UOsVC9IZeoN6c0aa74H8E4gzL
CVKNfXbIWtXQePWgzB4ziKK0jRd4lfdX3OXn0cZxBUKm2eXMaUHrW7ni8tlHSpRI
Fr1NJDBQTaw3G3YlMxHBH/U67XCqFBKgaUTwLAqK5fVT4yKFwtY4NlEIqOC0B7Mb
cwifpLjh53l/gf2dnZFfxBZ0jmM7j6OPVAiwJqfR8UooykFsd05MK+wet84hPdZN
N6/9hinzqVy4JNTON36mANr6Dz5gJ+NVacVS9avWyz/9ZAUB/SvoiWsYqHeKW3p8
D12dRZWOC1m+AMeiwNarHKgK6mPUp7F60wYmeg6gu0mi2QsHavKR7tUCIt051/gy
vRtvoc9pTfih3Eyv5qG+Q4aQqibvzU4AaNlrDUEyoygkh4wWFbJXTeHQvL7XT2rY
j4yDcFPIhiG92rn7ir0JhsOpGNet/QpC9Kh6VCcCDaFlp1Nd1FdCvBMIjLdMT8aR
9vcCieRhhUWAtm4nTx70rPslE1ND7iKEa4aehAZmEN/2bVlrCXaEXdB8NCdj+Uqp
bZoiPoIjDGnJVmvgHDDjcFFljfgVed2Vz2B4c/vAYAtqFbWPrHMgIpg/nxDvY0On
fhMeY369H/H0jRKa5WzI4tIHVEJ0rXybhVv8x6WsECACF1l3tb0j0h8A1fr/XSya
t0jGHsoCjcEYI+wWgxNL7vdFCTi7oOnFpyEyNfLKIwk2DlTvEfcNx2K3SsTx2t/P
8OvDNlqWfDQnXRIdArxnWDLMVYsbOHdxe0D2zQxx3qDgeNrzbiDGtq4A0KD06emZ
CYiR/CqkxdjduE921b0FzVCp50MsJqmLb9u5GemdoipQr9Kpq5rL2vy5j4pdCZuG
/fjs83X1YiG4WkbxDmXmb0alT6rYcSWXCKgpvGuHBO2FeXLCV7FGsvTEdYJn4Csa
GokAx2zNXBNqb67Bwkhjkxdt4MM9pdrmHyFOw7szoT19WEE5hPrvbzJxSlzDs1PK
i4HNUFufoIpEbVHHo4UmVX6164QFgPzK5yHpjzYMe6BqwSvyiw7i7KcCAPJFMIug
Lh/jdgE6cegUb3T5w99JKXRU/cXAojGrqKi7WQS6zpLMH1L1hmrViCktWgublLvX
oCgorEI9drAHaQs49hjrvV56yTIKshBC3mI30U/lon1qGWNVV+LsNzSbza8zVmDL
iCg/XkcbX1awb5k4FGPc6KYh1ETpqEPxG5iRk+IMnQ2fMaaCUhJU/u8VeaIsvTNy
IGPF1FodhtcZUWPRweo2Z1xhdm/GXDHbLY7H1w3cBRF9uuGqYdeUWnblSxDh4fcY
OpklFKjUBBE5VRO2RFyOgnejHsHVJ+GZR2gSWaqZXYUoLHcFnZBuvwR1yG95xzBo
/mpVQ9PWad84vJzorB0tEo9iDPJwXynHBX+tYAzEhwKD4ubG5/jBp0gAJNltCFj+
8vJuPfj8lOZ1f5oECzVcC0GirPnsSO5E/OA7tN8sjWm7Z9C3OmGjtYmx3zilUzNZ
pyslRVMV++Ic2vRL50mI8sdcdShNT8DMVKQXueHKIZiSNQz8opm61npaaRH97wVd
nSmwiDkw4IFxDZKq0pbmwxaYopJUiR7+jXWmIST4NjrkETEkFTrkX5Td2wtlJHNy
VYOKDsHq7RG9dklw4t8y+PYBrAco5vKoKnLFlEE2+3EiVfUakl5R4QM8+KByNEKf
z+SJMXW4AqyoC7swUfvRotLlf1wWDWEKhOOmZlH3IQMyAorf43XIwNfWvk4SEAn9
bbgFhOAiclR9KrKBfoK6jUhxamRO13QTvFd15AGonJfbuoY6PHdY7/OX2DG2xo5K
8C0uQhgjcx2Bk0B+lBWN1U/ldKNUpkij4bw5biIW/1XGlqurFPCC+ZGnvppsFmKw
YgUShVC8i3ZNbkO3YEubAVRs2BE0I1vPCUXsKZ3zRO2+TsU2qU172jd661cJe3iP
L6L8fIXD0hg58fxpB8uU2c4gs+1xshTsqxvPRuvVaxZch6iuZtrh2JNq6/b/e3t8
BAFviKwwroJ9yB5OODuyr0s4u8mxvQFQ0jgIIzXlLeRSCvJxFTnbTyP80NXJPdJP
zqpZ3wJTJCRiaK8DTJZqnbgXSNZ84hgRPhlaAIn8yRuFoWaUnkftpBT/IYKFa9DO
rAVWVIyzZeeEtVYt5KU0RCa1pLw7H3DQitb/KPyp098p1XkryRCFXlazUKqGAKAD
fGLF/CuVMyNPt3aGrfwj8fyF7bZLsl4lDBzj3x+JawdXHR90LQCNf5M9SHH5jO6R
x6K3nqvd/yGHsPh8CAJnVybhUJ6Q49r0nnfgEDF3EZOIjgyZtEtx5Jswxs8gED1U
ZFeo+TSYdRCsRjAiZ8cApTCFskelQ0c1lC82IhSQyoJP51QTRntGdARcGdvq4afd
k7r71K4/SlOORC/y43ZIVpHH9eB3DNsODt2geOEzbZZdRv9+XYNCkPhYzcNBrFVg
zY97jy845IwJI3E0MjP46IlE6xqtlGfsSKp37VQM3LQ4/vHQColpPl55BPrHEBSO
wszmm5kYqWm1IGMMzQ27kIIuIgLbxBksOidazwGDkXBAqX+R4FxR/z7uaMC/7xLa
pofEV3EGCjmKOG6AK9du+7v2wieLnPUtLDzPj4t85EY5dytQJgZQojCi81NsQzvM
uGG9yn0X1QYAt0u4sJs5Nd79eQ2I+qOUAgcSI+5xQ4LCucPgxWDyBxd+7q2wzT4b
z98P0L+D48sF1xQPKLWL9ttWjZKQXwBaUacBZr1PfaqqotxXoFJW9qfEDIqEUy80
CfmhmiOLq6ayDLRdVgkan9hcApp4VwwQzkv8LaBacW5jQkdLGQfPbm6273ZxxW9W
56gPI1NzHa78NLLme3d0WkekmNz5ygeIt91JAacW/8EgqdikoEeWKwpPHzd9sg8E
y5rdD5SUueZwT5l4jWjndlX1iyujF9T/d5cOCF+O3hk8P/ue89Oi7GuFs2DOmoMl
oLsUzCCYglQerNZFbbw+eMROsD5J7QL1THQN9i9yiZJTLox0xo5hU+fW4RZgtJDV
tplZ4cj8DACvpFaOR3NwPV6/aiEE3fyqmRoo3bi7tZzOOOHkil5ft3FvEOxaB/ID
2HKtfh/mNzCaBnEKU7SXsWC4lBJzKIrZ/5R/WCsZiQdCBCtRUrU5kTAgCIc3srNf
WZ9xs15Dpb5rdighopt8LR3iZgcUQkEtrWVoJI2fsRaIMJ01nb5nVSelf4XcLMy3
fW0eCOX52ToLOhIV8HwaJLt9lh6yOZGN64GKJqZEYPz1NbIprp7qhLpcD8t2915F
LYIyAL5CevBID+odqLHqzsgAt8Buxy8sMpgBUjEI25qgY35hfLFrRmkpBL9NVoIA
Pd/bSZt7otWtMsQHbQunnbBM1iSnzhwVcqKzSHDVkr7YnKLXwuqZ/DT+ANF3NKKw
/w4770b0rRFl5lAu7INfx494pYgiyYpnT6SMJpiV6S/0MOjlaZU3fx2/qI6uHnPd
/vIrwoUFaYi3Z81yXk3z44fPm4WZIs2txMYUA+dKdDe/RgZ9sNtgi5LC5/kZ7uwe
97DKdUVCiv7vQfDQOJaECS1QtgEg2x2b+WgX/Bbw+VS7/4fmsT0FqY2B1OIXJIQX
pG//ao4xsfIC6wDpfMzR0fKcVO1rYtaca/kpo6iAZHL15mpN9X2pgM6C5R4SMlUH
SeBLx87ulFggHp5XxU0vDpFjd6ryO7ioTW9HMUrkEHV6i6mvncFNtzoxgp5PKDsp
tZ4kkFc8GitBMlNNQNzXBPjNxXf1ddkCaiwEUNszuMlo9J8SMU9OY4ID2ubxDZrd
E6I4dqdgvIFaabmNQCTyC4MR8jbDKAZ6bwAP6i4t/aubYkDmZVniAHnFagxeK2zd
1PvmvF7ZrqgAeGQpR5cQQe84YcBawGhHQpGTKQPXFhDLpC5vr5eaQRqco97JmJri
NFGOndCyEuDY/MpWw+dTd7rTEGIBNyEmE2YVn5qV1ebxDXabT+Ded1Uj89KoFjue
rT/Vdwm18d5b8paHgktGUXh8DzmB0VE48gXSMg9j8Bazk5Nt1QX2tqyvuRuiAElY
HFqpYgH09Z5qMj0qhGgnYkwo46lzTljO98l4guIkwJtNB0wnhb2BBeZJ653jEqNI
adhsK1B16vnaNdE+woob3lWMEd71l+XyqhN4evfp7s6Ql09O43MG897fuJJkfBt2
ozsJXmLIEOY2TahF8dULXkLTiyQoClKSaAuAc99I66rlkgzKMKQYsZ0IAx8bkEpn
vmjdDZamJjlGsEMEkdI9xy1xuyvsuDMVNBuMvCofmRsOmYK/IaDp+ojKDTd1r0Hk
XSUH2T92Y/Hj8wvaL3et/eQmZXM2myeDJVmAU9TRVAN0qGqqdaZILtRsb2YvPXGw
lnVxatuUic1scQk6QBbUMUalA9L6kX9ljRBlE+uHCPwC7zM3lctoAy/DTwC1X67Y
oQWpW++3cVMD6pAkemu3Qq1bT0WyrYL7VBoMXXqk4TsuFw2qBoyROaR11esSEcCt
g7nZC3B2aj2pZmxkfURxIiAKLmyAyWwqQpu5Dcmg5yLem6h8HULFTZPeg9wzRJUN
bCRVeJul//Rnz+p5NdriYbJ7Q2Ou6DcWFkyjjmZuft3Isx+vnZNweYvLhxxU+5Fi
K32ZYLRN8ZWQjFvBfqpoTQK7VGqkej2jw3Lx8AR0ssudY0esQgnWpD6+L67kAcAZ
gcopje4ogZTctWPFPqOE1PSdVeKYXQPU4yqwVkk590g5R0jxEyPWam5Jf1p8XulA
YqllwdnHCHYJvMv8rps3WeAFSXdQGGnEz5s5zBOkDwheOXUMWyK3CC1QKbSBVSXQ
qtp3SN8PfwDjVteai3L/Cn7FDzqoY2DZ7oTnaGaIxzgfN2AEHt1K26vQYgMQ73sy
rrCI3GmvOJ4unAOBLpGQfb2Nuz4gf0wzf6PCy2cCFjGTGZJ8Vvkfww5mQA0WyVMv
Q8Wha08B0PY9HJF/vthkfbt3RKPF5DtvqylLdtUYY0mYlytie58qb75OKn6CZVBX
3b9/Nueu5dvz1OTxwH6jSU+mFlb3PscIcqQ0QRTpy67eFEwsN4jn19LjELjqZHEH
MAP8JnF0JWxLVTilTSn+jtuAZfGXETfJC5JkjQwobXvnmFrFB5v6VNrusMeJC6rf
yMl7MuCO9c7rE9cPeFHhh8FzrBFsq/wEPDtGyOojcQJZHLE2+pEoq0Xku2ayq+Oo
fNCCL3JBWS4cIjAq74SAmt6gV+yx+m9WBUdM77WQbtbrdKO/e7EOCruP5mOx/6cP
kvT4nYHPUBxFWmBDdhFKJmiafY76PMwt2rYAeg1FwQGsoSM6Gzubk30BjVi146UN
yMOERjnsDdTMUrDJDMm5DKSFYyius8Qw/SSOVWbHqee81NX18IUt3flcBl2igT3y
XsWXMiVw/cD+xo2WYBUB9RgEFFbLjsS2vIl7bmqHNeFAx8PLiPrRSR6kpK7xwQ0Z
DJmPPY2ux3KgP6PE1jbu5FPRkAznOun6YbcIekXKvnAdFRWEId9e6UWwdq91IJUE
Cm8SFgtSUQ1z8bwY6NguMjM9vFiwSHUw4n47Rt4orQQW/VYemZgZCw4TzmJahb0Y
YtNUFLDPnuRM49rIBSkSRBhGI8SBYuzKgy2u0INz1j/FM2Khi5o89C0s6V6IP2H1
fqcVLQS41BCyCVLyST6PUDEKNH4veeZmB78EucNwgbQQWjtZAifqmEARlKGSPbjL
/27hqCaumm/roFLr7gKl2wn+RHO8/+4/OzlAs+qdXbi4bvmoGgHl8LvYpxm9Uneo
/Ue3iJHRR558iiHBM0b4ye/RsJvb2geDp2V6YaH96zZrs1PkeJDoaC8HfOWxNSgR
rSsC3KdBsT9IB0tvdYlClUqC0GzzSDlWRAwtTKVtL+wNaXkMga6Q3PCmqSg4Epwh
ZM4NOj0EngJ9RDpARg9CfkbSasWHW3zO/qphKlXZguRDpNtRlyVDc0s5UuWKtZzt
UUN7ExUaNxmOQrIs15UlyeDCT1dz+bpXyWZFrYOJbqwvOhXCKj36WOQTTb8hy88a
I/bvWQ2drsND/hIAL1V/eMHLe0hM+5WeeL6T+yhMhCNsYGbt1ebcDmV+k8NPLREZ
HBWBu6W+gZfJKYXngKY9Cpkmub/Rnluoa7/X1rOeHsGb4XmoAXsIVQfL6Z8RhU8w
4P4TLggT8MoBU2OHG/MPaJpXCQ0dpEETSVUgWc3cir4L+iHXnQLrsi9yCBSPaIYY
SD4CjKYzBAAbXRL29u4dx1B7Nsnqnwo3lN26L0inG52gAtTQkkY8W1WaIy+SBVCo
kWvHAh9z2x8U4PP0RAsKFf4eQGRILTJHxiAPzwG444bM5YM7Kr6mbPCIpY9Q8nmB
dgBBVA4IeE+kBPCu65n0lrlXk860m3w1E5LwhlQA2YLFyZg09xZhiQw242osFr53
H+NLEL0WjHlchD9o15HBm+o8F78LTd6YzuTluGHp7bDDmpvmY6S40+oofP/nea2T
QYS9LSwQzbbL5pWrGkzP1ICwm3hkkiNpOi0ilMji2KCiLPBjSxNdspL53JOIwcdZ
dzExYHHViDgUvxuQB5cpcCufgtbPZuw4abJ4jbc9+FhApbENrXVfbXAcNJ7LnUGu
QTVXv1S4GzwmG+nGMqdcfpbVbCJm1nfPlVkw/aDRtrCyNTCd/YxuBLjJY6vLHTYA
ePARJSC8Cq9acpx2cFU5mfkAYMJ83kZzIl9rsZf8/q3XD+JhOr4Mz7Mdgw00XH3H
cOnnN5MJTrK236PEU3QA6LUOSGbydD+CLhY4ldMfiHbxIshRf0UtiL/vkSeIL+Ff
5z+geDzMYPY96rThvulkiXUrLYLpGWxJG+PzdsIe6MXnkZHvmp9Fu+GJaves9Ja4
hHVOrLibRMApe8y6PjJXfGY10GPvrD+k3hR36yshUv8Sj1+1U04WgKdsU5MkWQQm
5vu/mH649eh6bcz/FoynqmPIbb6PHaHMOzvHTIFOVOBbSIRynCdgT17n09uOfpF0
VgBzR4T85esphbJemEUcnNTjfrYIav+uLkDOESphLlOtx/jiOPm8abSXmepCiy14
oIUTlDL90v+i9zcKSGa4CWhZWqPXv6G7nWVeu6BNscf3ud1H2V1MQ90sg8fyG2tY
95DjaPCxif/bs4LOAczWRVif9Mbv0ScFOWbsufDuTSOAsT1/lvHyCCBb7x0KuiYb
JsmEaqa/OzhE/C4oyQ4c/CmRAqxwzvcJB9hsiC1n9jL++F+okVeXxaX08TIISjr9
677XYslgRqlJrkWMXCSR0OoMk2vDHwr/o6Q7+nhSfZJsMljq8EwpCXBKOThstKbr
4G1/sv6ayEvvC49Y2SGodqryyKhJl1Xr8DWjCKIGIcI/pj6HEgYlEoxApJI+wnsh
K2pKPk/IqzNmNC1q4drC4xRyXFFaMHABuT+JOwUXkol9JEd92kVPpyhDECDVQn+N
RbGVrfhVT1voqcQTIIpjQ1exojGYDK0anpgTGjps2llfh+PJCrZpZ99LmE/xEd2A
e3q+7LRKsjMF2q5wu2JDPD2K9icLBJQRsxVyEEeh5bYlMI7JYP/gFcQej81yQF/B
3JNIrfOpOQBsDzklcReTi0gqOMOlbXbwL0j2R0/CFIZ6lENUlgfjuf4gQLUJHxM1
9nUntwbbPgacQPykibly6EGby8chFPSQvABB+Nld7Tcl5vnIdjLPQP9Ibxhxvaxv
15GZ+qA8Zcv2GIb2Illz8OW9t720++T2sSVCf/LjWSeOclprO0oeiuIuLOUNI8Gi
DYXiZxPAJWVOTDx2JyJ08ER26DKAOuyR6I4YRjBHJr2cRyo2JUxWqbpknUrTINJA
f36pRoeezR39g/PwtZ/ZoEus51ofyy6dDi31GyZJMymGQdtn1UslLtjarxZjj8Rn
x3APGXarxNbCXF39zI2dEKHOs0itx5wDNQ7FUx/MihL2iCgQk06dOHqnV9DsF21h
qzgz5S7/am4TOdItNp2sekFgFlD4LPenO4rX4v7Ag757Bttl24/dV81C5XK/5hHE
36p3xl1EDE4QZ9qAW8BruW2vDJg3ritfyAjcTy8g6r/u8tBRDAGDihdPIhOLKCij
tFyY6t9itmNMB0fzVSBaZ3JvGHkkFos7Mi7yCse2Qwf/1syTJ3jl9PZVNkMQ+fwV
rDk6SEky8PrpnjvtKLfWsgZgd1PvDSpO00WQxCyAHHD5xsZRvMOWZP4Zu4Z9JdLL
4mXfcUwA+VucDL8ssCEp71EjsOVISnQI+4JSoz1Pazn4oJw0taI6zbp3t2+7oPS5
ZdJ152Ga3NoqLsBnixukO7efL3fQ2FdP5oahAjEdBGeabB1oUbtfEoegc6DkYKHp
k4VE9dYFOq0AaZ30mWBSZuWFR8ZsjTczDf/wejmUgVGavoB+lHsj4prRAL9KSWy0
Jtb7Yuh1qF/8o/6aLTM03hD8IJO8yaAvyKV0a44TvzXU/qUAZEF4n2Bnzk/INGYr
S1KSoUa9rPOsSyvmghpEFIRvJhAguscequE0PJAw5K6aNQ1mZNpWtRLWq8GwK5fN
6todWdevYhs/utItM/kPisSaNZgT+zUIDTINtqoDY5pPTcpj/BVaLDD/1+xnaLHO
O/q6A8hFC/tq/Il7X0I86WdRn9i3ZxXO76UlhWNPp5oBaADhq+HMxhVKZtxXLHYZ
8UAsHDzk0+kdCACie6/y/96CtvrB/V9UlqdFbbIgesuXlrlb+soDLBTaAhhEwzH/
S2vHqRmbevLSxkuBqlcBuImhBfzKpf6QW//D5agseKjv6Z6Um9AcblfEnWOewVZJ
6xrmLrCyE/YtaGysSMHeYtKE1BMI+Y7EdU1g8Koza5kTov5eNNQ5Mjlxe8C+bESg
2tSVJb7hrySYTZQBtehNHh0JxOjZUAXCgM5xtanOwDPZGU/l+NucUDJ/f/ZNSi5K
3PJoqL+z4y+s+8hJH4eSYHSsiRXeZ3mHYOEtkOrKbcCps/ECbXr0xmP/v9Ir5pmS
XtBct/oREERG2kGnA/3e0vdFVPxFXOC1Lsr9ZMMwOoThGVPfPqP1l1udxYzWUnvF
rlmONOLiLX4nFT6jmtLGENPs7VDqLFiSQQALIYCyd+M8XLrNiCC6Kit5sKByeSri
mFzrMh3X740KLFovHTkhGc2rhX4uzOnLsKwth/l5W63Ro4+IpvC1yJxH3n532M+c
3Q68nsdetLcOy2RtYbbZlwoeOtx7RY0uaxgNBc65M2QqtmmZiau4Dyl3jh0WYw72
4AGjawAok2zv55suzkoODuI8OHLBUktPwPWcNfteJMTFi4qHyXiof+pq1ggcc9mn
/LrjWAD4Bbu9veBOM0e2ydQVK9AZVKsjRgTAClt2t+Jdofu4Dq+6Wc44QbueNWrV
iHfoHUP6Z8Q8SOPGABOdhISNsbuvWg1+JJ/RSQAKYyJ/qFGORlWY+Y0Kochw65Rs
mUhsa5Dd4YMxkTjFAz/MDr2iIKLGlJBlRS7o3D3Qm9ZXqr2xYCGB2dwWvtyftqqc
fjsyZ9FhQH+Q1CUB0GDA8Nwro8p5z/OS6IX9/edzUGF+8ZS+hUYUMQO4/ZPoY1DY
CyFEc2zzcph6yrwAV5SwiQxrgnQRafiY9UQYjAv5KxAuWfejeYtBP6GfL5EiQXhZ
vrt8Lj9N8giJqWONdNvzLZdiU6RHFpqVrPaS4HydrZB+PlKVr3j/t0dazL4Iysjq
K5VxPYb44W6yveRHZpWOEX/iMHJfLyVXkg72vA6J71uKBBVKlXd7WKwKWxniuK1D
6oUEPhdS2cFx3SMcF/pRnButvXgRUJFSLKALZRKWCAmKlgKFyBs2XzHWz4r59KUn
8qJi1xZfk8fcnMitv1pVKQkub5efYmLqGceEcNy/El+3QqCJeKCTHpshsAhPAcih
K02WLrdq+2lPgZVDbY6R1RUUAROVrWg8WWIpo4QUGDci2Z4Vqu2hDVPet7n7TGn6
IRi4ojvFEH0laDpO6eBkcqnasTnHG6PE8kbZFMJgVGAhiKULXNKsnQIsHXZB+vZi
Ms21vow2LYCIaDwFnFZn8MUaQoYXsmaCQ1vxVMNcwTpi8UXSNCub7NCj+r9MJZa9
EQ/0QitQSBD9itulmmL+vTbI3nM85XtIwVinhH4K+2x/3jHOnvjM9i7IU34nWVPm
5yCuHhgepYsE96h90tQLx6EHz7rCO7PcIAnZqBCVZoyBBJR7lpZNd0h4JplWb1Lt
jsRFH3fxS/M7u7cJUGNbxsDb4rkZKNyRHYqtqBtvoT/s724HQoCXsI93hZFrImqV
mIsG9uns2khih0LuaFs5Gps0NVz91hg8xLwGY0cS53wWHnZuOw7xwgQ68XAhDH6f
4m2G7p+F9W00TVUj6U4qdu0mxxpmwF4HmL2831EBdAXspR3jkn7zDGFnGap5li9X
VUfT6Q+w6Gt1NFzCVeeeNx/Fg52jYIu3P3lras14PbQicb0iaqwXVEDnJXAET1GN
l2wkYeDvHFJaPMA9+S9CAKOndPP2BabJPw2gWyHRiv+XF4x/fhfeclfU+dgXNR7o
hmdLN+wsLsLBDpBINhTog2pXWMalU+wifIrvN9zAadPOfyLusN74GnPMKVKfM4yC
uNFjeDsxZb3WJIccgwRNU0awHIK5EGCGce0QfBni3WvKUJfpxEcUeuio41zGhgVY
+48kiATkgGfZHTXO3oPM1aMuqWHCJV+dmlmstGpVjDHpBXBApm97RTip4zzPVwXV
vB4lfw0HgHy3I0KpsxMaq0s3b2UNMdB+kuZzetwVOk5QrMA7512XjWQPkLF1U5Nn
jt+66znrBzRTx/4eEu8Q5SPY2yAz4shWbGNQgRIhFTje5xOAICXcfNC2vFbSTt5B
noiAiVm35avjDKC6y23fmM89lmdM2NGIVrvoCt15ECiF4XgmPjo4U3IAGwPkYwJa
YOSOdNei7VzIli1c33ZUMgU2pTCLRNdqiy0Q+bd7eK0CxbjLQnBV9f6oYbnpDTgl
Vbl8f+eDq72oVyESovtS14cwgma9LaG2TFv0wxu1HmzHOghqVvathqJssmq8lybs
Mc/4JkH6rGraGQk9wBIL3sNfvi+YGieQVaociFF4Zi2SVAcyomvfNA7G23E19IWI
H9+VY6ko/ZU5UmlBhc056C85vtWo3gk1T0tM8cEmZnHh9bBIC+jp6wADvF+dEyUl
BSXkhVSR8FOLMBb7TdOuMsTMpU5bGIvukKpDlsAZfdUFgqnC9yzOOrZwtd3knBk5
JdSIfF4i21mk4zYsgYRDdsadKxcgFozS9N+Xuc3nhoI0rR2SO0pufFfO5HTa+cJB
ky2v3X9p9n6es+T+h2t9B97WlHuoc74MfvDXyzSbckLJXF6AOGGqnR0FjfrrVBGb
Ng87ht8mcTmVUAfzGFwuXlksFnI7K7aNH4Jb2qR2wHmwkSR7tjg8Qi3rtD5fKb+f
CBDLXCO7946LK7FebaoyMX4JW671+93mstBW9xcl44VmBToSqu8BEMPohd+FyS+/
Jpo8hkW7r0fMtYszNpnxVoUK1qWGXHU+b+edgOTk0e3+O5zYznqnyNpQShSl2ktl
bLpkshyaO6t7+/OxJyQmyqF1pQugJUCGndmL7oH9q7QiKxq2MLQsspC3+qSssSXC
LDd6tygxmPtNqNOkTN8Oqr8NovZdOVEHJVHRmOuftuby16QExLLDs40Ct7a/fzl8
JJWLSjWw07N1WVrRR5JklLMTu31cDpPtwruuGB69g99mcK9bfypVsFokVpHuDRGs
d14zD6D5ciGdENMtKwkTKxegSdN4LyTdu2z4A57OdOQATowA+uUKBfzpbbBspj2a
m5CSXvDpZOHmCwhmnyAldQq4Wy8L6ohRBHt3ajTgPA3KbZ0rhiEzPwDM2UvpLM+A
hE/oTs8KW1n5cPmXsX75WGGyj6zfmP5aNOBX8h5Yf6SPXDAzrggNLbIIMsQFvFKe
KCDFg90sAYIwMXR9FQ19+iecMb/mAQawPncx3/7GmdMc6pHkAbsxlk4RyqeD9iny
5AcKomFv9Ni4QqrfVnIIa99PEPV6sLwqoUJ4YMs+CKX8xmE9+T7Eltehl8G/M7Zc
wexmTr88+0H12DNl9oFkZTAjTe7djRjy7gazKR8T/g2Zx7i4cPR5or0hsq55fQM9
K2LWSZQavuSkPnUqLl6iVoSVz4Mayj7QSeeQlif3dY1Q1gIAhq4Nc2jdl9BEnKnh
1lnh96V3/V0/d9D0GOl+kSVRphOoTPocSrDyIge8BkcsP9EB9cDewQDwKeN5lSym
qr980eWeEW2bmzrZWMJ9d7f7qR5dsqbrS1GhHl4RPxZtVRyMRn1hP0aiQxKmvQHt
z3CvEPeIkerGgh0BKAyk+hBb4Yx74DsfPvRnV7pIqaVl1Lh5eFIGUl47i5+yGZ/c
9fMd9i+K86Spt1MX1TWypkjqAB0OdYwzSaRFqD9kOnsjh4sPWkO6sRoSyIaZeeHG
sUXnx1Dr4XWcE3E+au0c/s+cdmq0Gwm6ieravj1heLBY6AXum1k7rn/DJ00Lq3K7
9QtiXYNI7SHs+fsSU9MoUuT9okRrD6X6gJywPYFYzV+uz9p74NZtqyErlZ4UxDft
xNuJh8JwxRZMUwIzxAH9qkY426wYRL68LmHqUZXuLUDg/OCm/XnBhkzSiY0CjwCS
yE7uEZiyIuXZ3E2a3KjugeSe6gZDCTYJ0c1CmNzgSzVff3IcRxuHLQccPdGHp2eW
ShQ+IIKFqtDUtP0+rQ/zCAdMXHJ3j59b5nHRNawr19fSxVm17Qc4SpaFszewbG+u
bg9kIP2rZgdNMB3ldICRdRdye/oabXW3Z5eaIeAfRlTmfESlrRroUNXBomj+coZO
2ZJJ6O7+UevrnNcsNDOZs2/98b3zORQ62yzSxHEU5HwoFlMSEl2WjPEspZH4op2T
t9mRptYjV3c3mhSyahIlD6quSVSbEKyMMGLLH5l5Ecx5im+Y7nSLvVAo8uAmvcST
Wb/huXW2ag2sM5hEnfa8Ox4BIQ/UKNMrOfbkSjv6o8lT4zd32yOtLDxSEiFuw6qk
uMibm8QlcjyNYrzMroTMRKzMAGiHXhsPe7QmG6h5O1eRJEqhH7HFar7hZkxzbhgo
Prpgk8Fww/XOSyDb4+mGFtFZYK6kj/oOKxcKhdZb5FhnGTXks+eT96wemb634Dkq
TVkvrwypMpuy1XD85E0Hl9YTs9EQ4Uy08vPoyX7if9oNm5rtqRw+kI9Rh+kL0oVP
Y65KKQW8wfix+kgUA6HkAlCd3cmxL1yoaoVTh3lMea0m2TuJEPFpakgmgrEtmYtf
xtd18pdS3TMTOWNday+eAPn1iTgvfeV2s/Z7uJxIYo/YejaWucvXccfGc0feAqPQ
8iPG6FJV4mFwWtc6Toh2Cm1uwiHnSA5RAgblbREJi3pJyGXOGkBisaXj90cVpAFB
skeLKGdUUPEj8MAAd7QvFW6VbTIGWSV2+O44ueLonEnazpNDDelEnA85x5x7R4ij
mspvumOm35B2ec72iLZ2efPbrAN4qkQgo50KsfoHp7wBQWCESjEH+y5BSy98Ko3t
tJK4Y5XlvKFCKzedwhiCEJh1FF0thI1MdyxM+VuReXCyhHUYxN7kZILgnu1T5XQK
vni30Y9Xm2iEF+UuWt3zDxsaXUOmngBMNL2mH5CtZfdesHuq8CRNhvQgnnIPg5Y6
35S6Awb9N5Q4/FWzNWIyBJ2JjCcfNghya3bv8E7zS9rIqqlk/bo2yikoeJ3TXdDv
v0WRmNozZsCwrR7wsd46jLlhq/LfabWltSOTWBAb/yPOiTybUtTyt9xroj5kn4vr
3nGtvHon3z5T0Z9EUd3Y6vW4BSqnH/K/fKwrCIJfa+l11f2m03DFr4+9uP6eTGKM
jPRY3jGyI3aKphxa1uX4lz+zGAsTs4TcrdhP5cX1R8++Tsj0BiglmGN67q3TV6GD
+q7UAkD1R/sQUCIlzaEPCF1D/pWC9hRfWruFIGS16gZG+MCsyLenjK/48MKPPKvU
FXu6WtYXLuY2p/fTFcLavwSdiShSlNiAcsSZaM6VMugJLUOjrdPQacXwxPfsU5rV
pdbk2cDT4HBp+nr5cKd4VbAjA725ge+YZs8C994gNU/y9wuoY1LxCoC3vBSzcHST
hqHaAydav1+baHYXneYQD5NM74wTOPkqm/NdOrW0QpUTWEatqgPIh3x4e4BGNcvs
6/vomBTaIfXDme0JqyrMZQJTHvdQFMm9USw0yueFWtxS1YyplVnRmWoiHx4Ggr9j
kOkCb1ZjWPZWbPkBqJCha/nZ+pj2t4sVg5kkVBA1gjk7n2ml4pBrjOHLMUZrcq3A
NgOtYK2exE87so65v4OcidurYmZU1fi37tesbvwmjsf+RDc/U220k39aZcJ/KUv8
HnrSkTXGdsTpIPrhgT4TaxuRhd5AwSLg6Dd7jjma6NMB68sxJyUFy8jpUGtWns07
oJFhpfkAgJ3bMTcCDgpXTqflGk6FnIgPWnnxKyvxACcjTcOkWTjehFQMHqjTsty3
9NCGK2beUDz99tXKr/WZitHvVhiiYQSyW8dfDsWZw27L4nTs5kthgH0JC1Zs2McU
8Cdsh3LJNh/q5dapICHaao+uzoDtIzGXkeQwSx2atK1Smg2+22e6DMEuraaXBzCh
aFaQv4zmBpQTwr+vwKeCE1Z8wS3SwJRaqO7tBxGzJGBMV8oPq1T56QvoPT2yhRLH
StlW/X7wIjEGMh56ZXnnCCKfqkRAbXa9Zy90yxdQVB9f0udCiuw0MvxY27Regbuo
9wDQXKfecemvDD/c1TCAD8JcdXQIchNFYxSwD3HsowbELw3qxcNlp5kw6IQCgygY
iMSgGxMOfkv05uB2VfMTzNUifk4JxSIVZYWycZVubDKOdgbINkFAijT9C7iZOnh/
kWdl/wNkBU5hQYI9znynUWpAPTSSUgL1aOzwuAPDUFJzkw7oFh4/uz8iv8U48WJm
c8Mqef45SmHegvNGcSeRYry4SufFjDIJqcLRRxVfwTxIfU8QS4drlh8Gf+9A3KlY
/DxbVIZTqiLlaKDZZnLNhxZt2Jen6x4z5D8YjKmD5Y1bsrqKt9xPD+eVm8sVC3dx
XHtybARxt1iVALCO8/SvGyRD6kc4aGNKsMENLGxqtVC6+WVLGhs6JL8I+8try/fY
S0zYUvf2CqNN6Z/Ho59x0yZscewk4FeCt+N+52vcxPGNr6dOKiNqSPLXrS3ebAAm
gda/ssbRsMqYhB1/ZNWX/8t5mslzbZEZgVy8S0nkwT+REI2E+yKG14mnQZE2K81b
Fck8MrMUgA5UUbVSxcqr0XwunkKoap9tA596BW+xMC0z8OtR/b7RwgPF0HQpRdEG
SEn+c897otCuDzOT8oy/7A3R2cswsw3gmOOJEL7S6DptT5f6V1BOA1xcRMl3/kYV
3sX5TGlljz+Y7EkfNq+UotLUqY33CuNNjE5ZzdEDloxbuEFlJWRsDo7uD8e4UY3d
aOB1fA7XRSKsGRiOWYSfGjFIILfGhUWgtGgPYeoLyfcoIUrFD9eakbWV8lG5cniq
tLSlQufTlbF4Xiv1vGDpRxIrkHR1W+toq1UhyGLa0OmuJNjL5OWkA9XeGeEZPRGm
C4pljXeOVOT8wAFsaDuN85aTQzGY8+WE2dXYCAnEF7N9NgBDsBLIUePXURRunAAm
P0Zzux3KeO05zJiPg/B/B583lbZUkj6M5fYmDMy3rQnhOuJpae/T+SlWGypFUZ8H
gT2faOLy6Lvqc5gAD56k5zjaVhra1S9K8/K91E6Gpzyaq1iGnSlpaqStrIl3jQsh
UXTHVC0HS/Z+BVxTVuRHcBjVvboHx5b3GWbpsj7sappPM1cBXWpPjinLzNKTtwme
cLzdTKKxy/CTZhrc3em2LBp+GUqtq0jxnH8AmLnSkXwizNIHH7ClDhQktzIxeFyI
47yw02npM9yBL6BPa8t9Pl0lhMZgycw5uQHeDxKhqqZtwgAt40ygXrgoRxwfDHmk
WCMlG+s0TCN1UpgN5CdJU6wZmQ5NlOffAktACQULH/d8J4LCsBH0fSBjRPpolWoJ
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNYqPUtq4TyjZUJD2vIuF91OD4MkGJeYB8LcURWq2RsCKGG9wJS5oLKNcQNQ3166
Wt39EBY+hptJ8CP4TBZNl6JqaxIqvKcFikurjdOKCHdlNF+OqJKSpwuvu0DthVao
JbvsA5yvuoNPnC2iDFUU0PlIiY4nqQ2Zb1liMS3ezH2v7jtvjDOSXCA/Xk7r3CuE
qfxJVpplCLZogJqSEt2SR58ax+VU8DdWWz8dTpX7VBzUe1sSuou/PNofwcZbxk2z
45oWwcb0fvjdZB/FV89xoODhVd38uMBK9oDl6q3LLpqhFr9in+9VI/PVk64mHAbT
j5rD5jc5UCXkzm3cv3QtT39+4hIJtN7hiUpMTPaP3w4fSGxi7Vy67uffHztluoFk
982Di/EUHBS9PX4Sm4CSBC8BDzpeSzZhMObyCIvuXI6CnxE2q0Dcz71IwwkT7zO2
7Yk6OjnKYiPuLrVCWIRAyhae8XnTr7o8/Gf3cxPgCMShJa02rtn1KAbTIfNrlwI6
/Gwb0sRBUXEFcsYylxp71B2R6RxwXo/U0/X12SqPwqm2Lu28wXeI50cS85WBwn1U
otnE84PMIkxYPFX1W/lAPp/tKhiX5DWyBnHDMbOict0ZNZ0Q3F+01iNayuAjO2vN
LZK3CGTQ3Iek7iRCK4wSQRONoWMBKm1ZhZMWASACZ+XxQ7VetCVULEp/qLpkwGDR
CJz6L66kyDKoxzhztrfd+rINALEM+AFP1lShxhpfyuLy/t48c7a9CYoDmz984Nlx
JM0V1iPlT5pL0ck9F6Ls6d7w+KvssMgF/oJdIXgSVPevkHYpHGPcAa1vWjTJYF+1
kjJ7WtGtpbIkSRl3iv5/Db16SBRH3NE/HitYQ7TLLivoXloTLj0Yms3o3iW2kAoA
T2MQTpIO/1QfF5JZYiliFJJsO799ev9Id/G7iXD9eoFHKnkh57OXX6da7MB6yT/f
VGqMpXQ30YMdobUy36FZycwLFpYpD7LMJebODnoILAmvtF24l36Am0KD4KRdXVbA
xiyYeKe2nHvOnJ3DKBekpWIryNg2ftfreY0WgPLTwt/FrdUq3e+imhvBthVudtNA
QhP0S2CPnUwclx7S+v8cQChYGxmYnw3UFQj/NF6yUjGL6YyN5lUX0lMolNlKAwK9
mpFQCmxaGdsmnifs5P3jSfYOFZM2/pETbnGP2xT+utu5Z0Z/D8BEAhnJkolI4KAN
GaOK+VL4zShWB1XIo8y4YidJa6RYT0lqdI8LGhBrnu4j7VdunoOra8xQ+e5ahKLr
b5mb00WZYFGP/y5XNcvHVslEycIJyGysd3N8ISUEfSyW03tE28JNi18TkqrDFI7k
nb0ox4+kI/lxwv9aJqt70UI8XQoEX0thlrPDpvAxj18Uui7okv64fwc+LpsoWlNk
FKkqch4Rptxn1CEg2cr0aCtsEO/ekvtPZWCPzqPRWLxnSEoZzA2O54DzZO76MSrP
BqOajk2BLBSw+ZRubrcDjAnaB8lFKncGALGCMekSFuYwlSPMgTNsIKrLHcl5q6pu
sABYiLSVgeIMMMsWprxaqZVSgreTYZvFfuC03CR75P/F9rUlOj0bDy/NAwKgyzXL
MuOXZAD9SrmeyAPm1rqX9JpfopeJwWh3xIyT48JSIvXgaO9MKtBtPSGkBZMzqXJy
ENjiOxZGYvTOei0Je1omu8pg2YyVK0vxL5OVeFkdQ/cBFkv5rdP96j/PodYzTSI7
UgZqz/NeVk0Ei4e1+mshHlhQ2/ZCRfNFmd16roLwVGPoiG8mqZKBhQpoaCg+KfCX
jxlUam/cY/soEEbfYUqo5WXUHU4/R5L1ldY62UYhG6SF8zJYzqqmE3CzXFqYInxZ
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vRJWKEVyu0CTUz4nr8Ca79vVv55EejAUBZGo96bCP0JcctL/pm51oiYFISMbp7oQ
TzEOppv0xxWFZ0MT6C44Nvoy1h9BYEZ7R9Kxk09Qkyr4EHDjSrW/nb4Pa5XrtWeU
h1eR1C1IYIWVRsatiBnp7kQfYZqgKAfEQHoRJkW02s1viwKbdDG13YeGWCsdRugd
y9SEGbP+idzOrLEHO3/ERLS/p70DyV1Oe520OSp+IpmnXjTf1w74a9FhSGWFgONe
IpgWq1dzH9Pb8aayTPqQbXzYRfWFQbFMm4hQvvOW6RlnnaPbaFqw2lpDbGMKOioI
6xDUoeF4vBKsIFcQo6VYBnykEY9BICsWvVs4gGYPrm29DbObsjumciYLXF/pRI29
tc67OIb62PX6hcvY03GrDPEln9eUhsYLFOX8xyVIRzAT6c+ga2DXZwAai4YStGs1
GEUUhkT0PKZGgU6GROSC88i3QleBkn8vboG1dOD8lMsTPDVn4+g1ZAE6wHrcZy01
5TE1a8FpzFi6CU9wRnHtoAimYk0Zxe9lc6BtbWZWROXE0UQ2/KjIWTnnRFX2jB1f
CqEyOtjJZym15nYzBJi73G1hOpqJ2IMJQTfejG9MXz8QkI3mgXfckZLyh5tSqswK
JmWIzPP6FV7rKq+Aiskg9IRVUYJx4EQ+/p0omlxATtQ3Ul6sJrLEXfE+4V+2MpuO
2883sBag6g6nVNobXycThlwMS3rzZ3fYE386IFsezocyPnWas5FmEypDFi/Dh3oJ
Fx4fdNyccyH/JCdAvyDbZHJr6zO1UBlDMMBv1JuyjDt/7xmgfQN88gTtdocWGEba
T+DtiNcDFpThKcPoGrx+VQc/4zW92wX6bsv7Er3zU/BlRD5e6RpA+Nma1dXwKPCF
3LrAkojwsp4kvOEzNEBkmPpQ9BVU4dH157++on4fMu1BzzPphchVNKDHC4f82iZu
kXv3kFGydDd19eBbAkE4PeLjdbIEEGC07jGGl4jfu9rtDbewdkjuAnGT6OjBS+Cc
yK0lJfs3FPjvKmtm64hOXfY9PSX2Wz+YTxq+a4Wi19DJGQIfena+WjNKYt3QnaXE
ASB4yuWKBToeJ3/dx+gzpNhWRVPiCx9gJY4yabnsuEo3fPRncZGabC1zs4plcLtk
YfxVnTitsvE3ZhVM9vxaplNMKCEPsyhtBEqbn4X5TIOSqoqVo0unVuhovyWa+PKz
QVn2jTJFnshJ4wGqunQtXEr6FfUYzGtPduZ07js37nKNvqfFK6LdreWI8MtIunBk
x/sPq7U/TfO7iMvMx0AxIymreVanqC5J0ZddRejkzzcRimZt8JvgZEDRmNJnAqKq
qLVznLY4b4bcF0/qQMXst5p/kw8TwKIyVsGOPPypuCqicgI6CIJPEs82GlirAt1x
p+NvhNPwMHmKS6svEvWeoJ1lHbiEPxJoloc93wn+WU180m9Tx7sBzUtYHGnhOxIR
oWdi/E4KJL4j3AImupvULvWjeSmNjiVq1LqSYQ3LmbPB8o1VpY/17LJga0xOW83O
s32j2C899Xgd5Yc/LXdiOLm+ERHXTGoMqu1ZKtqlmJYEdnWvPBv02r8/dMdUS2M5
UMWyOyjxJWzVB0s3YQlAIJ09CVfOvrhyhBEJaVbTFdKL8SX6DSz19w649s9L2oO4
XHuqY4lHr6AZF4hvmqdvHA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LUh//Pd2YPN0R6bG5a9KqX+rWVrFOsEQYeeZegJO2PUCbWykJUorkoYa0Yr77vVC
ghuRd1h2JUh6sbSDoO/oh9TCYzQHB8HMb4LOT+8cPA0L9L3a4W4mM6uzZb1guXHA
2rbBY9CrDukhYSMXAmziA+g59hhj7347M2ItieniblNqwL6NnZmUa0kaKbRHXmcB
4PCIHzBi7PTcxsesiZ62C/71CYgoO2ceWOfmK1B7Y50HcwhDhOP42Jfxo/kjClHn
TW7Ff7kwX0ePeFo6OYez7vGh8L2CZuTEI+RlVOwCunDRMMdohXklajtGZQ9azzRU
RbmOys3DGHGKoUhpIUJq+ImWSgnrkVYhQmZl33ApptuGtxgX0SSCTqWxyHGKU81X
CseUKu3JYdlIM3wDQgGReUdooyCwSZz3ga70hsOEvpCgZ8eUw3Fjy4X4icsr7SSj
ORRClbjfjMDHfvA3VLzbWXvMvoJPv5JRoX2penP7vOQT7CI4BINJkQQP3kpeyM3F
utAXp4DLCe+wnv5aT8ym5oLdd55gD8jq/G1xH2CNIZiJUKlp+xiLmSKZv6ehvlrk
Bj8Ofs8vPjqm+sdLsuIa1ql72GDJc6d5UvHg/oa7DeVBWsVLhMjLsOZ1x5JMTCuH
JahDsEqYFyslJFf3kNWtP09Jikn8JgMgAGp67AChJpz3KeJJ0MqNj79elAqEtKms
qwiEmBNsA6lxwNiBAbRo95tSemLYv4ahlybhQGVtYQAti2UX3DlSd63HIg1xppnB
vrojPWJXonp8yZvXjex4EVJdT+b26J3qSaZKJ9R7moEA8dvNa+3Ma9sEWECWm8/M
QRDs/Hld0ZN1tpLgDz/PBLZqM493UNgUV8QHBAbulgzqKobHGxxXma4ddl7UISnz
8xBlRSQYCBabFSiPi3WkeaS1BqmfWi3icK8Y5dzSopz3wrpoBgnnr/JagHdIvsMS
YBgGvpvsx03TqZGLUtMCzxeRrLtO4gGuzbr1zdfkMgh3wN6zIcfF0tJ9c3cmw28S
pBZ4NQRl8HmNzS+0DlovGn/fLSB4gse13LH2SVJAyyoMH8zUU8d88+LOUHPeaMKM
bOFSliMdIeKBV+q+MsJmegXxSztNzNYNeLoD7lxreD2P42uZdHJpSh9xIDwI/BeY
4EqXwnB9JAhX+leg0Fig5RUqQbVk3hrKvcy4VNwB5h71z+yHRt/X4njJEjuQPKLz
sCOwB9e3bVCBR4fi/cZuXDafP2njE6+2hRnMCk0VpezMYB/REr+JDEncWwSU4Qzl
WAE1gyVj703bNrw+KIQLcdW3IMZjtQtIZTBYfBIQUAxyBxir3prhyVOHh3I0LbXr
tYmbbjPRCI0ZX/HDUKaR6Q==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yWJEESlOjQpSA+C1Qn9jLY4irJTFEHZZEtAiGx3UkmPPKk40EQYBmZalP7huJ2Ga
NBsz/9nPYsjDShFU4fZiMbVrNbIZ0/oYKlUGlxkvJbFMLMq9G7Qa5XuT0bB4ul/x
lHL8vzTH2FGBSFaeWtrRZpEVLpnupvWZQpKAP/Z7vs0Ev38uxCNZz6iUpdOkhzyB
FcC4kBjI1Z0jrJzeGKMEI+YzKB9K3chq/hM+OdWMNLfMqkI9VNNVUJTPtOmvMkOn
aaWxUFJT6jvJrEFY0jUHoE64ZtFqQ+RWotn1Kwc9mCfUunP/2PEO3B1rGzuoy0ZK
Izbl8YpGLwnP6/PzpBv/ljgPIge+C+pIvGIw5uOLsuFg0mTXZ/mozowe5npFJsOu
8Zgu5SsVaT3jHwzSe/cAR+qPlkVUif2JF1+GaOP2+F1lvxWfqyFp4rmSl6Yl/Y0l
ZxCtlZWlD0Ff6avKVWbUQsgI6oTnNIBTlQP870QbvH2r9OljQ0WrsTQSPEXtAVUC
GH2IWQKKTUxPQ7pIa7nO2G5uJX9ffoKkkBcE81MxD2WJ/0mN1bYayW9Pu+qwkFVc
Cr7nPUYNEY7K60oSeFOpIeWAXmQPOIhqCMOKTDCjFXt9AXKxu0Q3vR6uzWLL3BN2
lCsdsif7WoOZPOFTWEOZMSHMPcB74mrgo6uGHrUIfqvT3OPsstAyjuejGCtQ5Yg3
hchKVLwrTlxGCBEPyJ3ddMG7ZjVhYNI2iOyN2HMWVbndu9r7TLOz0N3cDTy9KIVB
oFqn33IdX+Ul6pe5Pj4uOjH04K5NK6kWMNezko9AY/RVoU8o8WJVczNcUrf6bVu4
rAEG6rpqXcj+Y3qAJd6qTSaBOikiYhOuJlU2/V7cCEdWUll60Su3nmXls+lCi03U
G1X59Vld5Hm/TF2wkpthjklY5sJ2/2oPKYMR2jZXbYrw6cglJUloPrr/J48luTyY
wAU0AmJzl1jFShEK06OqrU8tq8vGSKjg2kZfIX+5KaKrnFZGitaq7FIvJVmoGQyu
GzhFdVj2toFWGuPBeu8S8wz7I6nyb8Y6LnyOqEtAF00HAj1I4aVxyKGRVxa/O7Qq
4sMocpgNL08+/Sxi96/HjuLqoyD1EXywGtCn2unKBXg2zVOnVi2JG+4n++SGo7xy
AaobDkvlZ913M/L9CX/NOJGpVq/B+zJ8vWVSS/BzY//jAzh/O6KnbJl/gAVYA4r3
LqG3msiZleb6eC1o4WtaOQ21R9xQFur4KDjtb4hYYS2RYdy0t8fiTj7Z9Uabqji1
2lbiGatgfwoqAeU6aBP1hmSOmF2ZMw5dAvrg4nLnKhkKccANiD1nHiOghRtr5pIq
R5KlCQecBbOVmIeyVq0rbW1hpCjiMPDDjxybu3QtkPluVxNQ2k3ehlyJ1AjAxyuo
eOHv7G8TmcTxAFTFHtoyWnvykfrai7a8bPGi7wSA5sCR5IAfz6R+iKE1wbIjEoZh
Qhw1nDWpM9FLECqBcPw1wFzDbIdLy5DimmnjXz2pn5ZF8WLpnYufyqw077OPM4fy
VME5X0a1QulG1Yy5t2uS1niFJzRAXd5cR1zuP7cJqZlqTAG9HudPIGuM2syFtUxy
tjZ2svZvhlnL7qO7L9sDDQBfh/N1QJP8KlCqMHkBrGGhAfvD8xK/DY4NasDKql3I
RTsE3FgC0TycQV1B70B0j8a/iuUXsYx2leLcs8Nu3/y7+wgfMgA9W8BIrFQM14XB
Bvfaj0+oLLq2gQ9qcks/VkAPBG7zDh0cvW0CrpT6wBeD+wTO10uV6OrEhXVq5sLx
ZkS1dg+AVqogYEvQjLtzv9qIBIFaPXPvHHOtCaS4jSelEra5zuFS34u1/OokCuwI
CpzGiqJEd1lBYwXCHDMCQQmwSbF6aPxNS5ccYoF7Eu0mWtxrbapfSTdo2QREMXFl
zyZSLkIXSQFhF45NUO4QoMecUllA86OqUUWyWM2MUSWZ/VPzPwgPBNk6tVjPTzGg
9OkJWBMbcVL9lefB6Td+1etwm1SInbsjqXKLXzK4z4LSQjEAE/SLoyJ0WMJURLYJ
tIwIkw/wt1tSB4l8G50PJYqHNsaMEtkkf79M03cCPY4Zmoywjj9YVH59FgnRsneL
RRhVpHw2feCPz5SyrYzdMXzLFJosMmDUTdaIbXi7PHD0pmRFJxH7GjFJ45Ktbeyc
BkqpD+aCkt2YyIE010LaRfLl4cYPmkEsGjSz8HK+WAO2WO2F5VyIJyA+L6VyQ+eB
AIvmCgDwv4cbHOznb3HMNzNc2fxamsr4SpS/OXjDCQKpgzWQA2v0fcVQYbIB8vh5
Aa1t/hNbKDd8hBCQuDMON13xpLv81qekzd3UnsIhbRTDylcYqHUVW5yjyva+ZBP9
YmyGyLqDaClK2lR1nMzbnhUumXdPpzMnVySHGpFuncyZ/dJw6yz/iN45UGUo/mj4
WmTQeRFux7ie95DHkQRfSyxNLjMXx9pPSfp+sf0aYjcOs55oo2QXif2a34tSQKtK
FZxqZ6OKo5JF0+P93TutjLSm5uC1G3IwiJ7H7ywZmN89pPV/q1YuMEyZ+6Y8uAtZ
WrAboI2P6EakKQo0VzN3tUdijyD+y88LBfHcTYAoUp35RR44dMHKTprg4PtsB3B9
3MP5SkB3MNcb2o/JHar6iIUPeIjcbTYDOpej5hh5XeJfnfJ4qOgg61Y9cos9yX0m
RwY5L1ScGKRgatbLEhAUg9lcsuY48DzexhoisT4YgtD8zsYaBJhcLf6SagwV9u6M
3GuyIhs7R+wVI0OQdStSCrpeJWyz5XPQLLvBXYK5KkJizHKVeER8KWc4VShoVarW
zmjiHT97NFoS/evLicn/0CvAS11MhtFAW9w1abkBPk8/D0gm9lHnXV5ZSUP9BXnC
8KvHy/JjUL4NpwuaQm3Z3uqNcdiiay1xlmteCWgQJFgGKvdZLF188FE7/4vmG1QI
NB3bqxGTUW6OsozX+jliaAn5RCK88wwu2OP+610FlLIimPap1PL5rgzQrWwTkZ++
ivURuX0uj2OrjVNQW6fm0KcpfNkuRk5075zkh3qa/WLRGNMcQCMP90kh43PxA0iz
CVt/DfnGnewMM0haDK1VFzKlLAdXG37zQAG0AdzCqEhEgFZ8l643jz7TX8FJ2IKG
T/WQdJWGKEOxz4yE9dXVQ3iRiEXixbQ2A5UTwuoUima4nq6DlDt5FEkfyXt2Pzt+
poh99xuNOSy1DHpt1aHPcH+sALJC7jjNfnJTLRKhharRpUfdQLbfArMV3PPU6JpW
qcT2rQe31vb0YeFkPl2c2bKoORK9IaGnyzN6XtduwiV7Vjblye4CiNb+6KkprVD5
f/BOooF3Lcv/I5g+r0KLRvn50inSr+kPtcVXC0QQonxRqyhQKC9Gn6OR+vw//pv5
bSdEVx92YyLJCHlEpfU+rnaMbWZbYMULs/ooCUI5Lhm9qCpX0DSTlTdHW1uIzDpn
hm9YqmN/iPYLu30dfS46kFQhLd0RPZohMdln5FUCshlMAdAFrYAEuR8mXQKoXEmd
6CY5tMQamNr2+QZa2WhB7h6prIC9eIPjSBz8r/DG6tlIIA3RapErzimT97me8MyX
+xPKmnRk2JsUYvEvHikz6Tb0vSkQnoMKn4XagIIl4Pu6/ekBkZXJEDSTyKmac2Ww
lZ/C2aVPDWTyv5qnWG7whbXzhtcz0ujc1GQDDRr5NPteULV4/PvOgId8jSx+6ovE
MMKt3jIv84I/D/6ov0Eg3bus73ll9RuFZCWzeEclmYnArEU7cZ2NBvmrX4oiqI3V
oDtxJrhSWqOb82bL/+lR8i1Acp+ZyHIwyrgTQ2S3aK41d28Njs9Ekci5SykTgtpv
TpHpmxYyX3491Iu9ycQiH6jtH4wPalI+rFD/3W/GP+1AfSuEyLLs2XTJZCQiujt4
NY0AszkKc4jz/R3styke32DE8nGzEj0k/G+1sBkAWSDANQK5waH6R4o1Oxd4Jsqx
Tzzean3mP9LYZqslexWP8/khBiK63p172pWnwIPVDWedhjVf0hVMRD4d8rCnOyWD
SOE+ajCbNhpr1xMuJQYIMkIRH5igobpYRWxIjY8C7gJtB2X67cUZQe0WNpSSyALm
fMfz8OvoSTgVKaeBPbocfQOkqJB83/nLO6qaiHUojgoOH+rq+wy6YXoPiOtFRegm
BlHSYOQdil9jT39IMjrjI2XEdiWex6ARMM//XAfLIMM1y1fpiosQEFDFmwluQvj2
wM2FOZdYX2xylDcl8Ii86ZV/hBxw2HNCLC02ZBvwDtMhZN661oFHkicpUH+jDZew
4dOkABMUSlBgbVRTuMjesOx0u/kFmj5DpHY9O7xbEQNQEAFIs1a4XY58YufGzsMX
azf2vR28T6PswOVjPXNjNiDmoLpOXslCgHWgTcS97H8h8/nxe2lHIKQ+ADszIx6b
8B7e8qhCYOMH2kv3N113jpWnqAwP3gAq0U6Poo9RH4w=
`protect END_PROTECTED

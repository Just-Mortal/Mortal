`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAACLspVB8ZssQt+qXsmmk5M/17Sd0pcx9IE4fcTBsDUMrem6pOSMSk92NkYygAn
Nzm70GJ0kujEl+sw1BeTZKRGXrIN6hZc83EvxGOs77fdy2zSZlTEF22fWu63M5Pw
ZBkRqGCEd3fj3WD4n9S+2MHSSELqIb9nV9bVrzo9LU+EspTE0Mn3PnR/loWvpUzC
VAzucZ0nMLdutEwjMVxaOGUMD3lv0certzlYjsuvdgVPdzGPJ3WoomjaZKzn8/OY
2TO+W44wjxv/nTXNQbjJH3t6Mang1VGJQUn0L5eVf0oNQMxcFu0XPcJTeA33yMuP
Q9JYUr8Jws6y9nxD9ux3hxFy7vV1FMENMZsgZb00jL+D7mP7A9UFxOUQcRDCThCF
uHMaiwg+9EAoC9bmtlBXd6eOqplfTO1k6BvKjI5ZcnwqfrdOA2uNdJpqovdwplaP
MBJmr8f9skpjHwYbKMRGeiDDW0BAfgo+OKwe4ctQbTDrc4a9ka7LLQU3Kmxzj212
feD8uHqzUgdGu/TlPWWPx5foWg7ixQW4bd1YfqgaNROjRTN1X7lppZiNa9tAOp1g
dGlo1DcetrDZXVrSdA9OoHpRWvRmuIiMRFQctfF0fVoLDU/ofMm7sob8KO8mZoMe
6GPMkMb4e/IcDEXAsMaPSusowB1orR0bM8gQtOvUJtuKOuDq/bRzXgT23hNNnsJT
vVoknZEBPzHPtm5Guu+6pKKLbhYOW5ec23GbxcXPEmf5EmZcduivd50mjOXSgKf+
WcdDK8+QEyTkEiddzIQryu9CkKuiD8K9cTBgRiH5r6ZaBL5lj3hl60TzYQocP9C/
vlkGfVdycVTaE52zGDDMLl+oitTpNUY8ngPK8u14246xIeZD5i7znIvmYhcVWiyB
t3pbtc8ev0Jp31d+PRrsiWozZye3/CtMRgxcgag5zkXk1elFpFHURliY4rjNT19Z
pu5Z5AytzSKfwhpmEzTGRWfuuuK2XrmMMVXSyLkgjKY+VfU1G2UtZ0Akq88/29CM
yfZd3J5Z7v3wn//d0KCHhiOUuqz82DIxKkWLfH2LSl0ZsQxAazD2JNvTszA4zdJ8
4sSSe/OIlS+CuETkAnjxmNxSyKzlE3cPyhCS2AJwKC0gnZLnr5OHlGLCYPL+RDF2
W/USOeRHWTxtbmsocZDk0rUkEZc/FWy9Lx4LmZ5BlZM594JjqbsR8Ql3NLqQU1jX
4srOEpLeNu/JD0J1QXI8t2DTTX0yfC6xawrw407qxBVo52PhcJwNTvHu+uBiiMWb
S6wCIgEd1sBN/ujD5rug7NZl28fJdyOpKb/kQtp9gc5WUeuH9x4Y98oeEMUH/7nf
dV6iWXcRDPq0jY7qBHqFRy6yfsujtQgARK8BC4HtHcHcIZoZHiL3dDWi9q+lqkOj
7aJec8Q2Zi6P+dYtgiKMEeTneE7DyBT3BVE3Gpz0oki+hTRsI7meavCN74UEdHMh
UAHtW0T4YRZ2wFqAwK1UxvQSIjUMhrT66C0zQgkuaVXXfpjn5sSqOcyj+H4moqXZ
sRW3VIh7Xh6mujc5zMsZ3lxWFQQt61P1dFiwxfhJDpTjUwfsGxNFRH3oN/9H2HL6
ASNaUw9uu7Byv2XMsvfWRZXH1Hf9LVNE/8uXYe2i8Mv6qUmUFjGaqHSUFUZM67Gd
Ywj3d+rTQBNsMKDshVK5Xwhwh58JPZK45ngXe5vwzFZatPx3eX1VxQ05tGHTDRMt
2RJj7OuiweS6z6S39hb7/JjaG3YfB9T2drchGZ7lXOgYOQv3sZUFzPowBqIommlZ
j4JCsfpcLnURaU5jNjpx44OOk/f3l/GnJufp9w/6jCo6m45wgHLx/3ylSzJAH/60
oZnw/nFqVDPr8e7lmZql1jR7QZRZwDes4DqOvP4g50PUkdwa+r22x8FAljR7wjg8
huGMQeUd2xKrbTICIvqZRnQhjhh7VTvBRjWjMN4TSeOAZ5bI+tabc5c3H7JU+W4k
NxyDLFselkmNG8B7yT98EqkWXeyj4V1eGV8k3uSNstNibZlqwZNEbCQlMWHJO1ta
6uZ8laUUs2nzKqpdeczm2HyPosJ9x7AiT3lqRMFLdvii9A8+xCxrP6akWIKn828+
lasq5js8AI6Ng94b3kGN0jAs831O2jEMiVISCRmpbXaBLyS7U83nmm+IR/GT523T
T5LZLMdAnA9pysTFhj8/SwPyplChHg8lK14bc1olhsiSiDpUxICp1YnHz30+/fWm
93huKqcuahvXYUfTbEMxmY+kW4z16s/5UwgdW2tkIf2sDHOcMoWuCRXMyIoQO85r
Y9zh85zDCXyyOPByc8AYRuVAnFNKpX6M5yZ+3/TCVVFj/mAm/XjDlaDZGjGE47CI
SqK1+F7fZdrU3r9LDduZZMgKCREee7QyrmVRi1hJ1/w8JjbWIS0+ibzTJ8tVs36U
bldCP9ev3I5/qCO4NgYoFlRZn1d8wYzTluJoU3XsE2lRYbiSoZJSrkqqJaYqtNGI
FRoFjrlAzDaRsU+7hVxJIOeoniB3/DeCtEYvKPTdACmaVL2ifUEisQDL8OtkHTrc
f2Y3lul7UcZIyVAZ6lel9w0avBQf2dQkcwsxGzWQlqsD6fbl7RYK1voHb4EZL3+N
pYWcskEVtVrpvkP+g+qRhiEEWHJ52RRfW5C6+byvVVbDcMbUd5zUP6CPES+gvKj8
MBr1MBEACI2Y6skwZSNWYvOTituIP5U+eWQjsBYLGMhvogUu4dx6l+IxMljp3wNM
Ojb0O+chf+Hc8FoIyIHko0bv7qXOiYTLUYr+aFg9FfMXyMa7ayMurVvlk2qUkQwx
F8llMdZ1kF771YXL5Qna1PbU+NFNHgTST/4YVOLzLtcE77SKa+KiUSymiQRYNGWb
j6JC6U2Ij3HlQu4/l7z+ctcy8VmQG+YYOLlAAcWPgs+IKuWJKT+GiewTeGKzg0iC
6/UbmGARzzdCJvePPVL1Z8QJDapwPVE7IcAcaWwPiRD5hZBxvMilv44p0wqCxE55
pw9hZ7KUYBeea4zrScuZywR0HjlFscV6kV3/E5Eu0JcHRwGV1iS76LYSftjwriXh
g3HI7zLGeHzJzwAWmAaszJDaPS0KxMkJT740QZotylnhDQnT7YASNyD9vZlWuYYS
6pFIU+ExxeuoAAe4kcB+3U26hUPhWIOSVueN0gAiUSlABv3vN/gQnLuuULc/E1HX
S050gclzJqIKQoHNfQzXLdpmqht5qoO6DjV1o+EvEq/YPc7UGUZKeXU5FPuYlTjQ
9luNx5BbkktYvfFC/WipDXi5hC7v4LFNbbAPdC80XJREcMyLDz9QJT/Ti8gGdJLa
aC5yxPZHDpj3PvVScUKKYWuW3r94tcpnPuzMh7qkzwZ5TzisIQ7YUTf7UYyinW7a
n5zmexuutMEGdvE1fwQympH27K6C4OHMJidC0PR91kf54M/9XwNT7Y9O9Tjctpq8
BLVYmvwyQAG9ChfKeBdT5DL5JN4GBKGkOYst6zdB+5TfwM/9q1OA/fiOPAXoyd5c
GF+ED8OiN+7Z/sqBQp9uNgkrlx1JZL0JiymIlwT9qTAkCcYrr9VOogwERgvbaxqp
ByS85DkxpX+fHKvy6GnuzQ1GkFz0jNW/T5pfNmuXc82ef9n2nAhsjEz3pKEFdA1V
Ev4BUVPxI834vZKl3nf94mHXXfom0m1RlsI9CxbNBi+U/vmAZEmFQtwnOs9ZnFI6
fhX4B9DtvtLi+XDbwec/oVembrZPygpxRYFkhp9JQxuWia+hQ8a4cHjPRx13omvk
ZnCXZMW7XSlqdnyGO5hTQc+V/N1h84GjOdjB9Y2Czvh5/80g4K9+R47BWPlg9f1N
nrejWVLYV63mx6oCQEl4mBnJDDFoqRwq8kw8oIKV5WtRy2krDn/zdENAJLjClVZd
l7tBSHDM7m0O/9zC7axsoI9xG8tBTH+9NOYaWwYtJe8ymjS4jZhlmFs0dl88vg55
el5h8scdYUPfEdDZ7/lQnZor2Eho5gHHk3Vut5M93R6S3pYdzqaRRDqrz2xxh/5n
E9tSOFKfIkh4OBFiXyjMGiyIBCywmOC1lEafDMXE3MJt2cIxQYt55g+kyVSiOqVp
bySPMzDldTxztRmywaKN7fHQuPIdU8MFvL2LGpTnDW873Mc68o3YGl+Vo1OQGn7c
bF8fCGpLLDQjnGs82h++uBo6Cm3z7I6A6qkmaT3MmYpUF/1CFMSYjO+bo/xx5JK6
8buVcROMCLx45iMaH7Z69JNjrt3U5G/VeC5xlBHjXzePKlvBqib4fr6rA6gZH1xH
tpTg8Ua4j2WF0x899k5k/5pXgvBNg/iwK4dPw8c6uFr7jjofKWRjn58sgR4pExlh
lfODepnwtgMIgZzyc3cJPHUU9XoVZnTpDjdQaA4UMpGcrt4DXlTU3ooQaRv/hOiy
UA75TByN7gAkZ3hHlM3ONbYN7WDqfpoxazo/PH2enbKVTek39XyZrF776/pGVG/5
mME95VDHX+SlNGWH8UW6NrJz95wO+JooXNPBfXQ5YgE5uB47HG8aZetz2aGRzm+i
vC9XjcgaAqRHeNIPBCLKGzZbiyhEogIbqfOhfT0qDLzJ6nVZ3H3PGE2A27DcL078
iBCnhzr5K62wXbNsXUonwB4OHd6IkCZYAY92zp8AD/xJg/sMjZccf3BSCOENGKQu
S4uPOAixYHlsS2gOPy1JgYbfVb5Uzo5VFwdzpIbAWLy+IrU0yRuQyOUKtliODywp
gqsNBiLnGTKUUchpaiJQhl0L46zS5wkrTq4NlquEfrFaQMRlFNUjmtlS8HOJ4FR+
gs4/HKJ0E1+QwVK5s86AXEJLc2ygiHzyLp1LBGxKUBjKnIkO2n+fEMaGu/w5oxqE
D/a4REsChLRY2D5AgRdTgZ6+3DSV+CtbWorqqAi1lXO7sVLAnsr4Rn0XcOgdkBLE
7Go2ozM6nuVfgjPP4C7uSJBs9v+kNQbaibAWP13EK1+A01MT8al7PvM+2alz2zCh
Fikytz4yba5OXdci2Zy7houXmkC2ADsEEwAIen5EQ8g0ch97XuYbHxtVt5ncOUdw
OJwsPXClKGmdx+k0TyNKK+JWCebybRrWuErrKBaBUmHLLojUiwmx5mYXdbke2BKS
ZfTLZ6eP3DQZxZa88JWizTgkgd5zEJna3+ccoSROvZPCLcNICbUkKJ4oy51HLMOs
PiMpqe9PR80CcHKhGrkJsf6mtcAmF2DxyqmdzvsL1XMwRyRMDCVNe8o2h90TLrYj
AFruUGCfaV85vIfkBcUdnHEjlRWiFrV8ndohhow8lGsf2rsV9Nzp00U1ZYg8iZBv
p1yYCoytfAO/T+5Th5bSEvD8ezvjwKkOgItphbmyRKW7w/JG7NO75ENb1l863tBs
bv61xVqVYWH3RuRmGqNufYkrEyudBQX1Ju5a3uYiECeu9p4PRVfOTeWtFrDJgk/c
ug4WkiGZRIQqvtyY9OXd27aAu1PG0ynqOjOxLOVz7wyt3RDTgXXnnPswO/gFUtd/
UwLL+egAwWzqg68aoBNmUmxnIX6czY4m/tpcuI3Q8WSB46xz2Hz4DhVtGdfCi4tO
T02/1kFQ5TZwaB0eeobuamWx2J5jp11oXQ+HvVwDdCFxeXlLmVeO4FcOQzjOz6rn
fsYyligCSbSDBhfn+KHKdztEeo3ZrXya00u9eisYYig2hs1ymaVd2DFiqzAC7yXW
NRQ4h4fsQxvxHEiCqPEavzkbJVH9dYS3cpn1JIt9Pwxx6AagRp7xkX1+2bbvmc+Q
R+GVcsutigUJHYNbu7EjbhdvU4UCdzWco+KVpQOjlB8KeM9ON62VDaLZ33RqU/bR
X9zdk9PT09qSihDZaulAwpIP7t7LISKMufl7r4VosGWpYbNkyIapgmJGFZ4xlDhl
Ciq8uTj9j9sTKOycNmnt+pBCXTTZYNVRK8Hxb87YuXkj95kPkW2OM6tbSQ7W1Zw+
F0IeLt1MjQyLwtk7jdCYit5Zg8nAsLsd8Wmfv5NlK+MBzlkCmiiBmnU/8EiSOjeG
datM+28uDDv6bfY2E/vnLz3Ajy0EHK0ybgWgajK4A5+5JJE37Qm11rjr4DQ+HWR3
7FaE+mIpSR8Kwg0pr2bRcacLM21CHSDAO8HE+gx38o6UYUGyXGYVES5UWwFSz8qc
yleZ7J0fOnToCE2nINupk1H2Y0khYZnnz77d5g4jAvqraCAdw68lquRQhC4JvnsT
Y/BxWS8RXP6Bgrim21bUQ0q7WZv1qhMr1bWZB728JvjjN2MRXKPmZgN/zZxPP5/o
WBU/Bpo4qTSFqMMlv3D+DJYVk/KeTsGfLZZvXQbhxqJVxmXiKcWWmHq9J6k25+O2
b+rrvwPKCqewYM82BPQOCSbLN7R9qXopwzHlMBRtJ/3PQO0VJaXLCFzbFx/wewK/
qP0Hp70Un4oOQaEQT/ngB5RLZp1pS0nnCPHZyANsrW76pl34nbcdcDsCV/Jg1kof
pO/mZENHkWFPdGH4atqyM/XuZq6RatUKvOaEH3P8k6oHjRV+Td9knaguIcbsnIQs
dKxbjzjxqWMWp7JG739uhQrAWEIO1kke27eP1VrByTUzPpUETskRQlGtjSMYk1hw
2dOqoan6fdC+vWv1PRL/R7QcHp8VtcRTa2uGwnkzTzwXShzKm/i31nf/ui1+Z/Ws
CSIOlHdXAa8zVZeH8kLxlV1Vm1CF9k3ScKaNR1X/vo9uG9GzkexSA5jy/TJnGII6
7KOYZRY5Z85O1bUe3jpdQLM+uMuv/t2jLp7Y3cbageQLilxyI3V0MP23nPVw7hKI
UFdO30SMz2USyliWhlrOGuRd6Vh6n2hZbgdJ5UrC5oN60fDNkr/5nkmMPsz+bjbP
waailkmYXfgFAPVqy54sTisKWUAx4eyQcMDX52uJSIijVAjfAN17aWeIhYLfC+ZT
ZcTCbyHOVko9c57p6kxDv/VFydu4P1GIjPm9RVUrFY2nCMc60E/daYUMnrzzUfbU
rY3PI/5g+8Gc/lPGEHY04zUMnntyxiSyS2ualKpSJIuCezhNdUiK5ckUzaPC4ISF
KJjIeF9x2Yr9Iy4DGTBEeBz7PdcKK7Q0tUevSa6idPZobGa73Hy4TJSwxZ9l7xuu
jGxZT1bvdYggdW9NJoQkJaTTUQecf0MXLZ5yLMUsm/3/AymrS6DXpY199+TXupFY
IeIUVAFfIp+MmvgolRkPRc/WO3QmO//wW48/yo1hQ0GsGwVrBcVEzqBMMcZMXg4N
HVH5bHDCksEwlPAmQHgQgQK+S3yNgQA1aQvwjSodmfopvNUBcVVGEQpeHDHMBDV0
eA/NSst3NgHDtTRgeR6yyiPnVDpAn5pa0uvyxyoEP7w4AGN20HEVObCmrJwYou/a
xFo5GfTnlaK6wWSpVhfcfoufu/nEB70OJ48e3TkpHJEuL/po9d+ype3Rl8aW8iyi
0eGiReGUVXmHVIAi6BBxfA2gPoHsoVNiFbX0HdiwC5uYnznd0Zc26otHJCmthk4E
t/DT5DXVGE5HiLeU3v+9DJNHJbMZZDydroL16KtfforNxy+sx2VK5yhwDGxmoakL
WxAbhagVrWj++AU/o/0runF2tZb/jbzxLcSCSHHFE2jhnnggwC4N+o2EsHke+iT3
ZQRxIK2NJZG2vWrCZw5Ev1Qz+nUf9WFGo1sCKn1JPjR+MALLz1JiPKtpNO43ZvP2
akmHVe8CmbxqDkQjO9rdCYo/T7ttpi28G+LDDpW+HL6GyLzz0+muckSZVcJnLPbi
s7nRaYBNIeGWQNy98m8Dq0APNw5s2UIihn/yPEMZI+2x/mMgSWTqM2i9iiYdjqxL
ePQNq+y0JNs76wuF+yje3FTCbS24M5XsTBryCB490ouHDqGwXAVVKSPKo2kbIdHm
wHvBCEfUEL0r4lJUOJ4gHXPkRzQUHWnBPUCdK0GJrHAV2/0mlh5UR/P3YYz/7yuR
I71y4XFRcg/3j9KKJpoFlUZCMK3HR9Ds1h+nUj5O8vOhBXUfZ6Q2vA3wXmutqHG7
+ZRTpzDJWsuN1uz3j/oH1K4geqaUI1YpW4n1I2mL/NaoVH9JG5Wp25eyWBacUVQT
JpV+ZO70SI8AwAoHukPY6h5Va+RUb0erVGCCE6oL15H+qB2pXrQRx5ERLeJ3JkIJ
cjFwRf8v9kv0v+f8XOCyQ/b/dXg9T7v8rm74hjbVL5f+8qpYyyi1oXVcymMueMhc
Dr8HpIGNXw4f1lY6cVJPpNA7MEt1aD5yyTD8BspHxrvas6hahT2U8k8cLDxKIX9V
dT8S8lLR/xA7rpES5lJKyphQUQGw5hIrHNpFT4HYDn7AeusZtWA4CEUAeEPvWyAC
w0RJSkSrgyeOKt4VD3Jw54aH48E8IbxIHKGy1KM5ve8KYRbrUzNgjdBSSYJtgN1E
vvbjWDGbhT/UwM3UAAEKfQIJiQNf0QQvxZtAMOQGCHv2HJqmSd6/cue0ETrBbvNl
KPwM3Ku3LZdS4BvU5nAW1KLr1Exv9B7vZLC/HQ5G6VizwGC+dgp+AyadSI2HxlCc
HVrx87ZwKv4zeAvMlnt84NDDvwZA1BIEacLH4KI45YMr8QAZxFkAHp1bXgpO8AAD
R2dytMKE5PJIY3tKRbydE3KrQEX9XG3p3uI5tHMqx5d4pijw+rFt4i//kYOh4S/4
eIgIbjFjyTwVHJRTA00HgRe1GxRWPh4RXmpaPPaXRDltuhVVNB+mt3OHBsuQo+zp
NVyS7yu/yZqN3n1WQuIb+/SfIZQ18R0rwnTObffpUscvT6xm2shWApc3M/b4Py46
LEBMcMs5al7Vr++PnMdg6XZ7xeLkp9hckBn7tzA/tOCypZzXvaWFhO635MCZQ+ak
XRkXzILMWnUytC0e/hrvmeOOJ0cP50Zp3LVoTvFT8d69gEYv+oy7+OFXtQo2AfMr
S4bHLCgs1QHgHjxP9gDj7ikXc8rvqrZ3wK4joa1z8qRSDcC1+SFjPv3z2b3+rY6V
X+nD5/QmeEQI39BWJr51a2IXd40ooouTwTBTZoRQxAw8d/cXIlkL0/wTq/hIAErz
vwcaQjsJ5nXXkC0WjnmA8GnMAL11zoybS15ob1dyE0nvafN3SChZzUTMQQiI+Opb
+35Zs4aSs4eZ06dRXWvEOWdiG5FasXJ8L0o80oiOrdMbkwDlC8QG0Q2ciDYgo82b
2Mz2fIt/PWEd/ESQctkqPcTZXIgx7Hpf93XvTimSya+UpFrW7B2fxBWc5QvlFQlm
tUqRoQRyPDAdKERVeFIiq4ftMy44uXPqAVVCpKISkactD+b3Ua0QfhooGYO7wNmR
mf/HLwuiqHFMXWNjdk++1GojNQiXeG1gIFo2pyjGMzCbysR56oSRTXSmWMADBX4n
IyHSFZA4pmP8mPZ1yRl7euUerhB8eVjbhLnRsCjZukEwk2H0P6yelbDO0Ei2XNEc
F3Uk+h2vQhpT+4mp5dm3vffvJDpHpLMYHQ3Cc3w4LjvbfHRjjoY0cZbjz8wAcY4I
vGaS62wWce3J/wy3i9Qab22gTAlU5uq5pbiIApLhBjrHPdxT9ttN4Klop35WF6gD
tB0XvTlGGFBNRY16wFz4s04vFz7u0JuIRIR/cbO3w7XqIS9q9BSWbwzzaYT5JDjs
WZCZNeqaEEqkMTMUvBLqrdhtC1NP1X+weatggfufqe/XTqd/bfPOkeaE4YIOB0hp
4ned4JUc4DS3E9y7F98cW2qYxZcvAogpqpDVLbQi/UYsCXUf8viz+lIvwpKK6fWu
CWhx1cvPYvanWPXB3YVMI1N36JXPuPTYF/ApQP9jmaAjllUoOPR4Yu/ZwqeS117k
/tO8wKrBXYoIK8AKHtASoG3x8s10QlObF8evgWMVTw1ntrT8MJ93gX6hCRN56Fwl
VMwEmzzLbX9AaErqLqHblW/pZyHGo7SiLtcy6N2zyVyHtBnRrAps7sBJd+DHaqLK
9jZBUB1AFOui6vPgHhSkx0jrspiOnnS7XMJT2CdD5HGZZHQMZu55Z5U/z/FNPup6
bxjX6BXDUb5I6LKdlq5Nc04aa98i8cAwAO2ol4i62F3DXvX+xdP7/AoSasVxKnTh
3tBAcpCviaqlUS0pfZww4KWKKXEhEqoZnmT4/0IN3Oq+xur8fqpm5u+d+IuAjTZj
bS5GoLvC1qofgkAHzKuCjJYZdLu91RCTZVwNn5bIruk/9L1OtH62ynJNdbXdvByX
EgOvjFlC2iS5lPkjBJrTaXlfM16N3kigOYlIzdE6ok/s1VGau44nhIEhZdSxmnop
UIvB/pZl+McapMqssf8FOf5Letb+HscZ03xotYcVdM/D68Bd5OsY7iBaMeMYg35T
OpD1lL/W9mnVux53IWq84Q4UfR53dETHio8cJxNMmu1G3YcDJZkggB0xcH2Akkb3
TsRPq4CrhHx9KMl9lrNy6uT/zHNnR4Ba/ZdNwKOk8CIcEeW6paGPd8QMYvR1rc45
wYL7lw2grxHWoDHOqHgkvqB2+PvijVKUh7VHMUFyzF1OrmZpEZPnz2AN56hK4p0u
0jgR2Hb+lbsGrp3hafaOwN23L+vClVOneICRCN16Xh2+T/T06RiXyWNduSDl9U/8
ghhUyQavJo9aH5zF3VVaQxqRLwY4wgz762l8raOGPkkMzmkXo0+/3Euwd11hWa8v
9KWHWfc1GaQc8oxBOv9U3CzftIWC9sYPJRcUcfdJAz+7Lgn6QTKGyrTvlOr20PN0
BGzOe/F9LqstouBCwvkIFLdbjqnmkQJaBUnvBb1R5AmxB21gmDOQlEtB7dEokfpZ
gKttdiswDRjBIvNctfZk1nsN7zrZBCJv2YML3vs59PHLa0D6vLrQoTbxq7WXCY0P
Ai0M3zFSuMbGDH4AY1nZWUv6Ti/uQWlksXd+ArduDw0RNAnEyfZPTYXvf16VB74q
Di02cBzMAAqh8XNFVEaDnSh3KWd6xNtRqjZIYxcoDmZgZ4qhgeAbntrWk20K7tyO
GNTQ3fdCNvZgTCzaawmFG4U+veJ9aEreVywLfqDLkKC7mIbvh2/DixrzEomQvDXP
BT2Vp5DnauKBVdypmR9Lk17ZpnTS27OSz8cPme9V6mrvEwt9GndnS7++e4QiTGUj
Pj+M0mDG3w4mHodzEGYeDTYHpzlrG9/rM2uB2KqHDHRSP+2I3MbvvKJvHChgdzt8
SQKDIZ2/qd+uSOCX4YWaAWnfVHuY0tMnjYwib/3kLR3SuguZInQBK6fSw7F428yR
e+ZObEXPKJXXWNYdRrn3VmMeAyoeNMf23o1P4bz+yU/9jToB/F38tdBUpG/3yJ2I
tvqs7szLfOwpkx2HQS8ecstwE7srfPW9cBuYFT3n8k75uUJ3ZB+wS2CkSfsXQdkx
DxFO1h81Sp/65wShU7TCgvav6yhQSCd4zQq93m/h9WxU7e5FlW0F5cpoFrWKceEs
UAfzYCVKuwX8iFY1Y+wqnDcahoBZGOuqzr9jHppg9HicraX99QzibBujKguQ8mIy
Z5+k4GmY1LeembZ250q9yD+RSMisAjd7cCHtKb2SSIcihCiBpmStK5sq8AUyMPCl
5JEnzPPYBkv8ktvxKIL1N9/GmrlZ2vxaZ8jViDTawxUef1XgNHWFGUpQho7+JdZt
0bqf7pF8qn35W5qWbaQdHNrSqg3a/e0tOasc7KGCRoPSPmZJweDHFQqJkNIxKFJ6
HgkWx5jmJ1SFtgI3V455Ed15vBUqmpqErTyByVjaXpKughAoONXt7ELz9leEmQRM
rk5usjNsiiFNmeMKUsM8a0KR39owPfpOwKyju9yl61w41stpfGbPBWmplNh4pK6N
VscCucP6g8YePj3CVA5j4AkG03K6SF29sMxmGH4y2uYEx2Okr/iy/YSAeEbPpwmR
NI/0tbfQK4GDiV73lFTaOaqQ6AlRleds4y23R41wjaCp6BPFbMzpQYbdK9CmE8HZ
A3zaNK8HZLsb4xPTXDtfTmItzCjUA8dy7o781GhLAA7e9EsrO67xLJTav9sjmmBV
8KwIx0ClFCnwgil5xg7yx+VJJsPkwiypmd6pBcUUwTImg0WkI5oMyo8uiqa47UUh
uvgt+PhHnXMaxB3ZPNaHxTrfC2v6HMDMSBAvjxkZHz0f3vL/hkbuJJVb8XR3kSrt
8U3wwvyjku611Nv3LiN0WdK3Z/nILjB3AeHbhbLfg76f7Y/elUOCfRCcic4IHacI
94nsw/FcInyuLOS9Q4gny5OCbc+YejoGxhPftjaf0mggwVAvxrVc6PKXt1pAsBlK
R2IlsHEEHWcWqvPaelPaSliimUnHofsk5uMfrhVp0OJJPO6CxDAQ+M9sxkEihDKb
XSyUIVSp5tI6+JqPz43j1AHKCMzpiu0ZP7FOp/ZgIE6t739ppDRr+mlkHZo4UGmQ
zldtmd8ezPjQ+Y0mXCTRkI1LzMn/m06QUfVI8qB3i3K4+dFQkvCWTn+YL9GQ2mEH
DIDqurk1srTjRRXWQMNzNdA4SBTi2tMF5n+97ozSY3dIpMYeO+IpaF4St0SBI+/p
Ls2ffr6oq8iRQnmSL7mZQUyHe271T1BP/jxE4+tpOqlN/vfh58ozZlKwVi/1if47
frkoIfs+PTd7lsJJw7a8IktTGXhW20tBJQFt73NhJVda5KTPk/tvYOKMrmpjLfSh
YVjcNb6txf5SSn62T6C/oNvBdc8cgvJGkhk5D5QO7yYUmgRakBLhtfJJ+Mv2w99q
6dDBuUlPj1l+O3LTwm7kx2X4Qr1phASzRIhEO/7rxN/K6EtdvNY5/o7SCwBOj4k8
X6kYNPedf3LBoGWF0rlPyvqKJx5LOYxIc7Z4dYI1bbVh5P9EFNrkvvKYL2WpVFUP
5428wtHpBFy/zlCpyuqN3x2o2FsVdkJ+fPK1eQDKAR8LP4pp7Ls1AzJ67WiFoLbg
5nYgZ+h74Kj7QBqn71749IAEekR+MuAgNZZKl6DwzRocOwSauv3nMt/H3e3i7sof
ohSQuzkArHhSNB3sTtXZtOzDYtr9MX7no2bao/wSWSwS1s48p68+pAwfg3gu2EN9
HLNVdLanQNnlP2h2SymXb2iwqmYxilefdsrWmc57/hAKCBuxSbEUpS8W4BMowDSY
ko+NInZSpTF+0AnRPNvTM/BGhD7pl46oEKZB4koMgZpHSOTiHJy1IE+JN+JJ8FRf
BJUgidv6Mz4SOB6VIZqZFImv1vTDk4D/cZCNwy7ccUxnAqW8us7xTVSW0vw7urDs
H4yDAfsLDfu7Sf3KADMoIU34Vfp3PP+p9WQmWqkQOgJ6hLFuyxAUSREA3/PhXPhX
zPWLngz4GISYu/10MHkxLmClf4RHEb/pV5AVrGS6sUavgm8DMAKzYroeM7rHERc9
sh3yNxoGm/XGNg2faNRsWhsKGLAbvRAXjuK1HcE+j9dFqhCVkrKLVbPGR56xQmce
MUSxOrx+kGjG+EvfazY9IoILVPFVJt+ez8fIA/pCWc36pVTtxdBQnD8qD+vpkCN/
P5OHPBOzltqGDn1AVc9LCt71aZBNFryqzS/xFBlI/2pWYuexonfP/UWFSh1Q7L4T
Eew0BpgiUCLoPhcQdK0BZie8QsXT0jgVc0EuVXlLxBiEOUgt8RDiL9WKfwiUWF59
yPv4H1YFArC69ZU6hkSHXASqXW9ZzyyaIf5X2jthd7e0LtzZxJZMXc7nH3NB1TrU
FC4avw29vz2VmgPdpWhgE3XdkZ5OoMDIftIYd68RhRMzckVVRStLeDxSN0hFS4H8
pofUNQuLUiDvCcREbHpXEBsJ4xl+s/vxZVBuUCl4co9ABvg9iAOd9vjfOCCfvLDP
8qC6rBXWtfl8tl8G0FCmuUXugTXD6I3iMU4h7wju7hZ9OkjegY2FLkp0g4hXOhc+
FVh35j5gUFw867H3cjPB6d5FYf4Fp2lMLjfVgoE5Bw13BjfatyejMIdYIA8dKhft
1EM9Kf4XffO2Tjn7Z0fSrd7d4HpldxqN/+7J1MGMA4J61grn7TfCLCfYdDimmEjD
YZDTnfp8th5uvDPj2BM89rbkjccyC8EzQ1pXqdsm08uwoy79nIJ3/ym0m/iZf4/V
Xd3UdF7k/04ZbUYngknNfZqnI0D/Ac2u5ESVjU9scM7Gux6WNo50MPEyxGOMWjmi
lzGool3HlSEc2/ntee0juPSPJqKKLakqzRvWMdUk5ezQMsVd/EeZgplLcn59ARWO
F/ijnDNvzQhP/R3ic5eFnnoxq/tqze3Ir5EE3WC9ACPpURhdXrewLl26aiXJ36nz
JsJPIF+9xjgeR9hT4+2KSQpXmMDO2rnNWPxzWuoSkpdtYhWsLePUaTyucpMuHgy+
hFCs7lWnUF8+D65dIa1/7S3WHmtmBvt7SR5KwGX52ye93iGkK9caZjNiDX0IUUDo
Ju3Le5fHLUQf8t0oASS0BalMpYu0EI5IgIsTwJ8rc6JGQosMhQZhv2DnnHcUPIFM
W//kvt+oKYxV6wBw9BMJHgKWG6ee/imvS9hJW5rb/RH890Sq+eLvA6hkP8zBXkHQ
Ewt9Bx2u++x20nG220ULlTmyjJWW9NGeWbVmCzchqBBqc0qFLlQHBeo8cNBJ/xaO
IulKrgVGfkRfSbpeWC+ZB6HWIzwT3HzcUwbtDqW7X+GbBJyuCKaTALmtgitc3OJK
eV7zInurne3ERruK4vLRlH6xZSLfMTkiDCdUGUcRS1g4BZ/7shbYG4JYBuQ/xjgt
Zoyk19rdaPtQ6/l2rvrqHVDwLo679vZUwTOYZ3nafqJICkCAFmrhNLVLFw9IDRmb
J6zPQIelWdGNTc7PHnHsVQYEUhGRTO1TfCugI4Rp22ryVUOj4/6hN4eYaVhDVSqV
cBnVTMlx0ldrM9juuNUr/5YniXgIzTDy0ITAAEhod8keAU/QETReF1fVjjPIFE1Z
v6n0Q0i31QMloVf8oIgbmbZO1PdDKFoXs0CIwQ75qinh5fobK0ZWzwSDtemYY7kC
+BAeamJaiopMPF+4D7i+oVDRIjNEjdRJRBLaHA1Wh9a8rx9R8WyCRPcBgvonVoU+
QbH5cpUX6HoOC8fcZxNvOEZ4zGBAUP8KD4Aspmaedg9ZCJgW17o3x6Td2mdQA8Dz
Vi01lnVRtjlFya6XbAIjxt/SXXMReinSHKm54uKRtsyYyRJK2Eq/hf67SN6ozHWD
pZ9oarawVqnwr6n2ttpEq7smhO0IQRG4icbjzlOZ18gJFsCIoqSdBQuAeBOH+lXT
ZH7vEuMCmY5Mq8DqxZDJGdFeJPutZ2CxTGWSafE/yQx6iiycQSIK3W0/XBpq1igr
yPCB6+uPKmaQMcv/wUDN19H0l5jhYTn/bw4OSZm95BYP6xfJjUKkNvnf64Fje4yE
yxTZYfAEuefFdtlcjhg1yT7AUFfBx36JulMjJRj6Jv80kX8bSR4HHBCN3ni/8Jz1
3kAsl5jsuurymcEL7diq3tyBqqXFy0mIvuDfcEb3Bo61rjIdyv/rN4+x17XOoYr7
oXOBOGj3Io8skYKjqX5R7b2cofnMBAgYPWnicN50unSaB1qjghB1zB8KJ1PRP44M
syKBnVUmfavotUWmqN5EV2Zrfeh1iamEvmt4KqHvg0wFUPHC1AgvWZKnZ2o/VVO3
SJDo2oBkcufS+54vvvyfpFQcZD6W5S5M/SMucH3EWzedAoHoEABDxJqgckaJwGZ2
w5RVOIWjhKz5gbUO8iR3lHpPac7yFyTnMxGrUbla7XM2Qdj6doigxzJ7Q1Z+6B3I
GLXCBQBtaJE6Ckbu1rU61Qk80hg0ybiDKvqDOoRyPXdOh+jjGwm3i+tLnViZX+Ea
jMEJr807JG7c5SPgqWp71JRXRXgrTfT1HCSZRAJfLuk8YqOLVIEahYvIZ+V4KxZW
bwfvRUoZVb4Ea7lPyUwSeKdzDIajZ/rFxCVrw8N/ukfLhgelBGmP/R3sLB/87c3O
e0lCqIWHzHeVJj5RrqBZd7kRC4+I8IB8AmRfaLazTr7idW4wZJKcAmwSSfPwcKi3
8tF7nqLNBwK6Ww9ZUOGHojA5OQmYPazhhSkosFIbAfjHep/tEF5Q+KaDiE9fbdTm
Jvy6b8tFMhzpoSajCN+9X/UmqegPZfAl3ynxsnt3prMaQUndHcxSY3l+gXxXUMyY
TrXlUGljh4xIVtwzp1r/GYBXOBpVbErV+fCyIFhxUkCN+J40I8+MNQkHcCqr4Xn8
T8VHbmNPgAO+08PziC2CHCiADylVs+lIifB/k9YhdV0hRhacoBeKqPjYdKDAdVNQ
DlGXkMhDbAehKnR0x70D2o+5oWMv7TB++qZkMEBIkPq/+iJnqfe/Fn4QwAimSyKk
mTCQcuhruWvZm4D+RLn/NgEJSF9wbVql8tmtFJZsVmwJCsEl0q8CaaTtwR+Wck0o
LcDAvAN6WBt9HdAq9M1jsaog8V8BFleFuxYQMnScaHP/wzEhhaOf67alL4JMXsdi
lNYlLPT4bT2rwgaSdyaq4La6mEZXvPIPN9JIWKRown2NsVJuZcnKlhFfiXB7fqtL
iKIy4oXlliWQvyedJltxYjDTk0EkvOhrEeGl8J4Z8HooEiwUF16bzUtqjrjr5hRZ
bbKqSnjIlSmvYbXH5IOpjKK0kSQ8CMhFQIpjL1CpZkxdzT5Aj96CZ+anhTjKBz/C
s8oViK0+J8evEphjD5QdaWkhAr3/Y2T1UBWxWM2zT0vq7IOILM8AWvIYHWgRO++F
UGZWKbPemIqgKABrDDyPa6mnk9GwttBeGiaF68kOL6iFNrKodr9QiH4n5SZpvflE
aPnlj2CED//IocmufaRLPotRr71AOXPrBd0ONeiT09Yc9WbBvFZ3pUmBr5u1z5jg
4hmj0L55POpyCD70J2WzXzH2nVqNVO/xlKdtOGMcz7H8gIdauNCuMQWodx/KVKiu
pap1TL2zz2JSNHkStUZr7vUMkSWIvxiuNavltKheYkfKI9xRr6ZnpQG0xmbAWFWO
7k6kIo4bMaJehe9XtteXd8asYiKyd7Rf6UrsqEKt7EONxyNk6+4/3GpWMUjFdMqu
herLNw43QahYhyav8QjkfSut+o+yLq6RCz6TkGjyENn7mK8cKBV+46y/IYfa+dGL
nyX1So2k08VTqlY/aO//S7effM0mHHirGJr7JtfQY3thEMt9HcSnFZlAGhbNJqee
gNPVginK0jhileamvjMvPReP53G9d/Td1ubqSjy3uhb+t2vdLP1hYCtww3ZlFnwq
uVAfTkrvHUARpldyK3j0FqRE042LxciVAFQcwM7hsOzhGEBUSVWDkVzvsApYmoOC
qzR86olzv+xkMlaDLPDIBaVfUmYtykcdwoet4yEVp1zsxUsEt51CE3KiTCPr6Oys
mngcG3pfc+tFride3raQ2M7+OOgf+Dp7qXo/R3Lw3bJcHvZfjGAQn75//wfs6yGQ
M0s12i11rLn+prLdAuNK/8d6jMNHhoZmUb9gIIKrmG8VZ8X7HYLvXT9WxWUjY3KN
/FPhmkWzAfLdznp2Z5fLmXQJG/LznFYBfFa5L/5aIQEvLc/n+OFgFAV2VMI/k7wy
ZNZHpRsFrGzlD8fJueyJ4DGEL27Kkkwiv9caFtCgqWl1/EOjeLfz/3Op9ukFz6Jq
GdYjPsb9BCdFrwXC2kPtDegHLGXO5xDDRx6qcoxNfLv0EIR5C1bzQmg1BKcHe9Dk
973rkpRrXT+TVXeo1Ns/p61rRzyPpZR55hkUMSRpGOSM/fOvuDfVRDx7W9JWy8A/
DLK6xdzdGb9idMft7IspxPJcXgjVXc9fJlhgs5XzbGf40mH3QoVX0k5BX3ZmGAyQ
ot0nwJ+wUa4siTTSs0QzIINiER2TdsIEAF7RSjAJDpxGVmnapUu3l7JqQnFtabAT
dV69EuRZUKL3QeCN4/oZG96V0CCjgKNChN1UEwWx40OQxfq7Nwn6yHH9daNWjehb
OIQYi386l4aHReNl/RWkvmMJvB8ZSyyIv0ZW3fIOl5O2t4SXp3c1AWsDflD84VGl
5WlzJWs0ZSrN4JFDaeElGHsBsmfM8q+yYq/IhfP0mLjUfY0z+QTktLvFeZ3F/WSh
jSELYEDLaYRx4jbo2iHYQJizpe4ykhlJxkwZtBtxUA6IVoU3QWXPxtLXyhKG6f4/
MIdK2s5sxx31c4L/c7/A8qFfkmWTLqUbf11r1QvmY61nhboHItYE6o49JDyduiTB
CQCNzv+59r336bDSXlKUTrJ8KrO/inB6xlQO7JEw/cPibCJly6ioCrCvrjgHHuc9
pUsaMEHkaJ76sBx0Dby7W59peGbJHDUSGi1g9p2u5wlzhYz/XajC26Nnn9bC7/mo
wLRIW4oRWb8ED+MGFV5/Gnq12+LzMrXDqQvR1ZdBnCt7tv6XdeNk8Q9JQUGD/oxK
Wj07S7cMzIgmqtfreRnUGECwMR/1Zxs2rFGSBB8MrpH7VjyP37I0VjjUBvp9cBFY
SJo1qH04mbschgwioGh2tQ2Cjy6RBiNEC/RJdMyXCRhHlSXeaGjGDUQh9O2bzFwF
VOUNmNX6YH/DXlYQQxsDfVL6pBrfakE9tB2Jg/HHI7rCAM7sKHLU1UMKLyfMvCIY
Vag2u4oQr0x+b6uL810T1K9p4KIDdmny3AoDxmqALzvSOH5Pw/WMWu23FNL4oEOc
Xc89i6PgXIDDtajg+1Ks2j6Rir2rT3KonXgWO9glp1iCBP3VV0284NxXtZLInUSs
0yS5mNnQVlM/ed90eOsI6uNTO6hkZxe2C7BCIvVw34MRAcBQDcIbDx62tgNnfY+9
QSEsRQNV1gRUVa9V+FZoeizHvjZWndp3JJm8xeZdRMnGmDcsgCOL3GkeGdsjS5S+
uXfIFgCVpbx7hfRtI9EGhV3sBdvwUoRYgdCADZgug4pGQhtpflHOXIAZCZw/LTQO
r+l0mVau7E87ScuMUcwPyNhdRVvxFcvNZoqthrYXV4ktsdeyUwpc3U3XOzAbQWad
3p3EXp8MI1yZNchdaNOa9XjDdNhqizjSDpmflnR2JodKUKsk6PgZasECPkW6Ogm2
758yFHW5nzVmaAiPfWDAt2Y/XJu9us83wULeFwl9dyEsBWzj68KfuSJis1zMP/xu
BsQ/Yru9RSX31nyBXrZfxS3LxxWnEBw3i7yNDvHdFyrHatIv559m9xPbWb8TSa8t
aazZUIxCLsrnkrU+3Avw6VqPMVb6tqzcG121+IhJNTBglJV9PU/Yl8f3ofG48JSd
O2PkQqBFIqdDoQFiaJNDygB+9oEr3KF/piaC3NoOAOFxD5HkTXiJiXu8MWqseek8
yFtFRonizP1UKOAvLwCwEKbV6DfrTN5lCTJc7OeLVoPCIDOIDrBvvHFWSUPQBl07
qPRqsdh+BN7PVxsQDCmVw5K5fsvHvvHNgKeCqxgRgqcJuwd4TyQc1KEr09NhPL7h
yp2y3hCUcY1dFYKiKnXtRUGeVRcznp948PQjE7u1dqssizDhkB1IxeXxeOBR3cHg
6pQA23PHCRzTZwiQmVW9dfkDhxYP5Ee901sSV1EkEntAYBwnFp689f82p5EL3oEb
HVRYC7+JppEy+zuAB960/AbCpqAcTtpLAV1qJMgswoVVnxEXZfnLnmmlq2Zc7948
r5Nu1yEqbOQTd/Y4a4OyzJfephz6Z6LLlOX1BHXhe7BjKxAS/o9S0nROECp4AZ0d
MZkJP87WQcbTVVramiMgNvmdo9O0ksPp5++x6+bGXGCMV4ab4jOCx5RMOWhhMpv+
ce7IxqnKGbtTdMTy6UXP1fso07EfbJLg9qqAbKxnCqp1X1hpLTPGeBGeMVaTUttm
Jb7aXooekLJz+Zt+c4r2MoXzsfgayjNCQAN60qiHFPWHrbH5Ngw08YELfV/fC7Rg
5+3RWW4LXvuyDWP0YJdZki9GCW+YgvuE+IvPLe4nB6sqesawFYTyY0RAbLr5wXH5
xnOmNP5GeiZPyuNzWsAPHGncRzPTisFqe78w1WLjxqLnok6pkbmHb0WFXehBUVmS
EkM5YJk4PJXMcIemCo3RGpm2UELtCNqb15acS0pEGqzvIGSZXgQqw842CR+BLlpy
L+qNWonXlNxJKf3lqqIM66JWM0W1Wm/L+TKdqiOiKKLzM3SrVJr3FN4iqrIwd+11
xGZiXEJ88d20gCvB1w3fGe5aUvYFPzxHPf3kHrj64MXiYxQTu0xWk1hn0H2TscEs
YVgPAKuQG7zraRdsizYhw7/N7x2PffXk1kKt7WFaERUaI3ebSdJJNMTlClXTd6jQ
7JS35A2IfPXea8OqjIFD+dwwJpWp6g/FZQyRLU13ur1Ld4hW2zxAKFG3zMUF5BOU
eZjah4VCpUfrPViWIlSSF3CBUQ+UXofTkbUBU3Bi/AiXobrD7K1aqnc4zsp5QTht
lI5aswL5BjmLtUI59Z30GJMF1WVJ5q6EUggaAhnGQ9dVt5L0N7TsQnSiw+0GQpdh
RP6dfCoMuY37/MDYydYI9b0clNaKEdLyh1AhSqIa739ciXWyMNA8ihTlkmuJuCTZ
YU8K6uYz2YF2O/sHmPtgIQ96ZapDAG2ZefbXh2RM66Dv9mQzkD5CMReA6HbrysW5
ttUVqHTdG+EKjkAH5ynh8Q8dNmsfN1OVZhtjHKZvA+oqYtEoBFRdl+zfuog7TR3D
d6UIzEP6Q8n5hajANbWZZCH6GvXAh84UXNBLBlvpOBQr48JYXf3zbwmYiuW3H9Fy
66GQdN2NRhpMn2GTTN7ZRmJMnyzpUry85qyzP5YjQUdqug4MtGfeujsBSqXi0Wp8
RYjS/mbMoyB8P9OYCfYJ/LDMK7AJdTnbW99AnbdzOZyW9lWX/UhK0B+M6SQqC1Eq
luumQs0BHOM0G3Td93e0KsJF1FE57Fa369QLHo1oDGQ2p/AYCl7J15e4rXsp3v4Q
Tq574Z22wE9g7S/hnUQrolbyKp1l7/n9ot0jkJ6NFizI3V5dTdApO5IPKSFweyOQ
cyLO7ohq9z2Ec0Xf/brh15MIlnCyXDrSZi9qG2U0y6zIW/+yuloM/Dj0BdBq4AHr
vujZM+Zw2mIWgmt4tiA1gtDrrsDQ2BX40AFo5+xQqqBsAxlgR7M0JBckUYmEbVdC
dw29XLi4mgA/NKPlUq+6zwl1wrLipEXwoKK6nywfkVGaM6ar45BN2Wzp768PXIVb
A9wRFK7Wvx++a9vsaffeQQhpPoCG75T0RByhFQBlutkau/oWJTHBzQRa8OQFh+zr
SQEmNJhLP/jSLR0HrNYVwtOkZqahNikxs+l6ol3LNDoL0gu+01KLq6LuHskY8ctt
qJ4AwLEAixwFSYjnahLbBzbPBcyPstLNw69QQIH3nK4FXz/hZavkkiCiztzZei4P
LhwKShZqknDTERLEjEpkB4mias/Mdd9mGK2aMfQUvp1TvJOr1qClV9gCR9juRlWt
+6JLkK6+o/lPci894jtfJ0ipF6k1XkxUYA6DvQ45Mea4asDsNDh4rD/OOrpkCnIM
PFqYGy9BVrF3vVSG3j1H19036Q9SyRjAFFBshj4CGzDFEhIAxbZRqIZ/UTZU4F5o
KwEVp4aIWTCamVWIAKh7kVcMAavT6WvUwX3FqFsykjRLmu9HCWU0xzG85uB8O3mY
jWiMg0h/S391qca0fHv/lBvpvYUabhFmYd0qxd/BA7wOJ5X2WNPkDYongxlCmY2G
qRoPesw8M00EMzfJ3QN/jLqhADP16SHiwLGDFf1misIh24MsJ42QKhuJDibDZp8s
xvynrhSYsiq6Ou+ogVyO6nkyrHjzE56VFjwop6NbrVXPN2fTDDjzWF8TicUFH5E3
a70tL33h4XXACA0RcFAhCpXOuOpuNwnd8DUKyAHHA4DtOyf502G97kxJ9P3AWUVN
M5ypU1749Y8CJePrlphlKNC+b2VDEQK10FulFmmGlKwKP96FTqU3ZjlXNUV96Uik
8GxIiBgAQNv7x2T1/qriQt2WYO6TfGppjj/qIOhSZLtPR/1Sa1G/liHBIjsdpojK
sAOZCebLZFNoiqdQ18JaTdbWkjsqJAp1gXzSoym26/7rR4BewRv2kxy+SN5NpHQx
vRKSSvTlnUjkd36r0jbFkS4DHvEp5c/KSuZDVB0kFQIQL8Q9OvfHdcRLvpSgpGMg
CmvgD0I9FDSKO1NKiyxGUK3h9SVfJsHg5c14Ijad+WZw2A5W9nVm2wrBaIQU/ygR
mQfsbHbnR1tr1kFeyYyFQgLbwFT8rWMvxr4bnffgsrkW7wX61v7sV8AugtI0gvmt
aZ4qDLj0gnsdAUkO3XMib6KFhUWkH9udroCro6h+7S+jTCGawnFBixeVIg3f0SZu
BxzXMD7nm0Q6qIN3BbG+ArZZiJd/EtVLLtm8agm/iHpLItdUrbif7jkYlrdwCPNn
Jw1d8ILIPTOsQb/7n+pOtMDB/k/IMU+BBp0J99AUU2qjT28ASKlA7WD/RjvT5Vjn
BjTDL4Ssxm3R3lkdd3Uw3qIR81aCA3hEDRXWVRv/xenKpMc1lJqRabXnKbd+5hqn
oA1waaXa1+7GLwEuTWiStyyiXrtV/K0rrtckpYuSbM4a8teFF3a37+f4uz3qzlao
RiHDEnJ+mzSqNgqcBA3JnAzA7IweaF81FYeDIYpdnHrxn4PBzPK/OyW6anxfQp2k
2ODDYmOGmBSGdV5p5Lh5yMMyfmLYoVZLbVyMSU+fstz6qdQX3MPBE1nV1M3PMlSt
RDSMgJ+i68cLSWUxbw1VKGg9OYTZ2Sg4QxIf0uhBgLfCsyE9MDdEv2yfT8DzPf2T
LCJ1PaD2ya8IUzEV5621q6sW5qMiX9K4W0eG3HOxkRnEpZyuXHuMh3N+Z23CVbg3
jC/BCZH1iXg9Rrjlays4wUzH/Fp+DuVjxVhPOqkCUJ2OFkeIs78jt22V9gZWi1SK
BUpDG5Cq+0tkArdgTF3CyzbSIvS2DAOzzRzKzmoCys5y+OPCIERkMmY10ewP5pK+
Trznq/5mGHWkHk6nwhhirfszaHL5oZMLozR6jYObX9wcX/uor8YRsx7R3TyDUF6D
91HHl4x1NHJXzEme3ZhjMnXu9FGu2sN8z2pzENB3ijcV0MseofnAOC07mYuN1WOX
d13cuMCg653Q66Ft0WaiVK3NxZjEhsPWBUjUX8Juu/T0MDk/PdfLMIfUn6dZWW8e
CuCoFDorAAFVPrDIjxKCqGPreMOHkleM8s5H6m1Gu94sjtLZ8EWRhsw+MwfWKCoo
zLCGC1U1sPEM+8b3iygzfJdEA0tWOiDEi3oCP2l8byjptA+W2ekj3IoCC1TMAmkr
67auFq20wIsSzveMJq69ply05SQ+Lc4GXdJUcq7EuORoFgXilHQYT5XWw9UQi5/D
sel5XyQzcU42iNIPYp+oFqNHbL37ojp9RwaIZ7XT5ctCsA+4GO5hyD3ig3JWSQPh
1C4I17rVssixg+QrWXSxuDh+74/P/gREXhxDm+I967FI3UWNU3szaoBFanKoLyRH
f35V0OdxuvASOiPhqVAK14ODRSiGdUJmvlrOB1p76I/tJyOWCCeGsBr+6pWux768
hDuz5Q8CuPavghGgOCAFDk6pSk9kTvZ42AoEKNQ+HtxRRd1poEnEP4SP7YRE/ZV9
1RisnaHUR/qWAM9gYYhz2Drorjx4lYjpmUBDdpZTq7O3y6jg3+7uTl7UNXtfaIRA
1v9VPRLhJHyKELrmeLUCr+Ql5T/NaDyUcLCLWvCpC2EziI4+8LoJURyq+ItqpBlG
8HddtEdMTBvZeaQu3OBe3ZtTEpeROnYk5rTtEXu4DkFheG4y/XelGF03HNp7mKjF
zqkAR8bqfchYOYdAoyroTVU+kbnTZvnOJeJk9arZw7vpjgZGZusNKJfdVOxcbO8w
JGxJcPSuD+MlAsmpP5H+bHCq5EIpZkvpST4woRK2URy++BIVrKwRB9uP9EqXQL1F
uuJV9Pl16k8/ap0PZYMCAHQwliHP8X2ppSqy8sBdAJ+pcyymuf4vOJnpqOQiZagP
hHXpZkzz92kExmjXa/uSBvK0q6PoKHF1nPWTNjKufmWGwqz9AvgfWuXD3kiMWTwT
Pcero+NsimlhQDxhFgAyhXFgNM/zaqqWvDt5CUQjWNZx5GsWiAQzmaU6pw6OR3U9
O6XPISAH+2UK/HEBggPdAEcw1LZ7Gh/fLQJt1OeSB99ggf8yqvMflU5re3nfYDLK
nNl6j13B1z7Guo/YmbGKXOLN1+zbWuqDRTzX3Z7728TQ7N/2RPKTrPjw56xh1yiz
e+ShEpgCEdNAKpEo8vU+N0Fs5ipXNL74Ng+eZ92DssOn75I25BNmmeiR9nv6PaSS
6cjOZZ1jpTiv1VYglV5Qzm9EY6l6i8G6laPIrprWdOMBrwELxh1ssLXwVdCcxe2W
X9+rKPQI/HMpO6RR5M1egi3ktIUAaBx/uOcAs0Gm+PuKxwVUgSkmNM/10n3YtY/N
qBD++NRsz/yw0Buy6f3hRqeY9TAFVdTCxR/EbvXcuXgok332i6BVxfARkFKBPl6F
2n4pNlKugdScnwy9jsg7U1yOde/hyCVHFLuihX0JkdRvnHp4BhMDsvHUEbZNoIr+
AYD999Ar/lrEPpZjz+7HvRiybX9c1vDIX+JJi2k/G5XBhP3Y3rf3Me+RV3ySQ7Ga
zDxqzyB8FEmkG4Mj8fiNjOyB5SzxiZQNBnXmb1izwgECSK5tPBP3x9TcGy2BY/Yk
QE5iY8VDlNB+0QkYpid5ZB53gYsdJV7RWadKm28doYhDMqFVrjadmPtz7AR7Iecr
sE0djw1ggyD7yVNMgV/YRi7JaB2B7xyk+6TTccuHxULPtQLnD8IiXEo5ncbDM/OW
MwuZK94XdPV9ZnxbpLzXl1ElTjQ2WtnbPMbyW1bGFZ4+moXIMm4tP/GUfO8C/wQk
7RDNuttAiTatbF9MG9f7TojvkjTMcDVRjhw6k7rCgXtjBIYi77OxPsi03GF2DTPQ
NeY3J3lzqD4kUjRhnrJMo97k+l9uB36rbcQ+xfwxf/9B5hMnffw2t+qPfkLFGRVw
L3KnByPIIsfIQgIuJQdSMJEzS27ki7erzkZNqTfR3kkLWZWnFYTqZUdhle2vSCeb
AkaEU7mI3jDMKRoDbEsgJ7J6xPY1HsRSdODbaHLlX/ic8wXmq+gnbfgvQIUWwQzl
dIztdrQeNoLWIU4+U5SRrUPNzletkb4uKNTeRm1zkczLCgU8ynZp7/zJ9OISbA5l
MSHwOS/p5wkIqUpu5+8FJLyC8XGM5ZNX0fQ1hwftLmtxIVEI+ji/q2UVZgs+t5sb
rMaezuSJDga78jg0OpMjRvYqRLro+iQWWDi8HpttKUp6P07ZsG89YdqPZQ3afAaD
9c2VLmI3e78K68rLRurjwY/LqOSZmYesISAyFhBqpGwy7GBFyMd/JHKGzwCYZk7j
8mL1PdcD/L8C3CUgh8neW56ViutpjMWvg8jyuSVkb08QSLtjAovqcDgL+TklXFeg
3FykOCS0vi0w8YcIw0A65b/4Ui0sF2lX3U91WejEQ9Yf7tzIsrZVKICcPQwMNHeI
8Y9MZAF1eCv7UVD/qOpovMViitbHA4JK6Hk6hFrTeg2thcJzMnbSlyxsnjqC5ZXF
9QpLTKSeuTdFzfMDmZp1sMCPYprfW7vZlJiYOFP6JPs8hvsHnbb6QAedtkCDdrNm
Zb0yBPYk8VivXS0eA+30CAhsp64YDM6Yy/e+lYx9sb+5QoDoB5bZF91p8qRJ+rN9
CxlabcS+UnfpmbcjbMrPaVDdFpqdMSid+9V1pJNZYlKrcQaPNKmkC0KbIXCQFFil
mcWi6N4mKWveZOzzD4WEQgvP/aeU4S1kOR1bNA30AhXAkg4NUvvEEsJG/iu6o0v/
zpnvxPbF1C8ytggCLfuDQbN+dYlAnVHTNJWfXxFSouRoVvjcXrx3dbXwz6ZXQMsj
LzrLSABcXwsUPLurXu2VjIUxDN46T3Ued6rGhlafdrwyjeiMc7TTF+mbBzVmeaOD
5zWiT2H2/z1Rs8/PTegMD5rlcu2PviviFV94hvKqwfPC7ztD6AgeqGVWxlE3U7IF
aq+rs/0LIlM/a5LBe3vI4jtIB5MdC9L5XdUszA80IlNxV6jo5CuoKxYFL0jmwaGy
fAJH1ATazyjwbo6vouEoZ8Z/kwWjSNGl9aWzvJDjC08B1FniB1FJVb6xwgNaWHQA
YYtYbPR2RE0286MF3GY/Axm90Me0QoIJzO3R2aWp2HSKmWPMguf02aDAzj6YEpJD
q5WsUFA4JaNwhL1NW15kT+9vxHDHh0LOUsoRNGXXSoEBxpPeDvCV2pwNm0hDVadz
c0Q+tdJffG7GvDbEllVTEwfclVpHtOJg98+Q+Rp8APA83FQHaQ52V+TVRyj0KNiM
QH7J2rtFpVDIJccIACA3Tfe5Jx2Z6KfNkiq6VOHQumLy2FyozAWL1jebIoaohpUZ
uSDsKPN9XdBobP3ggdmUWJMBu/0B9/+SNdUfG5lmU1VqZ7s8wbXhjQRbm5bCg/Js
e7Mj6mTQ5XNX5koZFhtEfwFYdr13IxO2hLp7aQtvZROxfnQkgqazJn5UtNq2TqOo
Hm4vKlpQpmZo+IDN0kNrP/9qOTI1A1Dg6XDqFJAU288MEoMlkCU+W6tcWjxGTxWV
mydfumrkXZCY1x0HuOSki+Asi4NEpfTG/GNgZE4fRcuntaxPO9gzNLY2Jd5OHHZg
LPOLG9TZgm4DabSUMTJ0H3VUSx33mTmn8L1FzQR9lzR/UvZpkysWBnEr/5aRsOTj
vFBkz6Fr1tkQnD2WHq9rc62MvryJ+hA0C0r0vrgfBEeDKEzeA+fGA1Llsadof6O8
wMSOs1wt3EWuhL1pd8YNqn7wpKZ2VP1vArbT3MYAvgh4Yv52+pSKDTOku+PTx3EN
T1fJkmtkqlsIInh49B9FFfuNsX+nFlFHGmuhgoKdEN0/7Mc0V/dNKtZjn6I+wWSj
91Hy4LBvATldDzIs/7gcD04un7PhDj+DbelmUoAX/Ql2+BryAynScSwnD3mn3R2n
H5C6Hb5RN5Akn9nI9vTTIn8Sld/g5iwNAujqWMt+UXGZTy+7BDpommUhCSG3mXTg
Mk1WhXxaVQ6NOVlnpxfqOhvFc0jDmi8Pollp9BBpXvlC/yI+1Clq5sIrRpuSN7BZ
Q3oylbq6NTBg6Xz954TPmriqZfdOzrOqxrqKkkOeZP+plwmNu46E7BcbspKJP7KN
Q2qd0oiRgxGGGvscCf58i37oy1Vs1kXXSPkkT3McXIpKSFQBYXFK284UVIUK/UHL
G8JGXtvAmIArelfJhC5ucZMciNlbCT9GD0lHCjuNdDrHDjjjZWfS9QFdseggmLPI
FJOu/Hk2/5pgeY+bBBRfxBuyHeycxEWdRn6nda7YNjEQ5/araR9scza6R0/MVm3J
d3HXgz4O45XNeRx8ZBKt/WzXoxohLzQlkhtSXqHisx0LcxxvO15y5eIMdO59O+qM
N/XOX8Bh7DPBmYzuUkazILsijoe3TS86KlDwdCc16c1v4eJ2tz7UTJktDg9JxCEJ
Bnm3aITFW9+LC5KVdm+oJlM8pPCM5VL1jl3bihe6S7p4aZt1ZSD0Cy6DGYDNvg6R
INDPJv8S+GsKdpyT609Mfyy0wkVZoNPKm/XtYoX0fZrPeObGSJ1NrJEMzuC4mGrJ
DKQeG2+rorfhFG/J4Fq1qgCHm/cvCKmnJwYxNB4n833YMTjW/2yugWqrPZlcG5od
wfUjhecuPQu+NrDTQYkWZpWOXilvC+pJyLITi/pD74/T73JAoeq5QrwNbYOidk3L
BTcMoXo/ttfvC0wp8xX4Fx8cp24MkJ+YIf/jk7gymg/odO0vBisfCw76Yx+hfM0h
SCNpjyQ1sIyVd6mlk63G/jDmAercfjKihGeNhSrwke8omNj0MONPvLeqJ7tDGOlA
aiBI7mgdqsLXh/kHwNvAakqudYowKMXBoNdiJujSdZBh1cA7kUftI25F805fo3T8
idfVXWUl0sWD9AjiqAsEUb3J+dAfPV4yQYm68qbkvptpUtxHzBhJM3JzCa5nhANJ
05zn+t8LT9oFn/x7iGuOrXuxQswYSdYxMst94fizChuBURAv0BY9Mb6lpCHqKE7z
R8CGXglOn4ZoDa/wceXV2OSSJ2Pto7cTskgahD0GpKpRvUQuYn7JNXN2Ps58gV6t
f4fUx/25v0npyyQteTAugwnZQIdCLvJMKx3p+LV1WhAW335igDLSsUxdfPrCsN4G
Lq6InlKYE/7EIRxOjfULxZXOlWKvnITizU2feiZd/0X2KVB4q2cM5D+tP28sq6yZ
8Ly1rR3jBxPtNTOD4EoG8aG2dDxqw39LAvzbIRbB0sKp0ilWsHzAnWn4Whodqjy2
gsBypoWNcV4PjHqbFCTr8NHHBu97VSVvJFmtx7ofSZansWzN/DeIcrr8FCtjrv5m
sWwEQ62aq+oSW5xwgsx2lxGJ9zGQcHet/jT7NR7GWKbofEILnLz2r8EH18aasmlo
0dtYzUUHR4zEL/AkSav/hdBERnlaVhV4cysON7R//MdKMz8agGJFNoFk6L+gXeAJ
hTUud+8wuCzZqOkIKOcdeP3pDzdlcTfZYm9RLDJyaCFST/44ZlIEymHrrrl72XSr
vU5/Fozq9t/vd8Y4lB5/msqlTasNkz4Dbrg3jLN8kKS7CamofcK5gaUt34l2Gd5B
CJiSC24A9eq7iskF9qEjjBdngQBzFepWm09VfcMNR6dqgUiSvzMvuZhyOTCDzwKj
611o+g7XqDXc+CR9g3edyS/cJJt5OnZ8YyGo8qX+QKpBJJuyNJyVW2u02rg/o5gB
cFnR8vCaEOSAqOSrr8OOHLSU684IkldABWvIscWDQUeA3Q9ir6MA/xD8eNkPx+QZ
LoskyYZBsDVSYihCaVa7uaOfbBEaC0UIPh/xxY34u1tEKhlccQ+Giq/PWvTkKOXw
EeqN4ZISx/btAXiNv1LHkFHEmerhF44lauH7cZuHP8QRmz7wpr/PYcsGv1OysLkA
yOdmr+j0vD+8CViseKV9G4g4AswgV6nFdxVWLKEPrt+sDiloHdZWyMpolA6Pr0PZ
2EDN+L8NKmmDr/oNd8dpimNeX/0cMyvFXyAsE9BSFHPOrmEFrwiwPOVUEwBTN6w0
gp9U9XGaPbxcPmv2nWs0F5olb9yXK+vI0h+xATdNFOMn/1YH66XqJxzD6aJfx81z
JSKckIKh7lcRos/0PIe+3t/aTBjz/SNhSDx2AF9BTrbF9yhCFrT3szrLFdCx3PT/
0IKTBoIusm18VmDjRfhwvemPoXfsDonRUE/5OukdL5AmSRGo4CvsxEvuNC9KRcuO
s1MUclf428mdBgvAAZ8p6BwbhKPSIBBoHA5h0ofJgOKZya3J0fF0VpOSX0fKNWRB
c3VcOrbkXrPpLR3OwEqcEDxg8JFMjMUXBoI0eBSK6EgJwko1CyLVFqz4lc6Cu6OI
nT8MBg9JbnV+nYvwLI03ppG4yKgHj4eQKfejhmWO5zKjidfjvQ+53DALqndH2Bhm
/sPXJc6GVhIPIuctMKMIsV5g7tit52IAwdhslSHHSouVfJC04z1Pj8bBPh2T39Tv
32na+4UE7fiPH2mrUmVhtUO8Qq3bsRqYqu/jjKw7ns2BaRdVypy238PKaza9g5y6
Hx93zrEXJwETx/f3ppTh8JdbzPntueotGx1SR5zFEBjbidohBTL/jxJ36p6XxdJQ
A0Ke8m7rVVVRatp2/EoYGF5DMfMfWXDH4otOyhC+ptpSbyzkAG+sMNxdZECFcCaI
grwNh3GfE8IWFKAj/KOV0QE2D3bNkKDr5xJR2taAp0n9i7nUgegQ7PGH8jXUaZis
GtdBo68vFWI6F/180h6g+vnFz9bPYyhhSqjTA8f09236y8FY0JFb9b7eJzWm1g8h
cTNGQXjEPsdfRgA6DLgZLy+5FZAmlOVwdCltFOUzyu1FhFBBA0f4+nR0VoRhz/Td
ZEriMMXO6CJKbhtFwvdOHSB2uE/ww2NtnVx0HiuXwX5yTTWQkJI4Pldcdcld5jT2
Ix4Rn3avf50oOyeYwsabZAtpoLxJS858BWhJHmKOMRQB6p5ITY6RyjzAGS+JPtd/
8tpVwBpzWm0oQtWW+rOUWspaTtmAaviBL7z4b86UPZrt9Fra5iOq43AJCed8hKNG
MTi69PaKU8Fom18uxmwbWHLTSYMw0Q761Rvdrf2pl6VVJnBj2A72GZBVETNPOpP5
Lv3tlCcL7ml2KLB/REPH3wFIzCOowWyKmDrlFPhrFTKKj4jlCDBfcr+NhSM72Jdf
2v4LHSBU2LDSmLx3iM+2w4ST+RiQWG3ITHAxFnTkocdLkvHIYwQAo0FRpZyudIA2
W3/HhLbmiFzg1h3iT8C02G4/MK/leTYqnxV68MazQLpEOxRMpXc39IqaCQztq5fk
P1gIMBPiNKBT56LqV/rlD6Jg9W61GcHnKtvlWWwskJX/znSHdR6zSvDoaJAIfb+G
Gu2z7OPaZ8MZ+7KuwbaFCMvWx1gRy0CTSmAMMKFHJ1orjIg46CUQCs2Ewp3Qi/K/
oolQYTcPrhpBS0RPMDRK3Zqgp9wofb8xKF/ih6RiPzqVRDKQ877ABE0QwaprUoEl
2mtc3stRhf+MwBMraMWD/5jlfH9hmt+B9qTMiTzwEBwN3fLNGpIPWP7h9YutNMt5
N5AdhZGsRztMxKuLhSfHqnO6J+mLzU6KDgqFY+MBkXabd1ZFdBy5TDRY1yEzdadO
dNAXgpQDL5b8jx6zFTxWuF7TOvBckpwVvJ9gctf/C1fEwmb+h0MHKm6tmssOyNzk
ULv/iGGf5szY0Mo9cHNxolvx1qIaVGTogGO812BirKFPI6lA/ob8M851Ijd+0Dcq
RvQrQQHFruqUe7NpJC87s9ITckbifNiNsmc9CCNdCpkrjAFGWb/hD+1hs2SyvyXS
RHwHg+nadNEhq3MHYYNODR8ibhi0hb499XMadiXXQZav/yL1dlMdhpOv3uYO8r6I
ox+HA6KnjNYGokiaeCpZ6Wx5mxuVmhHqW+p+FxcuZ44DTLepo4YaM29sQiHbLnPf
fcOgMCenXM+Niewk4skRwIe1GfHd1osU+2qE7Nlo15jNieLxz3e7jCYHipagawx2
8fci4GTofdo9ooJu4XUovh6HKLLwblbvMpHuDq2lHh63C+T9ZOA436Djr8BfW9H1
DUy7rb+OSIvEX6hmI7SV6EuTbPz2oJRXGKU87XvJL0uk9AflhKngPZ+JIJ+trq5q
FWDWYgBuwFOUVhpqzT90R4n4VgxH+vS+L0d+FOCcxqefO/mPf4hIEd++HuytP7TI
emnZXiAApnOtKSA7/tdJf2Ce5h98QZfjscHoBtMPghEL9avms2xnQ9chRqBqRO/b
dBD+YEu/ZhW0fLH8FkJIevCeT3nQnBmDsiUYWUUb38IFc/ncACfzDPkXSckPLKLg
D2SHBpcD5KGNm5hMIOQFDBQTi2eO1m8G06WbMvNLMNC6s4/DJ6w+1ltU6wRiqR46
CODd0XO5Yd+yIiI/0l72/Oeib3CAHlGVgkEKwK+mArgL6NpgvSAebcIsTRHYDCa1
Azz7M7+/fZcnzwnPDX+pY+dPLsKLe/AWPiI0rQvdBR9U87d1HZe1wpDtEREy0Lyc
P+b+OBlugkovYfkQZR4HKA6Azsn1hyieWD1odkh2wqXl9x/sO5Mk30V0mefYqyke
yIZwfPmz35KuIQq/rztunQ0e7XYeWtqjs3fGb5c3rZDPclV+cRtRgAyrJF837pAa
vYRFSpGRtnhjdkpE7qtvTSwm0C6FOZNbV1zIGNWG5CUvE/kN2C0v99ZPuNfXz69S
JV83HDwEtHrF/GARUAzwcOtPw2GRCKsYaucuuUnROTetg6DeRREje3+lG6MC5rBy
J7wba/7f6qxY48+edWWFuYe6qZ4zYQ+VTMeEjl6KAgUaQ4nQlFYCjkrkjIGpda/d
Cc7heQpXf5CmaGanQ2wVDKHfASGv+9WH26GQaDbsYB6BvAurCcttztO/MqyOEsrj
2noq4Ot9t6o5jjH7SnU8eXxVapcwJ8ShbTxK0I0vGv2Sjo1Lib/T/1476BBX8kHg
ik5SozSegTFRtMHFANS97y5rEqMTLyvKdtvjHpAM2plV0NOoA+PBdhqedfbfMGy8
AMG4tsJJRtNKkulyeJYk7pHioB18A5yGuy+Y4wj6subPwHhZceZ957K2RUJ6mYTE
kk+431h0r0e2Fbks0KcbBiGUF8YtbcKUCDgS6RQ7+ewG8DAciGZH/fbC7GzHBQx4
OxGi+DXncWBFqgg13U6MeQO7t4WC0veE6YVmcvTxn0virtzI2m1y7g1i393slcwA
4rfhwr4bU+u01525l82Lp4yPFxOq+trL2I0lYgiT9q/mDl9Q1Cal09eQekRJ1Pvz
CSY21WHKQtYAuqM5GmtfQrDAQy0SB4Xry/1Mpi/th4mIkgSNOZnIKQAotRpCrkg2
4TN/AalR6ZLKAbROQWO7JFBcdDFTed/5EscK7dqQ3Hy9dZ1IaKr+vbwqF733KGYP
qopba3HPuIYEXFD1xusD0+azBK72U02nGSsX66CEa50oGhLPo+Jd+rBPxM6RjD8d
QXC4CxFRh4SLWWe7zsneY5axCdAsAl/jI8FAmepvYyHvs5OTSBNVOJSI1PN5YZ23
VYWWohX0uSWghi5XK4ry4o/SGrQtYtMKvbLi08jaWVeHnWYy8y40YxfjQhTAGcEY
z4ltoTT9mFc3MxUvlgAinpp3YUCYqpNvuTODyE7+I78+mdjTzfNmjxEnQGliQJhu
0sAhHUS/uOjURN+VVHoR8s4ekBn5JCRvlDzBp42R7dY12Kb5b9urSkuUh7rVCNE1
v959l5oAyDJ9MBKlc1zZgjoDIoEzed0JRNgkV/OOKR+/gTNCCr6JzTUVKiP3u4XT
ZOgAeYz8Qnpr466HMxTV08pHy5+yvNjGbrvp1vjfSr+WLXlKG8WjQNbyZWYtGVh0
54V3efraDIZWcOpTXrvpfiqXfSH2KkHA3SkFryx6h8BrT8DDE51ReVoKKvUVrwYR
S+Cr2nRTobQ/S1ZXeWs/pqbcKYoSrMv6pTaIo7PQwsb5KTjdq1i9S0cYb5s84FVX
TV0fpxixlh9m94hpJVfUOh5Mib6nKAQ9ezLYKuEr6aEdQfnh3W1gux7tgmtk2HBl
kl9nxVESPLDGJUhryp+e1WE0QLJqDw+mXml61bogulppum9xmTY1NKHrT5YW+Cf1
qaraoRlpthqKWgoPoRDZ/6dqGub6yo9NTjC9zGV/piA=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDchidqqHkmZDl/qSiOc4mU9VLEV8Lp0OZb+sPaqLIij2GYheeeQ96j4aPC6wzpb
TKo8SJj9hu4ka9ke6U1tOOj932Uw9Xp2ja3sDUseX4x6sIxElnI2gXc/wsm5Od/+
U/6O4gRbV7RBq+pvU9OzuY/umLuKWtdmqwtQ5QGESiFAisOsaZC+iGXR3k3reJTu
JQTEHZQIwjuU2ylvWDWK8otLLH4MxiSdrsnhJTq89Bwo5EaNVaQMPn1LSTCwU37c
UdzzO4DB3mvvd4aLrSYjjKqJnKMcOid0502ZOSNiAy0EzRWg+rLl1m8Y0EfxZdBA
t22/yEYI3dh7oZDeaj8FZ5BPe7hhwgaiQMP0sMNq6OS2YpAq4hpfDOo1XPr7IKNr
UFFRZYqfJyQqsZzoFzgnYuDIKuOyHOFVZR8jpSoWsckV1aUDCJXZkBv2UZvZ9JHu
L7dcfV+KkNhZLBdhC1mioIyG954niS/GkBpBv9RHuwwSH5rM/ILRsVn4fa5FpM4I
CLaJHE4p6o4vCCSymxB3Brdkn9hcFSPlLdszaWxlpyfU4itr5kOBVpNQxjvtJCrj
lhJ9wTyiP7uUGI6GHMMuiuVmcEGBwXTwTm/pN4DFiDsyvArYkpNfZDDT2LL5uH8f
8PzmznWVlmf++/eh5WgP5JMwAu20edNDnsHjRsHHwdCsbqSk0QWk8cp6v+qPbQ4c
KEaIZnNNDlYyt96Fle/Lp9mQFh0eE1Cyx2+xS7rnJJ8S6TZMKiZG0x+R2Ip6xfZV
V2fd/7S0UE9LfAu/6aRRMccpUCknrxHAydk8J8z1L+pLJb9dgeAmOEaLDgXr5ZtU
`protect END_PROTECTED

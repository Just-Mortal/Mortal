`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQ7AszDhlucrZKmnqav/UEz0srCB/LYP/TsaafkDgzT0z/z5fTs0TRug8B7y3Vpx
ObkCfG9vuQFpyKfOdDMFQFUOFGilPrm3gwkko4MAS2whmjs+qlMI65r4XKhNGdsQ
hyrfCAXQAzSK0jb7ubYj5qdnLsjJJUuaJAXI2uPh9j13NgYNQNasTfbiCTOSsaAP
XQYmDQUbgd5BmCt0C2hrNe9zT72ONwbzAOOmIKvnhfHHRAtWCpIsxGZhp0Nz2TG1
8Ea+FjHvYO9biu8H1jyBl6WngGNuokiqyKwABhevy4K3g+0207WsN8BVUX1wmgsw
HsJxQuZipmUPQRnqak8yxIdYr8B0CPIVrP4n/MPOk/hLdOcJSsGvf5Q6Qxkm0+xr
hrNL6YozUne6o7/QMH60mEKvMKqcHvULcKO4oMlI7BhcnX28vh9/NHSbSAUxxZ6j
gozckeXH8Hvv0jkLqWFuiEn4akyhLKr/B1CrNesdXNogDtTxW0EgUeTFkUjhrZL0
ZG7cg6nEhR8ZOj4nRw+i038JqXeZx5l6Z8gF9Tv65/o=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCF7VVn+x8gf+WWut3xMilwEF/xRj/1q4OiImFdR2qkDieRbKsXowKx7ntR6+EFv
9siH88KT656El9tbhORH/5mBXlbKV0gPahQhozUJijSSq9m+fvdULXGh28XoBeuM
pX5zatQ5w+NEwxy/U719KmI62Ro/sRwM48c5dnEYb0fQIoOAb+VTiO6KsPFh3VTj
YX1ILYwZwcLwr39emkEfS/7VFOc79TasS+LNB679+3mN7NoofzFh2P3G/hURNwe9
VVilT17N2CNtVC63HO4sqe+yU4dIn27XhvUG0d7GX98NfwIBcpRdCmDMlXms/QYY
3Ge9sMdkgMNuXVsC41Shs6J+gWV3rKybVycgkuZlQqCDfveLzMdK46HfkJUf6RZV
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PaFGDtTfy2tGUAD1VdOSL/o1L6QDBPYKUuyiaJ0n8iV8GuB1yGHyP4VXQrviSlwZ
ajt454LsHWkF26WXrGogROHmRaVFSpsXTdLUOzkoJul3xWvkvBUcqAtNuLowg3Jb
3Q48w9U/PsopFS4/brn4iIt+XC/Y3GAee46xzN5K4H7+jEavpkPqM79+4WdNnRpH
mdosLuM8YtQ1SCdYVJjwI8uc6ZhfFbTa93nIISFEYmQzN2LSMi4T92xFOm1vVFvz
lcmsgnuAVVFrgPbi0eaKayzjTr3xNdOPutn489YTw41MTGzMrG6o/k9ZKQp3yz8S
82RzWcoKk4aleGs6469cS8uRqheGgtVRO/KOo2oatlSgYiucLc23YPm8qwCWVC79
VLYPk0sd4SqD8EoqJDSHX5adoPz0lNzkuPhRw2fbE4H4CNfnLIQoMNvCFZalN/KO
rTonsw6sYjABuoQNgTBfdhpodnH0o+UQgn8xJ84LTPTMheFArDn1+asMufYkLKrn
2ii4KniWQUaT7hNFLUW1BYrSgUsGgBXkZWZlXVZnYfuWslypaf1l74D8KX3AG+A9
u/J+V/xar9QFvOLEfTdfkzutGrx2/N4pU4qJl7SSM6e4gUaWUCSlueCzyfsQrL4F
o67ENJs7J+OSNTtbEmsRmZDCVNo7aN3eFHc4nLHehNxDCaW1wwfp4A8xP60sQMAr
M7OH2JVB5erTHtRz2Bx21yC+4+EmH+GqN+iRvuXjBNTiAPVHd/9eUyeE+yA+iqMg
8qLpHRyC5ox6d47Y/vOSD3zkUnoUoLPoCef13NxTKe5Pmhnn9JfgAwDgTGGGd6CG
TX7leUSIg9SJlNEwzd0t4YKIS5rN9L+seiyVRkjimZRWnDJeuaDR25rrLL+FkFzz
aJJ2iVoCYNMiyQnFf6kxsnFgTKj6MIhd6Ai6hgw0T+3620ixXyrI9Be4H0ewe8xe
Z4tl77Nxwh2BCAf6fRHoNADiAZZsY0Ups0saA79mkPH1spK/HRv07aHG893W4A4Q
J63ac6hszB5ZvWZYf7VjaLUXb4OPazQu56wVlFU/0o8uRqfeu/tVNE8FkprS3FQK
3HqhFDAOr1dSJ+CqdBy2R0+Qh2fp12QEs+4f36xY216T6mOCertQakmfC0zirhJ7
Gr9K9wxBAAsP7lKG/skWdVmVN9MBMFd3HoUU5yFNw3uqbPTEhAL9meacHDFlVbdH
yfA40JqyiAI2iB9w1vdL+TuSPVe9t6B5mOwKIChViIZrKkb9I+2QS3mArio408lh
qXstSHbK/1QeyBdXdIMssGG9WLTOJPj9sXfWLG1NMGy6oOrYZ9c52TnHJ1taQxiv
R4XUYCF0Cw4b05SB4rh3tw4LHq+Mib+Ogd1M+9Kwo2Yxh5ykkmpbbHAOG2a+oAcX
cvqdxytX5DcVOVwCRqVSiv0r1HtCvOvvIE1zYtTfOoORucTc1WXINn6elpjUeQiP
4bfUE0T4wRQfF7QOnkgXhuXHEORH8PZfeTiNQ7CDnfX3T5GAAWwpmmt2r78bElwj
0K9BV4vi7xev9ag0WmvwudpYRe7i2fH0UmiraJrI1GsOdB58vS4UNE8EAhc+ladL
7HZ+y61Gdr3PZVJ8N+Lu2UOpJaJ4fk2ZKcDG4uXNVUIC2W422szX80olJ7A+Yb/O
Z7GgLCpBB+cwWSeP/DTri/W86C8Iy3vTQvLA1y+jFR+C2SqsIvjVAuqtvTKj7L8A
XHM6NX8KsWBQwDi3dZgErdiRfjs3UyqXTK1xBUfGETw8/yVNYcwr0FQU6HI4HMqx
teZQ5QelPq1s9ef7Eb+JAf4MjYIcCUltjmcJ57Imk64Oi7PQuiSAJLzItUbN7lKX
3H/O5tkdGD1GIjSKd88QIpa5OXcE+ZaM2udSaNO2cTY87hyrIeZM/+/YAmOya5N6
ydTY0kmR8reNz7aEsbEXgQ1vqrd9nwqFrYc9EfyC6OG0R0nkDIgIT8aMZUavIaEn
tHitVBVG0U43cxNCLVYU696KpDAKXfzY0GLgQ1FHuEOnqlasqAniNe+42G+0/nfE
XsUBglw4k5+/fMqhiEpdmXAPLCu2kAXFwxmOyqKuZneY6wdvSbjjqP2XsJkXMBAq
IJ1ttbu/pQJvFLOTGTVnwFwL2hsCYefDU3Z0w9Kugx+Z3NeV2gUqppQqcbY/TVTk
tgg3bpocSj0h740MdL/lOBa3tMuC/rR6+uc2vHK3YGMJIHzd1PAFAxXFijfUFGf1
ABfr4Pr+X1w7Opz710bpLXOLQykpdGvWsPEHHW5p0haUEioKIvIzp28BwcrDWlDN
Y68ufXAhnTXepk/OwtiTRAAUckNDaI8v0VbjWycngXJxXLAVcJKMaptjOC0AHRfi
+2BN5IBYHYv+1hiArGbaCNX+zoK7sjOno7va1XbUij7GecyJFchRaWjerdFQxEro
Q1lDzW8fUPylY8eWErUnzdENMVSmdYr2jffKbNsa16xOnb9EUVO3mOKjObeNUUvY
YkU+/JldAC8IB/Xoesigu8pf0tfVYAl3qMeYTxZhLr9o1GicA/nB6ERGeOQKkMmN
2UevzdF8elhEMmbES94JzO6JZqdVEwhdwsCjvDlAR4R3HFRAk9PeKGe3kXAp7h8D
v1W0BZ7Wxyru8+Te4qYNK4EgFOIBtPLvMduQjOBzGwJeFoIIdIl/3hKHsUzWdmNG
qZNN2ckEU1Bs0DDZqZDVOxmhdPSFCPosBZeaXTi5hP5xcoBNDeujrX6nihV+nd+S
TLplhwyaPMnseB2giqyX5gPeHUpCuc8NK1v3djyYa4vPcA6RJ+F1tlbkQZClxJO+
o068v2T9nmkSDUpKwJjRqVe7BLasiXdDzMDjRYcfFYY=
`protect END_PROTECTED

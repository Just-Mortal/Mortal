`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gJil1ZmQvzo5zUboSMN80W6kJTN1uVTNcJl5YRnZZ1SzAKftjUC6n3GAKa/maq9J
HGxblZwR02v5X3GdvLbf7v/R0L7E7M+q/aw+5vvsoZtWOFjBlfZiMfdD6BCBAW9q
jiNtMoSiFkaGjEA5JUhAD6sHkw17PVPjaOW8IM3JzPxI2ZkstqzTNQByc/EHpD0A
KFQT/bHK72IUgX1ZrQwiZLPR02Zvp0fwukFhKsZgk8UTG1xz817gl2SwpPZ/zlpJ
MJ4mvUXnR7/ppaVLWTVLh1C+9yZh1vaUv2hnPfR8SwnFheuNN2RdICAdBw+23bLJ
OZd5WhYFlc8iLLIAmiVndtZA+eR1Y49unkj99cKq6UfznzNFBzp+/kaYg6VjuoxG
MPiQhWaPvpS0X/vwEI9yOQ==
`protect END_PROTECTED

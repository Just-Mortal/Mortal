`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o7w+N8Sid15S+IEdZNtwlzHgSUVj+CEC5vXnrSQZcN9fR1JOsZFU4B7qNEN3QXGw
AFXUoUuasPR9Opd2TipjHuAvamNQN0SBdLsG5VnAHp4IAXR2reTpnsG8+54qUA1p
KXs/nE0BJs5xBwq2TZExemTE9UB0fzilXA5oSpIpsJUwPW/EmmMJ+EyOo0izua35
rutc9V2qXhYjFBOo3tyK1jrCRQ1blY88BAse+rsrPpnjm/sXPlvGaKbEWtbm/aee
pwXkXE12WGI5Sz+ecrU8/t5WAOM1F6e5vR0me5AbZIqDs8N0Avd5IiBJEhaPS02v
bY9/CTh0L3LrzRRH7tTHy8jSc06NQzri/eac9g3XBlypwVuVKIxPtsQl17bmjCzG
zKqIRgPejZhF2mQ5W+945MtP04LGXNseAvfFSVVPuw3buwZ0TnsUaH7Z+GpO+WyF
f584kmneYlZx6FqPBT3UYchj+LSmjJHb5BvnJQHNPe6vfDD1moTYgcGBjNmdzTtE
aJAVru/NyZhaPkpCfxj4rsziRBgzwwWkwfOEgjVCDs2Qhv81jKUodCV7KD2DKX2b
kpvMR71Nk3Hl0Oc27gW7u4UrTrRMC4H0AQcFxKPmztmlzjM7jdHOUQz5On5nH+EF
Z2YqgkpuYeeXEUBRHkHjpd8gfCX/YHkO4DifKDywjpc6ZhZBQE35B8GI4uP0YGq3
3+3++ZpvaeuK1CizkfUqg+JCBS3NT8rDzOOnAMDsc0Nlfz+QXPtkzrLsMdCM6Mg3
XTjkE/GkhZmyoUKXl2S/WoCnaYY9uoAJF8FFKbjwbkv620fw+S4Li+gsYd9jQVql
EAmyw+cIeRSCaJKEC7k2UC/pTs2oOmhtEyS9XZ9JCsV3MoElhlI5yuHZiSAsfgBu
ays9Q6VNGnQJ3RlTcReGt9QRcYU5h55zmx1aZtEIpHuCYDffo1+Fa5SYY29CP3ap
aznefnaSIVWpgm3kZgit+uWsm8FG1t7RM4uBetiQpSYTISAkoHpsE/ZgycQuJDvu
SgU2QeCoqyUhw+HPKhEr3eMvPfeOKsf5gXHKpze9MWLi6kpfuNJfcezgIxihcL0g
JZ8c2SY54kqHGnAiC7i73jONXkE1x1P67TaC2es5TIkpqu5Yt+ASMsQmkghPeL6Q
ymKOFD1KrkKYGsgOOf2fYyj/ZhWgxJFlCQcUQR++UlQxUMrV/G0Hs6/0S3Mm2l1r
dOK7KOtXIrcHeqNWK7T6F2z+yTaMT8C8o/w9ZhkZcqnGIIjHUtTPX2MYUyNrIvfx
0wksICsgg5xjmhehOG29eIxgJmjmsL8BvBOR7UttKP4o9eL/qjnG8TwvDVqE/rh7
51hFp8srpR1TsGbXsdBW+yD24mAA7LuS+kh9sDb335Gow7EUFjBbNdJ6eEiPPavF
/ehdZvBi3rt9szRoK7PrzXf08R+JxWRs511Dc/hmdxH9ytx45v748qvtb6VD6Gog
AkiRVZiy1FiHwQ1jLRbrU77lBktB3BKWjCuFFKo9CU5gLlIAOLZ1TVSq5V1PAaz6
By1NFXzEXBHXM7vsr9qOQMr2l8gyyjgWcEpH1FSMV35ytiuraIMOmvmmzq+Ju3M/
GkKAXtxgQJ5c9svxeu8yAVYMj/iIIPMUgeNY3q+MhnPQxYPe/tI4oP9yJFTKx2KK
w0kGi06w+y3K8jxpelUXr224HLNqTgqUeMpBn58IfEfTncKU5FeWgUt+zWpQyk7/
+g1GGKsDB4NHaMh2+KTZm1V+YIy4i2jp4WZxkXmogwZOU7iA6r3/GKjJ1fJdRtmz
0KFfgJvczNXA8X6uyZeCxnoIFpOORE06mB+iiiXIsutsECictk+bGjTS5Ssw9tED
Q5HK87qidZFEB+VRVBnl6LTV4lPs3EVF/GA4Dqa/mYFsFecQqcsydkGykEZKwyh8
A/5L6h1ZG+6dx5+Df9LL0O816krUN1c0ilHm63x+G1n4LkaDmMRWMHKKz0yQ4APn
guA8mycR3Z1xG+3lv8J9+yM88wZ1nVKiCOZV7paiRh+4PlsUh8UPPL0e5R5l7TZU
iPAnazjyBqjaX2OndMbU12AU0RaVx84SNaLXp6pbidJ/sNmXoml3LUE7t8yPeWRe
yP4uqL7lTu6v/+Rfzm5Qna2yezSqWPONPqgoYZ8KCGVMd5tRbfNpHegJLMwkqCyC
crYxHTem44kuPg2NagDhVo7O3Z7yo1dl89/JFDD69+oJGQGTdOuSLTpluCRQkYaQ
SHcbuWp/AvOBcDpgWLteIQggHNK9mP/YT9MT854kHBk=
`protect END_PROTECTED

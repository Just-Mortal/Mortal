`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsYPy9QGGYvfNEhlciHIoCz1bp5aPCaAJ+o6YHBSUkDfviWBA7CZ17wgSZpQgLRB
gn6yON4KGy0IJSXLyjvHFuKG1/bj8uU7FME1qa7i3ya8RGq8U+KI5uS0tD3R0eMf
51nWASNYeW0Hzt8xzZ0sxRoLMX0TTa7ZaGPzY1mmnRYR3Y4OBEBS1kt4oVgRdJxL
IIVODomwJKysX1NFdBN11Rxlu9pL24T/zgkDsJiZvrr7PnSEXEN83aIjGRME9LAI
6FE2vX6kOB4gxrftX9Wc0TH63RSqkv5l+nPMCkPBsxAzR9XDl3iB5VTrNgX46Q+0
e38bvPfVPukL+ufX0QmT4Vgh8xk/e40MGy+DvJ5Fh7I7sRmtzwGd4Z0es4b/u36m
SBlkLdBUCq8P0n8rCqc9XxKMUrymZtaq1VDiONbUYt647+ES6S1amACkdWzFLyYR
EN98CzYdn3HxUIB/KI+FxeXvLf/C6AHEXhAvF2Wb76xRz7Yec3JrMIQC/ENXxrM0
IatNwHcHUnrHbetsIcaU8eBdoAsU4d5LMxmEYd/tFuMwgaTpVggjO8hDrE+h/X2E
MKvkau77XybcmcdSScFaiSybEWB5ck7GKWsQZpk29OPsuSYNUXQljAxUwtFpar6G
swBdI0c6tSJ5u6Nr8GKQ/jmdk/XKpNCX1u40SaAtkdtulsggh6q3M6t22Jy/WbK/
BZtfyqP/8E5REmgLjZ1D45oAaTs79GrE1AezJU/kylqpQ6XglKXxcsZqfosTPGX7
uDFKh3xnuBLUvWBCD9vbyT8oLChooCAJCKlpndC0B/DFrDbQQQ7gdOEmv8KeJ6j2
XPGSE1jcAR7Md2ObJoIBgO9JET9Xh2XSD2EVbvIccM2UT+Z2+b3dzcqc9DNGcGzJ
AQfyzwzT7pQ+N1OwBXo19eHypkKFx4RumCxl+Em+DeZ6Yk1bgurGX6lQSAZ3bu/U
EGBzjffBy8by1pInAmET7U0yM+GFAUUKgixktTm5THu2umsKzpDfOx7F07TxMs1G
jYmm2eUVimS4/TM/+pHKRy46VCoAi41XDyE3ggiPv3bNJbQybqiJWgFHe0ntwDEr
CaMdoZCK4xZNDXpydnE5LEBAZolO5ghenVBInSCNKkfGuBirwFM0SkQuO3j5PN40
Uxq5ZPY6PLnP3J2KXAzh/MpX/c/FO/NkHTeTIefRBD3uQRWY+XKs10BBfJaYKH+m
HeljQkNVqCWZbUgKvHsXYVVK7oyWDVDzn/CM7SN27APk8c4GTdundeLYEyCfGp+x
52UcW7zrdRRWxhaXM6iRDdduKgLWwSSeUTEw6zj9zWanNBcMyADkonA6uHHAVqSj
6Uo6wOR/+CqLD31hxxOFaYoJ7OsULf6GpxkVYGdEbmYhNwvsx58hvs7em+RzDrGl
ZTr80FcNxm3eixqzwMu2rFKbfonLIcSdkpk6sX2H+RZb6o2VMYFTyvZm/FtAFUS4
pUJPbEeM7p5kuU9PoeOuXCoyuKMohQZcRqQRhdu/D8jxIM52fUL88o3m8L/2snh4
UEWrW4rwScxJjWb9th+iMn4j+1OysIGYZtkjtl3Hwj75jQJJb1r2VIV0Cd/mVh6W
AKOoR66qJ2lI2m5puTZFizpAlQLGnTH8YHQyEeYSK+Fe7CHv8IKClDtXLPUppT5x
djfywTPwLsXKvje8noQT0sg8BHRlKhBzl4ToxTL58ak6AVj2RilVfOVVABO3UgPt
y56Gcb/LckNUTEkeRiqrHs7mwWwfIt6/5+gMKxkb5VXli3VXx2uJ1DtaJ+zVJ70B
Chb9XDAG4w5I/8/Yx5TFoUBcVIrVSmk0lmiMq/VUYbE8kYobNW17hmJBVoZmhXaX
T1HtMtjV064vP2aFCgvG+wwo+nmEdkZL9ID1cdSWTGv1LdySDM08IdwWSgi1OuH9
XbzJBg0hmq0dBSsc2ddKnHYa7u9ye65ksk4tuROYktAgxAuj1Pt3CHJHIp5E6MSB
pjAfAlUMcWTPhfOOguU9Pj6bnmT6h7g4NZyKgUDKLUmEypN6mV3waTi6cl1i/p1T
oq2uztq0yYdurNpXzq6oLx/aR516iJDqaZlxWIZ1CKM+zc+3RDhGYC0sXkFsXjtU
GRYKLKg1eRoNMwEa6AmMWnySuaYC8zkLhfhHZShAfhDLr/Iy9t13Tjekz2665prA
jPXXf7bDAAGZkUkxGKD+3H0e/5grp9NxNKwFFm64jcaxSgT9KuLgV0fEHo7HCtY7
z8jVAPsEmgmVylCf0hU07WjlWWf1Wgg/1NI1+t0OulPMz4bLmRIiDxiTQSNiCPwb
NsiEAMT9e7zRSfpcnxvTRKOYDAq5yK1+nDc0hWG4xuBHT6/AEvocoEEvtIMxTF8D
HUeoBfYOy5rDUJQbFPm+t7D3IOXk+l7J7aIjCYjnD5SDzVy+17j7DjQraxWoCyut
L4TU3o6u3q4dAYMBRhafJjz/wdtWWuaY4o2YQ5iH1k+sl/Q/0HYvT6oWww/ofABK
z04EuTP/zu94An4UxoD6GCdGv5AefdsRbBDV/t50j5eSvyiBsS1QqHzEfmpjJkz1
arV6jX8APhxoQtcV+599lWXv9eWiw86+Q/oepR8gQ0thQKb3u861jxMkQ4CznOQN
c/az98WNFFjtv17ziwJ+rObFBY9zsZwycl4xnL9ZEt0rTK7iHIgLABaqk/g0AjGr
2eRbgucNrk1ktoz8zPh+Y8U62gQGdRqbsWlDjm228ziYmJFDyS2A+8odrTEJ45t0
RcjfDfq9ZllfciR/lnD+GFH7dsPpNJCA3XY3W+z/lVLl5A9j9LZv1Cev+fLP6eUy
YrIn4AnZZdoiHp7nygl4qMlo45tU67GeFTEJRouctNP98sOTC4CV1y/R3UrsRigI
M0WKDrlx9+0sLpHv9OQFkFpTX0LdXhIwo2EaTDwOMlw=
`protect END_PROTECTED

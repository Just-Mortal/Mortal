`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tmu68WlZHUkEkJ+Q+ctnjbqkG+UKCv/voGe9qpOKl9dJzMPDzcTEiJqfGtAiLYth
D2VItL9grHvLbV3eP3G8wjch+JHoz2Eiehxtb6vSTl9ja40rQgmvg/bMGXOF/iq5
Kg+exTQcmbUQCfXU2DXyr3txNeKKqebguGq09UxjQx5gK6j2vb1QHV5AlD+nBlY7
+nL1QXfoHBkDjQm1w3Q2La4HBg3SZutKHq0YaYG69JcRaGsZK51SLf1UJpbwGTJl
NedRC1AExp1kFXtDVSnxeiNLuQ2mN3dVTS2BBaXnUEkW/v130bVmlvMx6UBtmTBv
+7aD9azvObwjCA7H3nkDjeJfYJWgJ6wae8YFVj7qeHyVO3ENWQQzV+uhJ2QPHPao
STinJIOofiEWrbIEN+e1fUJMR/15QnGGXdMJF65lNIE6lGYw280xMEJXXCvj4iex
lp8YtQFqi+ATZKDly8re0gSFkJZ5S6Ib4dKE4l0n9yuPMmH6c8PEeAky8SLy8AN0
nf3lKxAJBuoR/t9uuF9q0tOSTwopbdEY0jDJYK3Jym+XqeXEILmTOs194tp0wJhx
hAB5FGvHCCjIJqiIWCpkbby8T6CtgBRj+jihKtIeYSVqRhBIXpDmujjV5NjzPDSo
W9TwkAxKHWJCI2zcRsrhDA0Yt0FatMBAxKAHBSQaa/CcIA2uOEbQRdri6kzOtqq9
X2hTVbNz9jah2O/QZPoFqoL7mNre0jMGXe/qrQw8KnHRbSDoL08d+i04esB3BBoU
dA6qQGmUnaOa1GUvW/jLvzQ8P4bWQYHpXLmvihRa7K7mkcCS21tYFHI9ww7570/8
itFhvPqE7HKXknNKyiLLfMBa+Kd6FJcnR/ROm1gQAe4TLWKOuoUxjKzSVsC9qekq
O57AfiAQOhr1iXK/Ci7t+KFXrPveBxpAfDVEDyCWDv1Zki1dMA6E30biMoAVRxs0
H2zOBikHTTlR6FRgz3+jlTMENAmFJxQAYwvilGiSf+8SgfX32LA/WW3/B9/ovB1I
oiCrKr9FCG7/FzOB1c3HyqE4keVIQOWz444sjtHmo0zD7xXrlNhBNyHLQpDZsBvI
oIgn3dXqom57x7SDyORJGl6tu7jWvWsetcmjvQGZP/iJ7hDM7w4NTKCRiPR4PMYd
1AhXmFubDvA7Lvg/Qh5Qaa8eKrWcA/uIf7bCPr6zZ2xydWGPGawU+RmCoham0Cp2
mgUR7Rsp0tKYxnuz9TscqFcLMu7+kJs2/8+ieVyRjsrlpmDgdqk2amyiKkjH4tYV
Tf1OaAWBndjU/fnZXrrWt2ymuke5WpldIe007foY+eYHMCLBdl4TEfQbE9tQXzHD
9xwJKcPMMeMX9R9mvNK2uIuyHBRn7pjsXaAUs1izSSAWrDnGeHOIdSMQDWdvs4sz
bMsSbhF1nBGBNYD4j19yvg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HAyr8+05YoFdl7THeklrJNhtpj9gR7NPorM5S8ah369/N+5wim0YoAJl+TVWrK4+
soLfL+FM9/MOlHbMdCkXljF/b10dDSKNCGR3ygjRnhX7tA+RWiUvyz1ERQ8DZDWf
91DJteRapzgxOzprxmU/wtr24CIPaPhvgSKdMmw5HBa7LTG1WmkKHaM0GFELWRGt
kh4mrtC68JUA0j8CWyTJ/3voZNUoy05KP/nS8/otILcSFz1QKtjWogyDIO3hQjkI
PxMbgPdUzUW/QPp1BaPS5ssht82do193q3z4mXpCSUWk//ux5JC+VHcKWkRWSVjK
pRmUAwbnZWmNHvH3eUXlerJVjSoSJMG8hmc0pL9m44uumzV/jP5VJd8f6e4tsuZA
MBbZ/wcIuUiVwWg80UVVpYRgKv7AFTvkUkzEKLKPoeH2Muw2DcowkI7/BZkJeuAa
qPcBFVv54FRvwq6rK1CI8THmrpjCCGB5aOA0rHhqOYhTnj5U7EwFveG4hlNaUpyk
eaIDgRW6jm0UlU1EticsTtUZbXlw5311eCZs3mRlhTQ4Sn8x99mZwlh6Mc6a//lr
jDRe91BMCKYgKfOuZ0laiQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1/bwI2Z+yANMVLNKj5trAqHO7Ivc+vR/YIgtcRt2L8So2j8yFb2Xw7yoE5H1fWS
VsPFFQxjR+fnonCB4H3kUm774nAdXLonoAScplWzVLTPDVfhDRE4ppXmr/mJFCs7
VB86N8nP5Itu/+C2blOMVtJ7eZMuYXsNgr9I1h2NHu6HFV41ePv44AD6b5GQLhvg
vmrJx77bu5gyastvPnxYJnZNBmMRX4dl75kRDTpzOxb5VGO0fEinZ/a4m7YCxLVP
A8CRM6sKSJ3ZR57Wd0/RY33yativTmzClv4Oya3IzS0JhoMXFmhgijoBZdxTavFv
2vX/DTFcg4b3hYeMsi6l+9AWjuExYdP3YQ4X5Ixh2/06+X5UXc4qmhk6+91n/IqR
o+YhdpJ7LSrD5yG7APui4a9JIZottIovU/Md/a05iOI3UvpL0AcvUz4HqoU3m5tz
nINfVaTzXBLxtiF4ur3OwDwHi3YWgm3TiejhRNvYOWh6mAy+gEq4VFHn7fPhwfre
HLIf9DSyyyIvDEV+JKSnvdfj/KzT+5rgOO3epUx4jsnF5k6ybNpwwRfgWIBqOswu
MmP3Sg1aQkeyNbBmLBvczBcb/M3opVbQC4Oxv3w9gbMpTPZHN4rovhZBOynLZkLm
pA74hV9lZYEhmYyrWEYv1ZuU+h/71DCc8LaQkTNQRC+d4m2goF00X6hpp+h8wVsO
h+OAqwKlX29ikR1zU/v6DtPIMjGwS+2Jv7aBC5wv7qO4PBPaWTFsuPchkAiPnLIE
eHTEMT8FOjyC2jPZo25pOQreR5V7C6c4sCpgz+qGw6/RchaWC/ks96HdqDWH+k5O
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DM+zstBV0sDMFvRy84wcDYaPgQ8OYTD3hBGFhPDD16b2wyQ7wh3nE6Bbd8T5Tg4
UtPg8KboBvVg0Tc+jRheL6mUHag8my1DDIUK9B8XLYPbmKy/bjD2zJhZR1EE/C4I
4kSmqEPP526p/bia1qvRPbPBPRBs0efut73fA88IPdi6HDI3P+XgFlw3f/ubAQQ3
uc3cXeJwKZ1tVMNtDjbDzeL3Y8UfNC99SgLi4pY8Aj4wDO40xIuvr01vs6om8DE6
f0RIX495Aj7qJ95ddVVLahJzGNeHz4Dx74W76iFnprsV1UpqCfqoRZHgSr5dtljy
VgSEJLZsaY8amzuJjCNG8gGEnIcQokMkehJ4ZnMyKc+lVCTOJtSSWoYChntT/c2B
bswmOk6HnekqH/0sRNiDOyIbRWJSPwl4pJYWcg83Du7lpGMUHHF1x2NoJogm/ivF
FT0cIsmajY9ypYf4kq8f8lnNW2TcFThW234S6hoLZ4ZFmKrZomUSsUB9CBMFvOHY
p33XS0251d75toKIZO6+kLpHPp53PH+wXqxTbpNcj701RB6IvH9jXHP0Of4fGBsh
jwoDkBmX99O7H3xYS0B7TsEVvO0pWKiV1LtzmyRBdFdJhEudyYpU4uGdrTwx8sym
cYAry+/dfV7PMarxLnV0dACQfikH73KdT9OEbWpEvnulq3GImFfeZ0pCqkXEw1wC
NMuwZ7tJeddJSneRaSvDaNrtgKndgcNLfJYDmQJYarJsjDMhlojx2FIGEj3+RcJE
tVRkPobjQZb8o0ETOmicCICf+rbXREGy1fzsbvPPR8qdWMS7oC0FpdY+YZUtirKk
Tn3kUeEzxUHOfr5q5btjAHetdE3NZRS5icwMrQK6j08a3W/TuwN0XWKxl6zzvtRa
00bMP0ZLAWrUP6lq7ucNcu3Kr8sR/AuLuMVm1ZXqTcQ38iO64dkujspNZzfS5sBJ
hEeJpW1i7Zp2COiqMRdQcUw6AExYIuc8DdbKtEoPZM46Zb51cMa7ysEogHihI3ht
LRIYqja0Jpby7VBzrIGwSuUdXnkm8JMOnWTqrO/tOKfbnGFDuzCQgucv7FlZc88S
5CKQzUgXHOCCVpuO2Kk8EQxX6qyd1bz64Rj8RKukNW86dn5dyGxQ62Q6u060ZKlQ
SSusEViK7iEycRxexrGWpkTV5+UFD+KKI5p4NT0zDZwlFjkRhePDeIJviOkLqaAN
FjIExietD/Y76SFL/0fH7jfGR1ZBy2SAP5GQop3YmgXzpWuxC5RBwiXN+pWPMQ72
WB1b3r/4KdGHrrie+NSTtv7+aDeiGDo5TKnQrlxsM7hVxPlZMAQuEEErlizTnOhf
MhuuGgT9Rqdm2JqbI5P2O3OonpXXBSApfkynSkkAH77zDqgZwFLc56WuuzvoSg7Z
WZHxr+59mONu8JRFRRqdwYEoYiHbBZ3G5/xSF5koyJZqyv0WTreo92N+NRMJKZlK
pRirUHhNbm44dpEv67NsYmAyu/aXoGVnIQw7kUMdt776Tl11NZgVg+7KIvytwQNr
UbiD+aTOYapxE4GF/0BJA32E0XIiyCOJTzfEO7VoIZ9BQAFDy92CYj9s1TDyTmRZ
20uZgrMZdPKHgjzwVud1yIliIdd5w+MKuvJ03ww4+LVcTaI0VKR42zXOigD32cL+
Ku4fPIoaE98Op6Ei12oeat2Ecl+RhFD1tXl30Yt3AKuB01eLDq6ClpJkj2yVXw2T
HHGayUODrw74PcVqgXCY/uqK6vYo8wraARtk7z3IgdCkEe+gTnsGxUldR1Jo0NGT
OML1vjaI2waSZpVcj3g4nobpovGLjqNtTnB4G9P4G2t43W3pZuLl1bBnkATGHAbg
m+2aytzpT9y1wo+VI86aV5SyRsJi7PyZXIW4Ru1LjSevveSH2I/j7rzfhloklfWG
EwJyZ58ct8lIVmBexnbWFA0d6NXRAU7K0jp2domN+sNw7iUgL1thOImOLjPgkNvL
8yTq98KICe8VvthHMeGbHTBmVO9CFBjqUbKX1uWq77BQzRe6Ev6pGAD0q8EQ2gWL
+jLGzbFD17wnnXaUn1OY4bYJyopwkxM4/u7coMhcgXHa6LUDz/JfkDW8c98769Ld
IoHg4lyOagOzZ1n6Fc5xkoYehB5KM2YOy/CU1xkMgrPhRCyTePLPLLDOADSwa9y+
/BeMIZoYiPIX5tT7iTwQKeRiXvLNDeRXrnfv229MzAkfePwtV/CwJrl6xiTR0TzA
cUKIBSmoTsNnApFS2gBXd45nHtMaXr9fCJ3lkhTDyr1TtIJhXTv+rIsmpJes4nTm
mXzQrOrNqpg/PQXH/E9JYiz2FUn320n5ZxI63YASYzyC7goFLp1Pc5Nz+Z84jnse
IlBe1uQTf80NZuZJmIYGnl6BhK0QMlhENj+jlvXCsqh0O+ccKaYe5qMrLOpKFaf/
Jg4HJMgN9PjzpvejRbpeJ2TWSflffq7dE/lsigurxNZ9LDND+98ZNAQr0nZgxJCC
Na8S33m7T+8FWLSL5aObP9CeTgPFD5Mg8wnWeF+mFZrJeJBz884hU5hxZSwos5Ir
yJjD5zouny/jgmDXBnd01B/X8JcmgZF1I98wI8tOqXPEbJKLd6IkywaYj+BO8OL5
2nXM/QzTuBiGJY2bGB1X2qckQlCnvMo6D3YHDTKwauyxnKpDdMZHWkvTuxf8R3Y1
cOow9eWkZSebmpzR8p8voiMe1Uc0qAdp/w0U6KVK3kdK1inURJFWYdlV3lGqLsXG
tKatX5vB3kE99pApXWB5H4HT2RnhWJzK14ZBYxCb/rrlNvLX1ltlRK3VmfwufamD
NTn0c+3vYzHGLdJvpFDhJwRI9/4M24PUNm8kfDIjB4LjnG40VbMnJm1XrVDjqV5x
hsb+29Mo5Lq+AhvYFfRpIq38OZj9Gj+yg2xqCaPBxW+rryEC7Knh0xbF771WOiE7
rjWMNgjiHPDFa/ARZ9rEaJwFfj9zo+A4zhN75Jkyg2qGzD/u5uaXd2E3nCKrlnaE
OheP/ROH3oMC6y7YResawqyWDV65cQ/+Yz1daxxHVhTSUyaZ8LWqNS6f382btl5t
7vkFKO7mq7SOzX4775xbtv74+KR2BhAruh2ynNWFk7wQpVtN6eQtmhosX4lxoBLX
9ZZIhuhB62E0obiT1qzE5/wPyDoFVkf8riKASDTXEOvRU7pChWK5MOEc3mRNWleS
Ti7Lm11Mbdt682OQ4vXMGXj2HVls+WDVfQ0NqFNVgpGn7zAreozsHd0+OK2L1iRZ
MmNC96FKsF3xiXdpgsFHroIsjDROTlsoEeY98AXqweKOvdxks0rEXJCiFFmae0D7
PSj7Ky5NFuJ7JuqNHAIDXi53TEbMbJ7+B99CZ8jl6S6UFP8HLunnYEtEzljmm/q6
x/tA9zhA/Vp9+a6WdP9z4r8EJ7e7+OYcAQQnm2ymEmxLOoTzGgDhvspHGJm8xkgx
rA1CuFrYp/jRmBQN4VKvn+isvDn8XRpEhlj9zhj6FgOwx1ZlR5rWtmNt2ke3oY1D
7v72t1oyLU+xWbLRK2ZXOm4qUZDCbZX/luSbCTj1KXWk8AeN+dAtwimmSLfiqSEv
qLFpPpapZMy8P9y08EdmRFlup6dvwjj6NQZ3EyQHf3ohJbkqPoI+6U1MEjLdbvQG
ZktbcTt9xCE2Jfib+eKK8G9mfSWAcNwkS0h1pK/CfvpN5uRaq9PD/J8MXjmYiZoV
LhVe3eH8ZK1nDfTH4YBpkTqiIC+Xo8pUU+d7zCkKx5vgaVvaD3sBb2Oi9yzYqXJu
38fz+BhBtxHdvak/LBRqGlra6oe7wsbsRofu+hsMgseZNAViLeSeXU/8iN5Lulcm
aNUXS2wY+sst455cOxFd0jLrpjHZ/Kc7vwng0j2DvbBIw1bl+qEqp7ps0fkyev5B
NuB3W072aM2c2j6hdt97hNkHO3i6w4mxtR5wH1/9xAuIeOd7zCILM+sY3K2uY8p9
T/ktxyAdUpDZkSK2DOpzTxS7/sIK+zM/UvGFFeznwNBMD47zYd5s26CBfMMFnu/U
RZWTgCxU3MT1NzQ3fPG1YmXZmLrD33Yo8HmoJ/IEwlE=
`protect END_PROTECTED

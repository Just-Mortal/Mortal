`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/p9jhjq42JFAOAt5ur04GApGSBtcWHTz4YuFDUdPEd2IvK8Tn+QuCE0dgnptMlVH
8ugFwzz+TZpbk6yS6W9hL70/N/ArSgoPTMIs6A/FADZyrUY8OmyyjlhXqUERRJE1
xSUzOC6WPQNTSpYgf/mJGDrW0SZWmhcjUL45hK3lxVC372/HMCB1EL/Gw3QBW1en
NHxgNdB+LWHKzyc7SP8lcXSJpUMfZYJ/1G6N7yImwIElwRS6G0XInEsmja+ew/6B
Z7ozas7UROfogU9CCTOe7jVrxtFsYtN/AC3uSglnX+L2/GSf0jbEWWGsAD2f7ayq
q858s+ExPyJzrPnEQBefn1dG/A5r2hhPJqSOX8DbNvXn9UogiYgd4pVfAWR8TVxC
5h7lg3yPFWhDT3wT3SDbeGZBfMMKSrPt4gahTvhOXffnJuTFWmbkBxuQFVhNgEWY
xfSEGZvZHWj1wZlTQsQB05xZ+q4SzGefLUpM4Bw6sXb/FqDL8yKckDmBDcQBtPgl
+bZ7wdaBiuzDxWUeYjeo20py+QaP/l8u6J/6ZxqP/WECBg/eSNMSZhO8MoQi6Wbb
/8bswjqW4PqLyHq9KbbDmGpmWakahzSQ4xcaiowTlG4vlhojcTBSZm+qzlwR8kc+
HHN+fEH37S7RCOn5uHGy6CQvBN7zEflA8CeAmU/CF+SYoNmbnslicrb+qa0jEDen
Z7EalBj0htHYxylxopXocSLvkEKB69rR5dEsJqr80VSm4Gr7NodP5aMVROUFy/4h
nZcRve89QEwfgV73UAvH/HtUlQ0CLrcCREmwI7otqgpSg8C9As+A7MvjUKaG+mcy
vOerS2aQKXfH3Qkr+uSP6Ft3ErJ9U4MkFJovQLGnr9nqmb5fp4XEM4tv2nISTwqO
LigaI4WLYRTZ/UOekkPKPL2Eic088w8gu8ZLPfuX/fhgCWPaTgLfTJSV+CiIKPIQ
Tzu0Sjv5bFk9cBGzIEjS2DdorwOz4TqYqVxL1zxO4PBN4ziuSYHKZWdZXHpr8Xzj
sKMUlL8GemfMat6pHMnTRrFJNK94scE0APoR2rre1mhh7RuYpT/jVk9hsUhQ1MbN
AbOvuvT/UOLclO2M6fVSQOlAgsL834QVfJCXf9W9sj7q8hScg9akKsJgNhlRSS+t
s0fuyYXB2iOG4K5r+PE1KcwkWzXuKB+C/vMyJn/61AxtszZJd04jgMhCZlfdnFyH
Hngr5nHqZioDiN9EDNkq44mFaiFx7kzYRUzNZqkRbhOtMkPGWh6RXleJvGzwHKxF
cQJbJgdytQ/gg0pTtht4+ByBU7WWOznH/FCQummn+e8zUuim0239C3EP1PEKc6G+
w6RrSHdjsvBh8F+C4OV+kHit0pptksAEd8iP5pA9eJwdzm/hDZQ3a5d6cBjjbKJc
eK1w3c/TGH9RqoyMJw5FrPcnnXmgFhE5U347QR7KQzuwzaNFLzTq8SPiyywRY3L1
DFFmBYSvToLvOnbeRlqk8gZU4u7fRzpAQg4LfFupYivPbXVC58dPZDnJnqe97LlG
RzuxLpx+lIVThCwQ7I/Ty7fm4/q7RMfHZWXEqEnR2ZW58L/6narCRQWJHo4yoOHU
K0K90Q4zBkjGpgEP6MyDmbZzf9/DvZWL2siH7aUORmdKsj3vxsnnP30m0SpIIGdz
EMRt3Niyp1ogj3WYTQ+nAMrjvGyi7KTR3i8gSSE1I9KdqWfeZRI1ZKQDlnk2pYh8
Rh7ZE25rFDfwxQgon1mNLcoPPDJ2/2ixzaNDvfFE9uEwIbLcXIXLvn6nOqx0HHaE
vbSGPtIA/fhRJKMZj7dHDcbVbL6ddsGMNFmpjPS8WuSyjCOYcemDU+NBjepLJ+0C
zhyqEtIsls4FYf0mcWVAcKOVsBHwXga9mTdFdMVUUKeQTwEbReMQ7s4ysmlE2Hh5
ZF0F64bkt4ItmooaEvfTp3sXG4uiAfPjYHbLYx7N0kIPeMUBXel4gnXSWuQEoLLg
dFX455EyOi9thY5cB9MPlvSdmvCs249BU2HyM4soAC5mnpqlvai5T6Rb9duT/cGR
WowMQwF0HwCzYvJdxtt+KYVU1RLF0GtH170IAN/Cg0gddYobpULoxbcGckFK1qid
XzLYQV34eOfO5MwbL+h65Gjhq0Qai1kYHy5LaRkky22EPBVqWQd+D1TdaeWpIZSF
kNLSrAbSWfywPQuZmgc9GxyYLk6KhDQbPGHGQK4/p9hDouOX+oAACTavOcMFjUtf
XvdHyLiyVaD3UsApC60B364ZaHCJoZzBYCdg8fWjCPo329hgUjgk2mtFYPzqBSQu
V25YNtlWYBwLtDdCmMXGGRGcmc+IKP+D5AVVNSpPXrN662ygQg7QqGEWr5HFfduq
7fOf6sbGpbCxlixpkLlY0PZw63Y9hkOF92S45ivg9rJXmefzjaj2Jeamc+tCxy98
XSVxK1Z4gzQOFFCEdcFUl80MoMLbKmtuaXHlnkpt5u2VRK+tpFvzFsBhjytH4Dmo
FZ7YGFVIdHb9Ofll7Bw/0cKp9Qb4d3R/5rE0AAthKUu0BgK5tr+wAUbPNd0SqkZy
asomzuNmwR0+WQB0Xznd7TldGZ2/tSnfCeqSFUzO4BrVvFLUphKBmP4pD/2CQOcf
nvx/D8Ln8uYMEujNgU45PipYWKWiYHoA/oXBwFRUI8WZ2yK/UNle7Xl15FSl1Nrk
iJHRfeKYepkmN4rvTHL3Ychwevo5YXL2+35SI4PHRBIL7adbTHzOeWifwaLuUOvX
zqgEzefHp8c0n09m1BmQX3Dr+Dt4YB3TmC41F/g4gEDmiQ69C+AzpMLKnC9nrr8a
wgvhN6j9Uqdkuz51sdK323EWO8vxsQpQTSuuuPPUZMeSxIkuV6Buuni863JMjBAN
zcCT12zKgkiC6fzUjhYMty6TJupdkeq8d739sQtWIAQJ1tEFwXvskr4ImDz8j4P0
YuFTiY+TvbpxWjJz4K5ZdhnZv4MB6DXjyOBS2LWS0r/fYIlCszi6pF4iuMCMCmpb
f7DUA9GfybTwXZjVDemkPKG9LnrKAMvbNGu4H30FzLYDg4mMVnttrzSb8jHV05cK
cVIvOgPDeMgTQxNn+HrpnKyV94JQNU3+USsm9uSV8q/SxWuhx0fwcCRBF/YMr043
l9TFl7mmgqq8+QZob5xdXPy/efCVhB0MmSaQNf0Hum1rf5jSUfUUdCQ1pc2q4yrI
84DAa5N356pp9OWYNy3BFyb7GGEnz+d4Qv8H3CjvWWSurRbESncu3F5vTurLUl17
IO51PE2u0tNuO1qUbSysVqK22rfac1wPH7KPUMJAJPyS6Qm2tXHWsOefaK6xwYDB
GTOdD1mQNSi28LD0oT8rV4DUZAQtbUrjVxosLtaTSuMLdAXWng+iLJCcIQBrIiN2
+3ixtvnArtVjp8YXhs5EchVU1hZQJfZNjbdn6TOIr6M6Znh+EAQb/+X/nouAQQiZ
p+QgZcWut/BOz6TBFC+fZj4uXehT0DZi0jimhAgg/Z6aGFD8Zmhh79XP0LIGAJBr
9vCYze19TdssG9a55+zHvqPIErx0Dp3P5bIdYwWLxFKd4Hb+4G4joXbv+wjCeFlu
ZaL1+RXBY2hXJ+8tTsFCOy7jYgtO50DyrpD2l9/mGcgdGeBa9yZT2vNQQdsfTGJO
BGns/DIHTtmMV9VN0DDippwx86l9I8ZiGDFdd5+k8n+OGHxX5+mSaFNk9cRDJFGu
vd8k8Aoz4jIxdu0hxuSjsWptaqaDH/tUjOY0QKdTLs+57UevAN9zztt4nBFKClio
wVJ3tbrswVGVD79bR3/cc1n2gq6RADX6YSjv7kBRUqC/MnsxaBb9l5SFtvF01hOJ
J88rL5DAJ5rSJ/GaZj2tIiFE7TXGNgw87aL1bB6yVySE4wptCuNJ7QGBqCRdoEUs
Hw6sqBDRosnL51OoacKYJrLNiPaIB4vdlpeY+zij1UqSi7QOlWDCbzCifDmicnjF
QUb9RCBNKpUQxiikoM+YurAX5Zq4JaMOlGTGr8AEBWdx/Y6NrDB5vK7vto+xs550
NJ9w7I9utyi0rJiF8doZZx8Yr2w0h+xlRJwq9/xrDqXdBFP+qtO0ysQDeQG/k9FK
+wNJSopo8+H0inX+LyaIyr869abtfl5yU0FBlbcfp9j5Eerf9OVBKi9pUFDeQ7Lq
K0qnCWG3yp00/SzluJQwAPIYpA2HjxMm1OayYH+H6G0LsRlqMg0vBfA2UhrfYpHD
Zq1sLEufgR/sxMjaqpVNeIkPyurao41+KOX9BCrxIlxabcjlSviRdLCysx2ezguo
77rtiMImjA/6s4l6GDxE6iMgicZEIu1drz8dM+LFtyn6oYq2vWhL2iZjR1xuhx28
9mTqADkGEew1QuOuvfcOmdNTyyZtYPYV4rwkK4ZlPs7rKzEHgC+zXCjKRVoc1XF0
9H+ou5lXbrTArE6OFz49EyLQnkT4LQ9i2HryAeeECi4+4jzQMCgma7MPaF5B0bhT
bGn2vbNXXSbnMUUECue+5a0MhC0HFpBI96A9TMqBM/F9kXZFnR5jb4kqTXtQRn9T
GRRdAISNLyU9xNoV4Jtik63Jb08FZU+I0DP8pVmwojELV0dMlDAd4UeE6WIfTI2/
gfeZxsPv8+sEVKwomP3HAVrxoBvOhX8XFgs/izq+wnB4wmTtErd4ed1+azCvxMn2
Hm9Hx5gk+qoUCRAWsDM54wuXZzr7F42AhT7BSIYoxSCf+bKleKp6IxrQ70d7Ogcu
49F2+2rLMYcGHw02okjSScEVXrd75kBrZGNHKvfQKIxOlLq7vsRJPumXi14edlOQ
k08jIBl/xmv/97I/gFe7Wkda8mMxG8wTVpuTQv1QL7cR/MhI8Zdy37apIS6RLdTO
DuvYKEkR57vx+VQ1J2qph0bXLuoDJ1cuzMG/1cpwZRVZUWuic2jK2ohmFaWICgV7
ryGRdD7V7vHN+NsYIm8C8te5M6zlmBzqlW+3QYQ5sfwKnUQtjhL/v/UVsmwY/fWT
NlXrsf3AAWnTmkvd9PM5FlWfmE+MOOAJ3zkE4fMouklpxsu9FreDCFPSz6XfsF91
py0WLWnKtMbg7lynC/ktsJ+QJosMhnrqmSMdxPg9TykzusD0GVAyMpIaB4bFDzVd
kKkYUswXG0LV8DeYvRU7UgjBSjopVDhYdDFEU36FawH8ULLVYtR3uKSYGcaZzQxe
QRCo321j5xXIT2oiSQ96R235RJNNobcPD8sffFJ+xmDJcA41X072wKPVfOjNZMKY
8iZU6B+6uGmsrdXHUyz0T+eg44WTegA7JOQ/8Hg8HBNbS52vNrtHeEKl7sG+Ckna
2bazcTlEuUNIe3Yjizwig7wvMn2aUVs3t+9ddrplN+PYhKGg2TrIpwgTTwy0GWf1
EiPVQs8QmR5VR/g5EAWuRs8Cgy/39CdCfwETx4I2KXMWysSp3yuOVK2aNg0XH9jK
y8hijVISY1qBuOm7eHjbbag9FeDDjYfsNdmqckzsfYuAN+I2qCqWMNeiAKjmxSAX
JksKjMjQPzZejDRBsVERH7kYpR66dL4tIqtcYMaQpMALePWJknPs9T0Z0kfjWO+8
9vcA03GG91cxlooEI9N0NJbk957DYq4IuiPJ8bJ3Ct+YyXeRCLGCtch0aI8TFu0z
PJltC7HaeJ/c4rZ2aAG2lAML+Sg0FXh/OEgzYHT2VuU1ITxcOSZCKsdzccWXWNGH
P3F0NQo1SIL+vwDGVBhVVZYqOlExiumCv56tl+eydqUhORS0/TDm/pt2OIFKCRhH
WcHjx+GujfEHfzB8OsYQLp11CCB7XvH2fhSnpF6gP4MzeV/1dbn6JFmWUHIsZRFE
XYSbIX/ogeNhLM1IIGDfAhnNWpQnpRM6H3714Bj95TDjHTx+DZzZOXmdi4INZ3OY
LXSn1lzqbV+OTuws0msCGtfYmcfdYYsJ2KgZ7OL4mGp8nOlp+rUf3nMNHJefMX1B
pIzsc4spMvWtZGWCS8zgCxUtkTCnrtT4IB/kKMmVfHx1ctryXSGazXC27SLcflDV
R3DlcERxARcz9zc9Si4o1y57pQ806SZVxATl2lrAojrfJIUb3WwuheSd/gUZC3sk
HM7z+o3AkIin0GlsR5zIOi6Nu0bFcGE13dCi7/rywA4Bkb0BjsLV3QPBTdMxsw/i
5oito0UaX8nH7p6UsHMBTcXUWinphCgemQosIvjRQZd6v0q99NGmhrkyIDRLbZxi
r1tS7R2xWZxufov/8eyMWhykv08Rth4qN+qDO4op2wD/aLPpOUfK7VpA8XTwv2K2
rfTaPINlRFyO0TVre/1e5Y+/XwGcMmNdAoH13b2YyZGrn+NlWXI1IUlxWmL11H36
980MglaEq2IVcSRPhnCIMZDC6tCOxAuTa9jU8y0w2DEYMQlvrbmADkDZ3xC6rD9k
MnPZUeCGj2w5puwz8iB3EiZlyZfcxUTat4mjG9gnXDYbEGeYrqPmcfK2oOwFIPn8
d7KT6nFHnilLS0HOq50bBD5+Lfw90g0kL1ZnTjb2wgU3pdaLJZ+qQ7aQVKsfFnoR
x/mQMeXMSOTI1wY+RU7RdLUwLwgE/4Am9yY9b5ROZmtM0m70i8WCToBxNsrjVXID
FNZVJwsFPPjydkwuzk4I1u4GSrsc8SmkExGGlAKLxLOAvDVHZ1Stw3tgxgOp/nLp
18i66baKjw5NHcfXVAhlmI5361PbNmyZL1AafNiXzwiw42SZjTxsICzveQyaHi3H
GEZMDtyDPnJVJN5sqoEWsYfvhXdVhGViBwIdwnjrSaS1tZwnZaWpdeu+oAPUMKgn
2jUVwA0T+3TiHXNBpmfW3oWmSJUITp4Yym0FZmnerp3/0266Jd7u6PB6rB7sL244
qq38gO0WG9XHu9xPV5SC72s4Qj0QAj4UWU7JwiUPqx2aShnZ6ox5Qwb7zfZPhkfv
G/pIoWyj/BHlegvxNJK5v5yLKBy8+fdstnfU8YFd9OuKIBChzs3b6+MjJVQBNezU
n72smJhKMgVzhRAYl2S7IFELM5aQ4xIjL2VT941mSQC4pV+uP5i+3lq+cVINN2AZ
mnWeZZJQb8djtV4aFErPxtxmou4zxTD8lRCttIjoLcL+D/FySvfgH5IFMCe0Xj6f
0QaPV0c++aUXWgf8TmkcYNGIWpvIUeQpjDquNc2v11ra2uEJjNWsmt81wD0+bRhW
qwMQPB6ywA7KOqHjsudB3k27iHa1meXhmZWSR+Ce7bh1QTRAs9Qy6mrcJTcEEsQC
Gh+HtYaDWyaZfelC3brlP5PRyO3cUii8UYNl22JQ7S1y2HKjNqc2VAMD+3eZURuk
Nef5rl3CgFbxDPq4V9ozanXZCflVaE13gYzN0/vtyj/eCgumTCQBqvK+f8KPhuBi
ZfzRZ34sF1gVRUJPbOIdGex9SX7ObYo9XA+oY4qZuA3cWPscfcwQ8XuCNkscIw7e
dIB0Ftdme2iuIMDY74HOg6qxnxOWbjphJOJHamh9FpchGHxg/+orlIc6nj1CmPZf
STZc8clA9t3Epb4uat6J3wqjelXJwzBX7YMSaEwVUIFeom0MTppO6JSDfgUhIIVT
ppWxi07UdDbV/WVxn8vpI+b4JccYN3od7utCQv5KqC+QJrVTstRvAaVgxZOYi7SL
ZiwSAeXpF7phD2OHDuHnqC6fvnfHTItM88CwMwtHyNUG7b+x0oSoJkAZm3QGtUvE
SnHhf+G7oStf+SrDw/JpDy4ZONi/NLplzE8sOkHeCdeLddtgN4O9IVU4FS/hVBcF
N/eHgpvObLdBIlHVKJWi/ZMlRwvJtxaiBaa9YxaZb0cuYYTrCkHD1Zf6PYmB7HTh
cqNA9oxOJc3GBRU/mKW181mx5yAZKyE6tr7/hHvtB+AvoCEn53dFhyWPmmMV9TIv
GbgBsq69ImQZcnmCBaKfEMQqLUVZSxDamFPUS2+B3lMfiY3k3YFUhsu83HKEm/C4
J5eEPVkT9hog/s7thiMBNLKdD7/9KY1bEqqjp2XN31txyVyBF18NoF0Q1NosSdQV
yQA0QC/z4icOs5E7k3qslAaB4xNk5ydtXsVu5EF96dOQBb7LOWJnt2vPIxhFZUFp
Lresxd58PiK0z1SUPmQRlbVZFngTGjZ5clBqMNE4Ki5xW/EtEjz5p2sXdrCzNlEy
0FMchjZNMl1VhLipqfbL6UbZl+d0cCm6/SBZ2MRqgff0vqeXnGIcYYks9wAW9eFA
X0Hz2ODpmpiZVaQhMdIlS6NyJQUYsyH8v4pTR1JreQVeWSYXo1f/UKuhs4y3y9EW
HCOrnLUdvFwDvL/CudM7fev/4ISH3DpeEBQLTmT0j/rp7Od7RrLskxuv0ZeOIiRR
haesCXyq93C5dKjdFwyoL9G8UcrbX9tclM8wAjeGpjRPdA7FBKWuEd4pzigsjYxU
po4jf9MkFrCRfZuamyIStVWhdXir3ExetDqLRmOEjenhQJ6F9q0YLw4rH2a2c31g
fOIIw3oTytEujka5Luc96EjBerXpCMUdP7T4zUj4eU3kx/KcE0P5GIHhBd2Vtj4o
lpslXieVo7loef/oaCHRmCx088uw55sUg2sp12aLw/GTgLGUIL5gQax4PHSoYdk9
clH0Zr/UHXnfUCBXyfKJ30fxZqzL6XMPOlqBbUpR8orDwQIvuSyN5Eu9rmTAU0Vb
BQGA3zy7J+euUrEVnKAgBsbaLpB3HPTYpzmik7SUd9JDjQ2pbcjAp5N2ys6Q8aUz
V3EQLBZkDMM36LdWLrnzd2T0BDBWOiYmJjSqFUd7omlxDekUW7Oq8p2TW4e2HmrF
uQa6TJ5cAdD+wyGCItxWKDhfnT9QpmyUsZZLvQgIUVuTmIUSyFlJB0tUz0DYUl+n
MKtB3HPxMGh924nDoYruHCnSVnQFDll98DkvwtlYE2Ru2qoFEnjQfxG7VUBK065H
V7se77++3VasQcNQgcIK0Mj1a8lrB4pedYyDtx3b8bGphXShVa0TQ4cnb5a+8ZLj
J37l1jlktnSLGo9l5yU0PYRI+cQddc3anJGBFn+AKEGHxNQapUdhYPBU+daH0KXK
FoNDgNYo1Bpe8h6t+oCHt23sNncH/EOQrpX4cJ8BgIssHv3cnRPeav2zOaGzKQrI
wWq81MdiNVEQev5ryHyjDK8TX839cFcwCcQc16TS59Pssse22oKhUkZmfQL+9f+V
XFcvwxr/nJ8W03AYBNKjpsy+wbUB64gWjPvhgLTQKEXX4v9GZ20yGQjxDesK7amG
qR54buFb054i+/gM5f6TrXJ86zxg0c06ArYEw6r7Ql0mDbSvTWLQA+C5OuL+kaH6
ooEed11KQCs0ojtDM8YjOWhcKtovkNeA+C7VQ9yoDv0vRg4ZZDkuoSB59fvDtaU/
6bQ8cYdkOBwLdRRO6yR8D++ap+Y8LRGH+A+FvIF9sgeEO5yIiNj60immA7fxAfLb
rVWwY70vCUrH+ep/Pd7pOjwDceoRU4Rl6z/Q7aYwfKGgX9u+SpWevExVoSc84ZX7
0bqVDPEk49dU7nCWg7+mZavAvihYdsC1FGKi8iZ2+Zpd5w3vyZRiaeyjxXLYwoWt
meyqIQHfnhTIr1JSrm6IafGbLqkh948PAYPPdqjnPNQmn5PiwmlG0X/QR5UAmHRM
SpYEuS2bwu9gcbpvsOtVKqHH2tObwx/0EkGXsCnz/y65Tzb7jEfnyZsFwm7tyZwW
GbJw3O1OvCri5IgnKqmBtri/AiBH/m6Z/YoCRQMkDZA1cgswRlKItojY9a3kiCHR
7cndFMahaMMdyJBeBPADSQYknR2VI8uduxd5kfyKNPb6EToPM8rzGKymho2+JGii
r0g9iHCtKSfwEdOBHB7nB9FE4tXld5oIcsxnb8MBt7kznVlj8VGHmAHz9IC3MjY8
ZlH8FtakwgWO4IIFEE+j5Gm6ZaJURp53Uswlu/OIfTYiNr0PigomrAOcWU16h6OE
+M8G6qYPAmXQ8DYKF5V4KlFltPRo04sTytZCou4P/KNoS9Q/VGIP8y4Z8j37sZTA
J1jUtgZFbMGiIQDTTC0maTRICe9AOTLKJgDiTc3rGoIS1nR0rgT0ufdHoK/aZhw6
+1m4qo2PVdgiL0Tv64yqeh+F/f/kfEGJ2QQoNlwwr/utxGf0Ql91dsNUbiUZcl2t
Kxxk/7NgamlQz9kIOuJWphLGIKSv8slHHRpBsXt3Gf0aDeYzTcawzCmxqFAwDrJv
yER02kGhNTgmAsvPo4c0XicMM0oQKb0JkTK/VhtCP5f3xcy5v27ThVcUwTBEoFOY
EWW26BDc9A+QeiJSFH0ofj9cJOgMlYEP4jKOFDRdQSsINZ+sySvs8xdH5wNJhIvS
FqL5+DuMRRz7EdFcUG4ZExGKvidi3R4p+HGPWf/qJw7TJDLoFnk/u449gYBq1+g5
xq9ArgdhcDTSEXwgJ4OBTgGHI+yMR7zDeFCYPkrVNfzt+3/p846919d8n8NhPXZW
QDo2P/3Rygf7T8Uh8mydeS6+VU3P0+PHAU4iHj0DOZv5/VgFAD7kM7UTww6uv9+g
SsejNWVSeBmtPdTwuFLO8v+XzDJL2JO/ft83HPAJK6Vy2BF0w82Dzhd9KA4CyD5u
FMixpgSrWaTJfKKVuwlC/ujlMQrEtG0Mh5ZVsGDg8QM4fZCSIIiS9KetOIITDIk0
3QPZxZyvNLJUZQn1ZuiwQKV41MdD3C81G0LTT98rcFSzVRaBMQbmESGv5QFCBlzN
D186Ckam2ZrEl7oCMMoQIcvoKy9dFSVLSzpdYd6/QXYLcVFupH2o5oNHFcWba2/m
smSJBN4Ea1C7JrZ2FUnpU20IsIh9UvynziNizLyKT6JxcvIIRYDWryTG3YtznEZQ
qERI7q8a8DbU9cyhYvO7knwNQPvtQ/8y76NG8bEN//IbFhYe+2yuInU5n453EbT+
SXSCQJvp9TpsfYb/++0h94niZ9EETkx+UKpXPrB6E/tYYSiCVsLQWtiENq+PWOAa
WwMi5bX5ofeud2yOgtKqgrkY8UBCeRPTiKYAKuleT6OCUfjbEIHm8GJc3yjc1IsE
lnkpJUA0TT6vBzR2bdTgwCl83AlmQtVxFUb4tSEzwkb0dSiFhimnJo9LoiJMo4dW
klbyuT1aBdCQx37CNJunJlmKveAqpjALi3NT8kUhl/Qnk+wA3VP/IAEY22Zed7bg
2ZuY1LjNttXaRnKFQaK9PF/D4P4i01dLKLXNwpzHxqkFBb+PClfFhOMHl7D+snWd
tLMKfnIpYCQ7pDKRq0m8yD/9P5vJ8DHAIzmjPs/m/qNC7bINqzNWgeov4cwIllZO
aHNYdKMfi2tJOaopyuiFSMswLlM+VNJQ718h4QMbjNd5WguJVjMreIiKcM0J4XCA
TgWSM0+OfqWjnDwFQlWdERFvaPYMhPf4pCKs2Gmw64I8+mYZLWIji0Ya/QP12op2
vEcJ6t+n9XGO6yyQPnR1ooZoD158XjsLEAT+uvmSbmsFBfTU+6vn3lSChFUChe4S
pX6tUo2B8Du1+tjt19uU7ipJG/6OEgRj8/qlN0mk+jpfG9yB6Mok07r+cOrG1WuF
ortSm78YK3if78st6P5SglNaz3XuqDBKDx5+AVruG0sEcOWM3BgYclT+riDx0XqJ
59mYWl3sT/kJPQ6W0yUqc762sQ4qg8LOIbMWdyMXuum4P/MBnYIyf5AGWKd21ZHe
gewQh2YOW0LvqxvcwhBR6oPH/AqN7wz5cd7HCE41DyZvNwJqB0g4/8zbmBlDzj6Y
YIKJu9U8XRWKp0lkl8DFllhomlpPu6U8DfJWRm7m6u1z/T7mbx28nP7NBsgjq2Wz
HNfG5RLSqQ2WdEfHv6Y0n28vNjicaI4P8ty1PyyAIbBZLWCwTUBOq8KXY+q7KlNF
MxVHY8AmC1FCIyIW/ZvGz6fDh8u6uyZh9wl8NzhtVvjdwD6lGIhEVgUydOg0yHoY
AKmks3vxWVES3QVquOvRo8+tGR7UJzPhdM857t7wt4i5IprZuQtCfAJEBvJQGS0J
vkYX9NH/zIlSA34GZCuwzWY15xSnw8PWcS8+35A8vtUTg9dB++3tGcygINULUdR+
dgwihn/C0DvF6qiTJK8aY4mttdjPvQHcizDtcgfNkrKWo8g11toa0dIr3Id3ksPV
gMGVOLsUJtQFGDY/fYQON58yocZUiQHRDiRIePzpe6Vl00gqQ16OjT2TK8xW0VEo
HK5ZS5E50bQXE2w7iqH6F+4Zk6JrBWD8CR08FqUx3jRu03p40PWGzO8/D+guE5GF
RlGLUzKuKEVT/JHfPXTKHvzuqI84je/IRwb9N/MFRddvMvS0zhyDxxgiqIhRTg/r
KwhP4yaCXgzJnUUeaWZB4gP+ePV4JXRYJdXzI+e8J3te4KsW44Mr8r6lfCCSe6tm
DLzFXNemKSx0Gb0NLgeQvdz3kOBm+QdQSCuOZPFuKqdnuHpjtO0GWtBogueS5SMm
IGuHovHxq/8/nwjoSkRrPxlDKwf9mUALpsL2eCZHSZetZ5GE04yzEH4GPrxFmctN
xdoV09rz90WhsH3XeVKND9+IY5wr5TpOsnpfWVxBvJZtyBKW4+Zvc0l/7i1Z2RZZ
t990Q3JBas7D7yD2XKGI0uBoH1ORFrLwF7F00WmNrJ6xDzIs/3zWccy9nsDVddmk
k2rdgmIeUi5bVXKMI0Oz46xO1potf0i0eq1j8yEzjywMXSIkcyAIlpgGdpBhKEHc
KEp7tF8Wj9SU6KTut6fgkFZ34HPHnCUr7bjVoIe8NOTaH4BtMKCuChk4xPVVyOQH
cAdlJbEW9+Wg4LSYSqMRXd8RLI+hhLyAHvgu6HeckqPFcdmzALgqissIyT6DCBo6
jMtbNXn3XyP74WgHPYPvT6RdioSSAopR0+aOmEyLYwxroQ/RyNIY2LOT/03HflXl
TFbZG80QAm1F9A08hstPFqnvByEGKA3PhCRYgL0xjr72KmYIumBbZfJGlgieo256
1ybyuuWYujKoZjBo03hjaTYW1NebpKV02kxpy7RBRzxuIY8UwNnFLF1plezGfCgd
u79x8ET5lDdq3MGpQJ+CECwFe2LkEPlI5ZSqrxxKCd7ga41Ksg7m6Hg2pVv1kXJX
mA1Jrgt+zhm8UAwti0z2ChKnaTnOGwyRJ0iGLFoLIcQ8s2PqL/OVZ+AjGABBWe8Z
HdQVsbxEKQuF34VfJA7aiY6CN5zZJsCR0bNLSQSVYWLexp33wHKpvROPcfJMswu9
W/KGOzMWoJyX++Sm2PnPxeYpE+JuI9Ljg5elYwhZtumo1Q6DxdZZNBHP27hScgu0
UZ/4+X/4yAh+z595fP3R1/9NLAxNokqXnRoFsqzxtSE=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4N4It1k21lh1qR1aobAjd/p6MR3OJOcAnSxozeOfWfu05i8YkC9cecAnn3Lz70n1
DObnC+1LrwNekpx4PL4rkY2R2b431RkpldCJ8ckkGrk9uX4ETeLBronTOVKLL8Nz
KUnrDpgffne5VXtQ8dft0IYnp2q2KtAGwJGtDaxXruNOdb5dGSBYIoRJJgVolHB0
S9I6F7RLfbc+Ch2H6Kin/AitMe+72i4bG+gd+nycNvnQ/ydRUMLeV1OZT/WuOQEQ
WZgRnDeQ1lJS3+uJqaj3qkG/wVGxRB1ubqcrR1LovyWcbyA4+R/c/GiU3SsH543Z
wtCfiZwgL/vccR9TJBDhSmrRCNFm1yiwCKknQAJ2lu/gYfYu2oMeiNLynI05lzBg
BJtm/TwNNP3u0wCGxgkzhm7ky5VSbBC/WHJzo3nc+2tO6p8kN0YdU5ObE/sc8tdR
ZjOPQP+KyZZSFI/5gf/CoXvDU8vhcp6VN5v7tE98kxU6bq89dW8NEFPH8+tCrK1L
OOOYIH5C4aUZTIcDmrYJASukEXhYRptwuhqnegdmouwKubgz+HhGdqk4LMiNeHoJ
qVkQjsc+0MDlKq5X3C151YqG5mivIJSMUrMRP3US28QTBop0RjEFZ+xAJC01BQ1Q
xJzQvH24feiJz2dm9oqr848cUQug22jOdPgDcL1EKr0=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcFiSZubzMOLSQy18yFK1HlJqcDDBmviFLg94LhOmgDkmiryiWvvPiWUMGFmeQRx
3Fd+1rnYYNYuakbPdr2Ov/OP/3qAOK2irwRZCw51LtlO/zXlfq+X+1eK3xlJRIK7
lbuiZq5SxPQXgJCJL3TkaLXb3eXR4YeuWRNRc/1ibUnGSxPC9A8KdcqpMmz4NNeW
7BllY+vWgg7gpVzELG5Zywj4xsGxYbybmZKGO7t4Y5e8g0alxftUVPYpZi7+Uc0a
yROwfOu42xJ2d3GtMedIQZLhTM/B9o51DL+OquMvZI20PzOt6I2q7HJf6JmMOwvc
mm6hZPNCSEdLHY02t4jeK1weulPB3GD99bgemYd1cY7zhkPVBi8I2L7tXwJnpsaq
2K+IWL6EQHEk7VZlkkOZDUlZq0iVFY+vxLhVLZb1gBVY35OMKMNDX3pwO+MlLSB/
P9N2a7INqEXmWjkyLUrmrUI0PdhUCPHN+FkKOuUeMoET0ft1mquBK2M67kDAPnIh
sYtz8jUyes5yPwORu0E10vi3IbtDM5glJx9iWZrW3F2CeyNW5kr3+3sWJurqoOD8
6QSFYUqqIknL5k1RYUIeRlA9xw6t7Ux5Yw+QlYn91cJ68P9vDRbgqT1fREeWa+I6
ygafTMCXll5Gj35xkqUbAis9GFq3h1nXt/v2hZ6CDDctdwlnu/eaxvjt4UTmR0cr
ghJyA7vrETO51s4WhMP3UbjWv6znsPWPReFp4dHG5MlqjLUxdWr/ONCBmfZrxm3R
J9pwNv17ViXKI+VPECNFiIKkwFhWFabk9NT/QpNPgdSxkIEVzY+cU6nvKbXq3i40
en+w/SDVsEREWfEwMftBusiFFNwJl7QNrOclei2/vy7WunskAmF/HljKVzZhyBow
g/6ae+jYnzABQQ/jpbF2KrqmJLxJ58IKYUlIqXvG14LGUroIx3Oh5PbJf7guyTWH
jLQB/vUi6G3S7SGOaIlXfv1itiHxpEI+0WNdgjRA4I5p606c86h7EQsCXFc+fHtX
qhRa1wZZI9hDfAJ2b7Dbi0iACBwT5orntppjPTzs0uJ8b4JABj144EUQpcMtD8Qm
wk3lQkZ2CfpzEgIGbsyziHPk9VjKSUW4ZAjDwHNREu6HJ2WAh1JqjXfQetCu8/OY
EdBrVqpQHwP5M12TxQJLVtmKfaRKNFiJ8Cl7Cgg2ZnV/IopOpEW+TwdHaenLQRcd
ttmEtEGqFD2LZczMzclPDZD7JLZwTioa0NF3dijoFAeW0I1VMKc/0SSfLUmTnJCs
HdEHPSnoX5FABn8Lo8cE/zBeEaW9TNwlr3pAZDNktddFelOAWT4y19uSXe2ApaZo
LdOqtqtdmH1cJWzMov2/D1fKskNkNZk/ZZc0I7Jg3wYhnMU1oOii7eCCMGhXwfet
o////vTIWRpoit9Vdh8UAt2zzMlq6D7+JdAppBZ9/ovSNKc+UzOQzzAJUJG05Eu2
ZRoQj9h0Tfwlt6+gwfqkkQ8FZsmROP0mnOPzlWS4kCRCyEo4yTkvOLwAVmZXrL12
X5WfGt5s8HcwYHLSBYJwFyr3jDxX838q5OqjmHqBkz+6rp/AsiVHzgIFGlk/o8ND
0dzGl82v8wzuPjgil/kWl7duhC6s4CR6GaGDUnBworSLIyoM8vdIabdC7erC/uYp
4bIKfuKsmrhxa6yYim3THPHz8PR4+D2Gp0LIGGBFKrgaEGm6y0meTNc2ZOtkqmt0
wa5vfNCnq97SAgkAH11sAYmkqYIAu0d0PG53vks1WnSup1qVcjdDuZ9WlilW6fDN
nOZW+h+R7WKl5A19lAhICGDYVZdOiUvdkI4ZPyKuUVI/HMqRAKFcZGbA7q6nuY1P
MdmecLwlgX1+NXGAQWrUk+MCB0kEs0dy4cR9GfRUXN8Wfpj11TXmU6aPUpjN+YUv
voiW5AxZKRDQsMpxfnyop+scOJvg7B6rF5+e9+zDmAKHWq5lsEqrYhCE5agBMl21
UvGKb9mgtkRDOV2uimxOCZ2+VE+qcHCwU/EKdGJ6W1HnYhka9EBzFwuDzPFbJMi9
tnIT8MX260PwXezqkLRT2qDoGskxtWpA8qq7aGmc51Cwws0W2ac/KvR2PziztNid
CJm/m4Rz1zJ0h26/Iu2p2WFQIw/FoXOHWE7jq5eK4tJPp4YbcA9g7b/ki7ge2pnL
PDGVHdcX2iKzeJbCnrwTcvZgj43pn0XoJ+S+Zx7DHxYaE6VA30nV39YVat/XZWxi
Kx/fn/J0AWca9uyRIXux4pXEfOeP+3ZZPMJ3Ze8hx97rP6XPtcthISwgT3ujU1mc
pan/W1DMhwsWJf6iBEkYBNnprm6U1AlXQh/dmwPr+OtnNjSWxAzJLK9uL8md2t4J
Xl7qvAhlZjcvw0gQB+d6PbcoydUe6xWo38lGRyOHVP82W3UsQYD6ga5wrPOa4CX5
LQdD/ur+u/eeI+0v3sZoQj2P+ektSlV89e+88wGIjrkWYOSz4I+hBLVw7hjkf5wX
ss+mwyi0gII6UhHAb2gBprIBg7Vetted55cp4p+dlJHQ0YDjTHOc6E7AE9Crey9Y
kvJiH67p7V8Ym/2yV2wRWAyM654ANwB9yXnr943Ywiqrz2T+snDFLXgSEz7SBuQ+
Qb7F0cCJfwlZRP69d0frFAoRElImvCZCsJh8rNaTvw3jTPNsL4KOp2SUsk/zrGcR
qlBtNqnAbFNDDrXs+NdAkQjRN2XYIbwByqwnHrK2HeAz9pROtH/QIwfj9HpzqzRZ
RVV1VpB3NKD/dk+oVi1IZJpHlYAFX1d9M0hf3hjO3+SZ+yFif1M3eXzN2weTK4wA
BCQAx130ZWaAWbKs7Opu5y+ClsmerYvXWUYpNARGxhbBmiWrpbZokT9mYMR1VkFk
`protect END_PROTECTED

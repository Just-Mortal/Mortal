`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9EY3CqAGQJVkKuk6OeafJhTBVnPdqc8Mv+X3kD50zQotzOsUKFjvAsJC258h6D7
5KmyyVW7V3/V2eHf+oFj97e0IUSCGjjFTAhxq/B8GuJAeVoEiZX2AD3w21vGuaaE
JnFqjDPJWpoaqK5A4LeIisFUvZbucQfCTYyUldE6siBTiiJVSC176T065tAF2Fdm
NPw/EELvvLa0oyugnQj1G2GxtIj9bU8ty1mCEmZAHDX7s71vfYsGQscS/pBRsXUu
2MsU7SxkTEdQ/5BTsyShrEUtwswvUMsjKDndlBRxvVYgYzaXMASMWvtHo8bstkU0
EXqm5hjcVaAvSB98+vNHvR3Q+NyUx88hUbiGuosTnUzlzqxr3xnOOh4kdQMVSgTk
tsX2L6Mvn+lAcDb/EpX7WyJsThQVe5rf0Dr7WkVB6++zuHgQNBYW5a1mDOzlw8lH
kYXKmKvuCjO3n0RhHl8y2l1D/JH41fjEBTRg4MyI6yMFRll8xGOWwfTKZUIdH8Nc
N8B0GzdlZ/mk36q+vdwDmG4drW47f36XsePK/JAYBmy+Mn3creO47Uhpg0aGtmBh
c5mQGpysc5grWQF0lCJh2aWm0dLWmM54/ufsDo5X2ur1XCskVhe0D5DErR9nYlY7
dywTS/eUgPwHt8BG2jmuGZBEVw1y6GdwrxB0q6qnG+Qd9OhGjBOeZadtTKollb7E
YbB3O3EO+gWKoRK43+FDl/rP69bWK5mnd0qMEeNO3GwcHA/LrnF91V2s2vec1ywI
CEK3exv6ukyry0G1OMzA9XcJSYsofrqEhg+z7UncNrqzuIinv5vcV2G+/y+mgMlf
M12ju4J5yT9O+iGV2T8XIf5xY2zROlkgPMIV85sSq+CceRn5/vTpuBkr3XkrjrkQ
tBQxuJ+FwcMBxHGOKXvO6IjwaDDu1p+W8z1qc8e5ZPFIlA9N3+b3dkb0vpMSmB5D
NsICAqE9CgBnmwEPOqkqhvuX/5+bPkklXopE4HuVedVpcL+kRCebudBezjyF0VBb
KYOJtlf4dLED16cAx8fzmurkzaY6SEO0wi2LVBY+DIiY+GTZ74GYw3Ou66j+6R4x
76IKmSCOw6W/tiR3R3Y7IeCyVjoHZk1DMj75S0qSYxRqhrSo5G8LFPn2t83lSEBy
kIuDm4oMOgpNK/UwqbYBKapooSJQsnH24pj5T37kojD/q2TS497jcjXpPGMuK16u
4njyI1HYV2tLapJ3bB7TyZQvqsLyCS0U3gZ14srnLuCdSohH1IVBI7ZNVhzkpam5
CJRHArAujSrA6DNcU1QLzu18jaUM5poYeiwHlLtGVFheRpYQ5TnPwTBXwhylXhEp
shr+0BH/wVtlt41C5qKfYBiaJbiLjJ0BfGh7GcEW1x6A6m5v4be8Ee1a2ZWpUbMy
I7GBfQpqe3oQ6De3MGZ9+H9jg4gZWZaVqJ+frxbmvv5rRtqLVRQMwcIsFYGfHFgp
NgpXV8pqW8yn/4vY87j3GKlD6pdbrrXT4eaAwAu07EY=
`protect END_PROTECTED

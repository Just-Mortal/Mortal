`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8YcbBNw2PRb0TxoIFPbEEAs1nqf495YL6Wer4nL5NS+Ru6HKyofCTxTToY/RXKZP
GXwzX22iVTQdPQpk4H5H3bLlS7Z1Az2/u2oyMfOJ7QN7Q9L+45dDtCjuP5JRIfmz
4ie00aCXM5oItAgl3TMPkWXIH/QHN7qOli/a5OUaS/GgmSJuxsOTTrbXOkvGUruY
XEDTb79saqMv4odMvisc3yZT1nXxnPNrlm8RTyj/KpDRImBYy3B35izqg3XnztBZ
AjfY6qgKiBtA6tysyI0z6G4A0LHNodAgA2ZCM1+t47cFHFHCMSZaL/xopV490F/y
EBKwqj9+R2jWG83LodXcQOMfFjhuJcV6SS5iyfVVRkS9UbveXyXaVn2qxXnRW2M/
dhRASFHBoCPQU+7OcuvEO3cmPkd8RaQTu+GZrqJjud02BKl1vTfkesAzY+oSxwtf
Y4SUX0ci9opAAWqQ9PjOddIq0cUnX9aVNTkihknAfdZE6EN2o3Kq9v8Zp7gny6ve
9eMNr4eONBSgSTa2zqKkXouTj+2Mu8BMNneUR74GVeAQDx7XeYY2IFeYtSMkW6wz
XAkOQKa+VXz4R1pjyDy95oZURYfvgMnOKHkmhIKi7BOoOlauM3IXVAV0RuMZFqPG
BSPVxt4kCTLhBVEkoC0L/bqH5KCSWvHw50Rafh9SxHg79i/MQBqpZm94T80tuV9u
gg86KwGsdsDEL4sz6galX2vM435LoNhVinP44F5U2kIPmMZfwbhEoqbs/EDOmVOt
okzjnnKVzKaZ14ROdtK+aPUEwaqBjqgCl4qGsvWIJX44/KO56Sq/oWStiA76zqZu
7fEx9ufFLpz37BUESMB4Yc82JXlKAozztK1WvuL2/Byl9WPCFpAwi7gAToMQEqzD
X/JxunkU0osPCL2e/50LTZWBZKNHIMsr5PdSmKSulhAkK2W1/iqc0za1v5hFuIAF
RmEEYYFg4njTgh7r13hpThUY8gQ8VLrSfPe3Z3TxyZYvnHhAb3YTU6hehEACfvMw
uHr+QYt2/h8IIVZPzUMnLr9P2s+q7nS5Y9ARlNlC3yNCj+Qetq8EJZxnIwM300Me
4u7h8iJQhcN+gib4jgaRbj8tPM2R6W03CGKQnvlXCkBoG1rk3AY01Txn0YONZvI7
Lc1JvHKdFNR//teaWDfkKf2b1aSWVpAKcBxEnpdKJMFpi0wzyJ3rdi7z80V4JtQa
7bSmMBkW9dXXgJGBtDYFxmgwndKMtubAWItC1J+0nHHhYEsPOWDzrVbaISv4lE8l
ZqmrdYW52JM12W5kJr+WGzZdLAqohCcvm0ZEVoDB49UFYPCAWsIEy/aCmK1UfLxh
1ug5C/T18uMNw/Cuh/07tKnmTncq4wSPZrE9TIiv6AnWhpqwCPhqjMCQxgZKBGyR
K3yrGdd8uS5p5KIfHjplU0YBCB/UjuFhsL3JnWgUsNJgILBkJbrIqLJXERThDgQm
7Yqg1cHgp+1xntQi6yDLJCM02sn9e6+o0e9ZkKCGdhzekEQHtUyNSqovrg1vcviG
ywsMOOcSTWiSVdCJm6IV/Z7NwC8jCoP90QcXlB6sU1RBY6zJe8NNSviG7cnZWgJX
F5dggWaHTr8oOOrI1Tnv1uphoNGzZwmKpMEGoCpqtEeATT0GZTAh10VdCWPXKGGw
ukH9uscIszeKG/mZB0LN0ecZRGcN5md7eW4oPmM2sOCnXhZwuu4AChX6f+VfFSdz
M/teVSL7+4+csjWaULa1w5Dcywd8tlAVIClmIlpv3EVxbV4vwR/VEgX2kvp5/s28
j8/EXTuBa7cCF2gziKqYepYXemfB38DuCobqlz8HI5Efof+MSmhpf3LavhrwlOuo
SmE5kMyF8i5C3vVNs3FbNlIVsovWSJtEN8i2shlVo/YaXRuS7Q9y1FzvqTmZKQOM
sSdiZTV+4ZzwUsY7d/+5ilP40/WOsoIL4ZSQHxN8Qx2T0mB7NJ1NLO20zPwNe1Sl
eLPfoDAbPCA/nqMr2EeCN+cy0wvsCk9k971B3IIS+j+69XXOBg/f4MMZ0+/D5A36
otWOKvMYHDuOWPiMZb3U3B8ikvqVD5eDNHfDpMqDBOk3mhYm27xG2U/ha2/x+Fd7
K6wYRdLAgfcz5XCkTC4OtiS+UMVsq8nIMOxtRPBLwQhQVZublHeA+TBkWec4nKZq
waVqMSn38tkcU0xPuUmJwtzpNrcxoKLKvkEPW854k+s01IIFArekO7uh/JwZr0ZN
GLyBNhILiXUS7UawfZN3O/XewDC7ilLsjhveg4buAflwiOOf9zc35yMcZullQ7Z7
CsjjLqB1kVj3ZACvP+X8WfagdvqBNSJaNt+DL2RZ5MHnqKJDujQaF8a7TI4w7L7P
3Bhr6+RVhXVld+iHBvTbWbgufRn8iIUFGnEuety87XPy7lQyQJqZgvY0g9FrWNb6
OWhinWz7kZIvDFyYYHUjVuDDgQzQr1/Gh+yVmCSxo9TA1qSRKfiHiRb13Tem2/al
IDt4FL1YTs6SmsDJgzi+es3+t3HhPMqZWpwt3tk5t17sETl2w1qbjq/kX+T2Y0jE
u8Nf4FTyafKxUPAZlrEaMhAyRVl1K1eCmGr0A8RW7sE/3OxUdPepkpaqITsjEoLU
2ibIxiqUb5ABhK/2r1lMYsNKgc5mapdChiXwNc0kdJksIZza5dLBiAUzzSWLptP7
8srE/yOMQUgwUn0YhY/CRBP9C5UkhYBEpWF/WxyH+rg1/GmPmgFTqfF89uGXyznj
WzHmxmDE0Vs+V0C906r/k0uzSPAimsXBxrEb9eqQE1IveoA8LdswRlXqfAptC5L+
BVwmHs50ZXr6OBzv5/4NPg7ZBq0+lskhWv6lTdH3hLn61yx7S85+ahVZijfddrSZ
ZF40T8DE1itjnCihWTwgOHBhajAmT2EnJNkVEUKfFT5dzqiLDTUORTvOuTnsNTEn
+MQgvzWfMps+71kx/TCRTTX+FU42dQEYxh0JLZw35iII4jKwDLkzQ9j2DD5iOQe5
VUz7jRx1GnlfseQubWmf3a3gSIY/RWMLPaJygQdeGahgDBxJbswSQXK6AtjIPiXV
oiHhmwINHyQdCJeF4yCR6nnEkaa3alpSb2RuA4JvsoXEjyRaa5luOl/0UShIePgQ
DMXBQYmV4YPknyf/E9ZQe0gQY1Re0J87EbI1IQggn56zZK+MAXWcdhpKvgjY1Hm+
VkAubZ3UNmVxw5zvLt8V6JQLKr7qB6NvZS4ylXQFvP1c+evSzhD0iQuu6SSA0QyX
DyVhL4ej1EMUHDA1EgTXTa5nVA44yygfukZj+VuBSOpiEh+EwbB0ixnEsiZYjy9R
8zbW1/G9XZRD75exnBdGhdu7Gt+qq85fwaG/fz24Z1TMEZtPXFSV2wI9+1b6R1Gp
J9Z26v1TtElng4SaRDAMURjgsy3S/rvXnb3sq2F94WFr12XhWGYOsL88zSPuQc4L
wqYsV/ugF+3KHKTl+9K3iHaaWJJewlads+HYRQMmX/QWC76OolkSPRhCez0MaNA6
ogB1nPGVSpn9NyTMNBUCrSkOV+0jyn0ExGvLkm4KDjDMK884nVcVXhXaFXzX+sL2
G2IujGlxMPayldDlGMf+YspmQxzCOC5gLy6BxP2P3CZtkO76fldTQlj0LBLzLT+I
DF/8t0foJkeo5iBQAbszobBVS4Pi3R1LKwRskd2d0CqljdsBN6ZkqhYDVy743cfL
1eskQ2bJe0jtSXtaPWKZ9siEB/pyExT2n5CbLsWk039ydodwE/z7RqTKwl6QJPhW
N6Q6U0I6Jny0qBRhohkwOAVRiU79/XrZJq7t0zSwWJDKfVcLJinJDSrj/753m3Wb
+JAznufdKJT+jOtSfFInc6twJlepnJIgO8VM/cXzho+26Vq08uDoGJl5aOnYA2+f
Xz1YkxO0O/9ifUDQ0Zd36dmmITSO6UrgRg5FzMh9ejViBbk8Duh8/yWoiAWoLlxw
eRLwrBVfumpdT12LFS6DY3jYhOBi3ZEr/hz31ibO00G6mJa7UhuVSNMv/OgJgbdC
9QIrXyDmaqKFt3Oe92bZWXlaWIF/4If7nuEhqkmI2WNhTf4CYywTuHLEcR3CSirZ
w6N5VVwOdcnfeS9m6ZS28Oio/JKumM6d3lUthmFG1kWG6yrND58WHsEmsN5cXwkm
/g0O69NtSAvZAuw6665+sLWLg2QzaKEhRSsnQdPJP4I+Xlx6JcCXYf7ZyV2xpDOs
3Sf0MvmrCfIzapPdUaDUgOD5Vpnsrjcvhamd8iDbp3kVBc1ujibOF3ftHgMVRx5O
oTaSKjHB65GrY5N8kGcMqAaVoRIXsvUn53FPSTK7YPhEGM5cDk/yvUJfOmBEONqq
wkvzQ0HXhHUd2PQqkAfFAl7JRb8taEliCqGjCkXmsJQCHd+EW2+njAj4UN2WbPGF
VP8XXLEKrSyyeHl/F8Lyza/O1ihjF8+LakmHIz4Nln6DCy45NSuWkaq0TDg48mM0
jM2U+ivChyXsI9AGyRhs0z8DcEi6iVTkypkQV4A4gtm4jR78kXKyZHWPObVJ0OOR
NGmUQRgwP2H+hY6DDxKvivBB4zGAE0/2cPV3AOFKyVVwdIIJG0r5ydLCAGHsC7k2
WEuoT83JClR0U5Se8jGH+upGRzmJG/HhSYNDpFLdzivI6VB3hy2kDS4mcxKNH4Xt
R/DdXS+5bDuXJ+HFH47bi7gW7LCmmR0IsgN4aDvYluXrsLmu5Eg/b2YXYisideUt
mIowLTReXTElnZlscpMz+xIbPrbyX54an+rx5j9wnkxMO6Fo26RtDrocpOZUvK8S
/W2DSctkN5iGNCJMebkQ13wJtyiPsb9EDb3LRVWXkVIEXoEmO8B7agI7qrqiP/ix
dCKT9vAbuoD9v9C/jquNr8Uu+i0MmHcHJCXdA2nC1CM6W4P2QjWJRmnQG9sTfD1q
n3mccyCdH7mxeUijRBpnParaITfglgW/vvxcxrzXDXprXhi6ik/WMnipIMNS94Oy
FFjBsTy0vACNkjbnyPWkG2Uv2+n97wFahZ5ZKejhP3arcO0QABlMk1yfJomtZqEc
b63UyWa+KVUBWgFA/mvQ+KbNC+qI0/OJsCyPCwd+IOyFtn00izapRXXqFll231jH
zqCJ8w1svraG/XJBV2ImMLHPjhY/wndbTrxziljVRrnl4OpOgAtIgOqmVaAjDIFz
UseInQmWAtrOvIEeUjW3NWyKmlzTIsjKTeeoGgYpTSDw3rVAPFxXqwolHF6miGnj
rt3U4/PcPJPO1HJdC1h7HT3m6jRspOjAGqRxDvO+TUi3HYeu815/WK76kaqKhUVP
Rz4wcZp7INWXnvAs0vxyeB+3n7qc0vAc5mWSPQ1/+VwfN+mPzlv12ie+mlQqid+H
H0FE5oHc3QEZxVc7WRsI7CeWA/BwPhuSSChyShLVElDn3SsMMm+wULgcLC5q82QI
U3DS/rypmyg9e+uXaohllb1AxK0qh6eektHOxdPXkw9tDf2b9Q3Ig8WgUPSjTRAi
T53FBEuqkcOGh28dxFSR/8AYDdPFA98MNO7Mk6XxO4GpTJ4CW8fTV34talSh1g1R
MgEXY6DhK85q9LA7zyBiG4gZKy+SlUZ46L/ptF93xvBAQLj5svw4yFaxftW7o88A
RxTsMmmPxQVp8zDg9EnQIQNYia/XLKg6Kl4AHpPwMsimo0hyQAGBtZjg1N/EFxrv
bwq2xWjd+QsVlxMondHmvkc1YX27NqjdVNeMx0K/ZgRSJZcCJzGYaQjhtDuhdtmw
a77dh+HgwrurpFF61Vp/zJgWRaCxRfv1cZF7cZhwyuj5lVEA+Rj/suFdyZDOL9GO
czV0X4PoNCWGSpE4ZDmlKcWsKnsUCGVhX1Ziw2U10HVa9YiZADumyCW5G6gvutzm
mKRIsCd3O6XsfNLpFMs00tdyK/vTtCe4azlel1BzBdIUopA7bWMv56vnQhCp9Jzw
qK3GdpfJgIglflHNRoAb5dNhKer7l+X2Q/Qv3s/9QWFZ4MdtlL4svmBVKLMX5w0e
StPmfPDIuvx32ADBlUb5j+O19ewNt+WCnCMbXfdM27gWygNRgjvxhFZpZ7cTKPrt
By3SxrYsL+dyIt4+XZZPLwDdj5a1peOAhTYygFA+Xd7w3jPlDzGZioJjGZos+nXW
qxZ6Aiygh/VseJxiIwuGAz2bcQmIyMAO9SOfkOSUXDz9dG8fd0PBvAJybCYICwt2
Rf8Wnw/2VP3EitHEGFiy5FPCG5uoxg6aY/aADPEXCPihm/BUwfc03SayTcNewHsF
NXmHCPCJByDD9U27KhKPoKXyx6Z8bUuzgXcOwwd8FqxAIEHT2enE+KV40pTkRsEK
mh4vBd9dKbBe0fncrHYqo2UT6G+zc7jX0+Y8XD9jSlz41+1grtpig0OFmwT3If2V
aiK5hGuI+QNlgycwB+ZZol7tBgl2wxHYywxU6O4uedASg7TspmRvj/ssxbWhxrfV
85o2mvJ0ICt519um5+8PqlsMRjIDvhIOF7g6WLoEwYbNI/KFvOJpnGlKA4p0q+sf
9vuXHB6+GKt8JAPtrHsYEgBIYgK9lsm5qfm9Sj08XQLN3wpQ2U4izAqKVOop3oaA
mT9EMdFz7EMguMSzq+wop/GQUpblItxQDwmokCc5yfLwQmZg2pKvCJdDzNVvbDYJ
0iEaR0hAjui1zfQwAcAQVgsl2kSn6/SHwHbI1dCKDEYyA1G4IqmL9CJejEUBFUlv
95JSH/nAk7IrfSD0lfxd3w==
`protect END_PROTECTED

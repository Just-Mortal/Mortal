`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ur9RvRk/G1Rf66uphH09vS99uIj3B4rc8uvYhUKyWeKjaYsTryX/Ob6E25xBlTn
3K8xxlGZxSnPEBDXutEjtKL1EZiIMjPCzi+5rs+MusR47LsQpgvPXacedLkLpUDh
eiWL+tyd6rxY/407If9hTjNjiwRx8bneWhKNWEglOQyN4OLuF4QdhJztFcYsVWds
QnJ5gUjPGD3A6L2iq2wcYhMWrXkkZ+LNAOMPQLkY9OrGoPnGdViUoqrT6U255B0P
miGf8eQWd2eXORt8zx2G855rDPl/+TRWonZj72EtVLmS4jqPkveBa8GhQKVaouNS
oFr8cr8+ISq4yon76Km8CsZSxFX1KmhW5hZywsN6oQNOhOiK71XtEyqkvA5yERtx
ImiAyUahDnb97hnFFTfKfvk2h6DrncLqUKa9dq+vXBYnhT0SDwVunWLoMylqg+EP
to/MwyLnydcDzXWeSThUSG/n9Dan40mR5G2UfJYwomBLNufI0LkXPxMwsRx+Nxau
Zgjxl20YLtT0rUZfVallty1WXS2QRYP4ptcE7WJnOBbchu6h5ItgDROA2g3KhVpz
DZv6nKavXghcrRg8t/zv50LWwQxsA/6RTKkH2bqz9GOMBFeAXSJYAQUk3wbfpeAK
7b3WU6kESx1rnRlbLU7FpNViwdi+auqrfb8qgnFmyKk5YRn6j0y20E8L+J1quk1F
7cr7/F8ckWR+lvjFQWLeRkUsQLYfbOpIVbqNyjbHz9JDKXwRG5kqkDmYQSPqKIlS
0Vs2Ke2TdxpEFP/oWvuMO4XdP+xBUgM5AO36B85NAahngi0l8KAhBAWSmVa9rDc7
nHmZuSFcipMKABqOAnEpOcCa6vo9JebzQ1NJlVRkXuZYRfogr/5Od2UTyBIdgbW6
bT0D2GpFpeL7NTsaQNt3PgVb2sQXkxm9aZWQmyOR8xQBZzQYeeOGX/kuETwYvzkS
0XSaWJKBbMOaAl8BsZiadO2ITBFVzPNTNMEEcb1LgnPrUCp0+W5lianxoMS/5v/k
v5UwVOJi1VRGELw1befyZH4H32XeMHT3LYvfDlScCR84kOVQ5oOF7CaU8AgNignr
3RsUBxwqXoOeqKe4yJp1LWPvxVY2ZGNCorf9TFHNmeHJ6eYWilsrbtFSiG11WCRf
DloIkDRK6SfZpiVXLLpMeHrsKUFARGr3ltY63faoTcelg1mlJjiSE+Dlmat7C+oQ
TKTNRQ4FAMKOy9qDIQI1qWtfTWbP5MPJ6UZjvZu957KPy/bgOV6XRCIWKc8x+f88
YrPl/NkwuIAxh7gZ+tAkqPlv32Im639eu67ZR+QPXK6v2jBiOpbS6Fnr27g3EsGK
SAAo9PYamVbgtz2PwiG0RAQXFyvTJZ98nbwRbH65+jGCSGMsRv7QtbkkXqSojYhj
h8FM1HW6UuDlJ/LSwWBsqhApp/XWQEzgFXfN2RFOUwmz8fCpVbmBK7qhDg38d3Xn
m7bB0IBjtGnD5AYw126x9F0A9FbN6EDwZrD/g/ZOhMGEsJ7Xlo2F+wPDvelZt3qX
lHSM65QJHwtMtmi+xJnPLcnaA+GUXt8cXa29OyR2CKnz/OPBDOvOG4WJHhgUPRZC
MGWheIAjUwNPk4mPQD8GjSUsugksbRnSDo4GMUELQL+4n+Q0AibHRNZ68OOyfnnc
3m0EyXpOU/t/ydaWC5uKzPyRy8ZIH/0nuookQHkAnc78Au6MyZv9b2dX4nM5SrPq
2XH+8Sp8Ry+nROVOcdVb8uLuOXTUhN39pR1bsmov2glwhCl62q9I3y4FKZumt81y
92w05uIBbiTQqhQkAsl3FhpZor4U8vo8v/tNI+6sy94QEX1BD4bGgEtKnnjESLL8
fedEGJ1EIXlKk1WYtFYa+jkv/HO4nOUGjPe2HqXpX6Hx8W2k6GGFDI6pWRmGLRmB
P9w90uYAQXZqMCCSudcPHehnK4dwQrEyhVFdxXkmLpPZcMfKMzy3nDXreFvCzuGp
yCkM5rZYh+TPkhETDQRcVPipU19690oW3ywrw8ilPt0GTMi9Voh0aTlVqfNDc4rF
`protect END_PROTECTED

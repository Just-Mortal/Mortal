`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nmcefIJcqRxt6/m5mJMh3dIWTIC6LcPZVXf6E0VARBe3uNHPvEvs+EezDrNsgIJm
9GZARAKlfJNoSc6xtV0twrOm2W2xcWTgKpxIStT2i7Vw5QI9aw4azdsuF387qI3G
cBz8TiVLTFPjkkr1Y4wtMUo1xfbRB5pgDsueZhjjFKtYl8PGjVh6eDbP7aOoVv8u
NobrKMnC1qdbnWTUG/7l7dQ6UOiwn/H3DoqEYMTmvJll98qx3sUf0LA+sBIqzC4H
1OE4lfS+1PP95WoPY8nJZTnpmRfRppT2uCcOa9QVUxJgvmph4L0sagA7i5iqBaR3
NWdL2eFHF+GC7XykMW0RGm1znjT4fuJwioFH7ojqXi6+EF1fzwjwrueP1lPFDKeM
0nrf6yFzqWIJlpBskGuwEaLTdov+eOi76Gq2W12Bl9uasnzKEEzbz38miSy7BUVz
kIhRK3KrhNTbo7GlihYXseXTbSFIPj2k+TnMeFb2dMn87vaERIWR5hCzco0xxi7f
t32gxwM3gOYrZVUD7PoYTKEQ4ogEBhkN2VjP5J7gqsUeJ/LVXOA6AT3+NINrIeZd
JCAmsVxQYmz8axaybayJQpPV5N9nF+g3HhXuEhfpamFh/1+tAgeu2z63sSuUKnWQ
NRbZezY0ETptRQ6ByrvSrA4bX2iBcDH2GxJ7PvL52N34jcxrznhxb4/MHhJrAK7b
Orae8XsRJMvrEm/MCxcx/HhtiTrNXxk29MlqfA9QCRE=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zoery5IZlQdV1oLCR4zz9RpoR5HnIKyCnFQmJcErNLH8GDB3IgDkH2uCBONbFAxN
UVHLltEO9VubwJYdIYsPeQ3k8M7iU0lRLocVmq3yXJudfcrhQNMZno1RLj0sDPQA
EDQCLvX/r1JHBFuFSrDVtbbnHKClbKZ/wmzBMFBDQLmmISlmjA0vrYpsNmITHd5l
L6SDIeaSHodaJdYRUakB5NC6tShZMAt9VTPPRbFd7gtitGce7KQ4d2HML+o8bRtE
eH/MXc65N8xf85rIqqIJty9kYwCsTV+0nKAIqWkU7VQcaQzn4DInfICByystG12d
dNCueIMPRDCwyvCxRaCV5qW6WUmMwICQ9RMCDjG/9ZUNKqtYKZ0YyrgROsY3Un08
XRG0uhQadSXOXS7iX5BSvukZy+4Yp1h+Oji7+uk7bluAXmm3ybxTNOYPkZltw7h2
ZHqzr/KAaU0w5mnL7CvMBnSQbWlVKgtYlmjlJ9FhOXKD6hBI1wPxJ+vAqbAQfuJF
4c8CRw2NH3JkQiB2e18hA5FBRPdaQd+fqM8wpo1tRcqRP8/FF5pnRO0iRWE6SmfT
QGJkiTu2r6iBFztn1GHp/wRIL7MfanW89H/162RNiITAuMEdsGDqAow53fai4PXM
k6+dtzs2gxPilmVyN5q7UWlRYataxjoUKeXPdGp8lUJpkio2tes1Xuj1GWTYG8Go
MDjEPb/HqE6GV6lgRc1cxqsIXvmt0553Y6qBOlhI+zk=
`protect END_PROTECTED

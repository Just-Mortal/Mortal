`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MN+B0abtJvuqkLVdcmspUsNgdZLBTNvpx03foWdRxY4S6Us51LcD0ILgjyoomjAC
0uaLDSnMJh0DqS+aUQFvSgdz5opWEQErHo2e/9nwk+4lnLTBY0oDiFoSCq0DoSjr
HstsBUoIXTkdZbfbnzLH1bduhFJ8kmeGMsmXXhHXjUhDJLTLP9kCfy1eRJpdZF3K
URH3S9XsjR1tRQwDy6VoaF+9I2U1YP/5dFJR+QXgX1E9rjMKOLQNIKy/Z4Q6AiGV
ye3ag0bju9d5seRZNhwj8+wjKTYyhhR1YiAdYI7Q35qUOo2IsldrxlqwQv/qmxAH
mFRVfPR6D9jxw8mtQY3e8oqmaLoqC9H5pGCkc+FdLxt4felrTfq/UYWPeeF/Q94Y
le4DF0kY38wIB0jxzs26VelayV0X8NBb5nakACqjAE1JLUYsrAORD4zltItU6rbQ
NBnrcbqVf84O6i/TO5v4ft0ijlkdD3GW2Ybc49iyVb5f4RvN2xFKhCr0U9ltZkiQ
zVdEGaVrf7B0l9NLycgqvNI4Dfq8b5Egg5nyVEAtrN1+B1nFxJC6SgizzE1fPYNB
C3YJePKUS/7Yic22uxzFVWQLZ5wg4omiNjSjKsbF6vTcPUUJeaANOSg6TBP/z3JQ
uuJ4K9zn0fCB0a7FgXo3IA9AEFP+anW5a1MGpqKxRUet/nOcF7qIIJf6AoegDX7c
0Ijkfpvd29GECPeRcqYn5viX5QJhiW6NGqnAImzJiqeRckxa5zww/USk22NCMpuJ
/xAakTlLChpao1MKNx69BiXeebXZFbPYayllOSltNNY4Hq8AwQYMt/6KCuOZGTun
qKikxF0OazjUago7mihYXBTcC5H25BDOp2Bz2vpU8iBBtETJ3HIxGmi6SnjVwY3c
OxlmyHTQG4T3QG4j01QPHdzspvDFTMDJvaH9nrk3bjKeRlgAzfPPrLX303HdLElE
HOlI03CGaakQeJZzyXvDeOG5u/Uy97yDho3wV6rnMyGvqW0PBeXag5W1WBPDaKyv
o4ua71dP948MuFag0KJr9H0c5W8qFUdl7LbBIEW4hhtRUfQWUaNKJU8TuaPya01S
wS66y7GE/5MOgvUGUXnoHA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+8eNrMIw5V6Cqwf2Pls8eGKnUMOPdna+HDlkokaUy4eAp5IzxL3KEfPOogXcHLI
d5FRDlnuD5pJ0Su3FpFo4YYbkYjk53gSrw+GdMFpU9XVflqfUc8QPwK/qnFOKsdU
P10/4GJ/m/tz7t2d1nLv1EgPBgvp9Kss4VXQdSyb7KqoSBwPGF5bhyo+qhlssQ21
jBGqa4oZ1hNlNW50U9vftMcWFn4P6v+20Xzn4jTg9Zot4Vzzx9obDnhW2Jm39Rrp
8VLBHzB5OK+Q0sijwf+NHSQbPNt9654LuZ46D5POOm6cEg1Du6y96pzINPtpnzE4
3kdI2mlbYWvB5y6VRxvOiU2iiI21EvNKFpxw28bgDE26bh7t+ph8+kZSkpeFZ9eL
IY8aSXiF1k7EP71QwYGH1YZPFS7vJzNmfji4niAarRoIh0Qj75TFYPj1hnlEyZ94
U3gEbD07x0DbJx5OdYweqT7Sv24T8NCP7jZYz0kvewbxTF5OPt1u8tMRi01C2Gc0
0Co5qCgP123wh01Wvb3d/HKDI+xePEQh50acDtMe+kFkPDgXv4PIrqBCXbqQthiM
H2RtGd9I390473eAmDzBr4uwcmYiVqgLiX5/73kkH7oEzC0NgetMCf251RC1cPBp
lm64yJQP+1ZYBiEnHz5OaZRsETfylbxiKtSPL9tJZPytruIetnvjrEqZCwIR2hHD
MMWUYp/sk19nlZr1sR+K0dts2GqnRZm/dxg99/wja6F5U4YNSmKaQHKmh8aE3TFV
ZicNK+jo9T/1cZMR2mF5xmKfwmU1y9LYOcFeC4FrHqpzmH3Cp+yfJ4cLNrydiFAH
NEcx045XIhi3bI/xO+c4wvc9zPq7B7IGqggMFyMBZz9sDXMvliRJf8vv8euwpr5K
jeb9pSp5zqwNME1lgKokHsLUQ/+x0z9DoWOxtfkgqR26Jp2xqoKrdFkr8ys+6+Dw
X6oX4EMfGBqBXydHA/RehpkrlqlnI2EebsafJ1J3TPXr6dlF4JsWbPpME/mRIKQC
/Y9DtmDOCiVDNUCJHuQ7/+JCi3WKGuoqiRrwVnW7HV3VH/NxeC8h6pRvTRBDp2WA
bCBTkaojIjMSbtAGBkILkEMqRK4c9Sc+inVBiE/D2E50ksJPEr3AvvTQvFKAGGT/
xkE0ytcd2Pw2t8NkOjo+runlg+XSG+F1hTLulFnlMiYXt8lm5thH9yaKrB3TW6CM
ztjImoRmytne1qDlwBjzXxsdqXOsbgk7KOwE3LP2eHlG71E0awf7QasEv3o0DVnR
HxZ1SQmz+1HcrvU7r4lFFYYwA28mzgvtdmpY3hHawOUj2Pe0uaI91/ullHKvgVgL
g98IuRz2EurW5rDvOCW1pAaCPpoTpNcRQr6IXaKrz2Feis9wBwOwNNzeYhH0tVLD
t1JF1xabx1n0kL7wcmO1zqv0Ag28fRjXsedxJZEj3IZebvAzmQ0bHN3LzcQAGd3K
/WMzxTzh/xiuhGBjaUTW7P0eqMZ1V/Zix12x4arfGiNCjr0Tgh5hBP66EyntSdt/
LYytrW48HR41VRZjG3/Y85x6gh156cLY+seA1ArD6NMwo4EStrNuL8TpdoHSSr9t
zqO7TW4v6Lktvzw/XTvW5dmtx8RlACBFgi7QSMwmDaW/wSNpXwh57KIP9ER6f1QH
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8pg6roOj0TCA/DfNzaK0GcV7nA7NdVCyCvZV6JfPHfPyeYq6SCyq0kRgcxr7u7W
UNhwTEdTMDYdb3o2DWJUa6Jh5CkRkKqDLsnbYxuMJbNCzsC2/IXZ+1sNqNYLFL76
n6VUThWDsGrs9e9CJZU9U8SqCerLgwrFU1CN06ksiHzndiJeYOWBywb57jvUDsTI
XRlNJYHnkERbUj3TjltGeWNBfCm9h2JyoBMetgiFHbUuYSZxeRqvVxUov17avj8b
pNHd7nDFl3pxlYx1e1u87NAS2jLIxHMZ/AC1G8od97HasRcxu9SRZo9zXvN3RuOY
EKnC+BxaSwEk6MWYaU9cZ+QBCczEdDJSdoIVc13fMFvJaNJkPHGmt0LsKrRlLEG8
Roy527S8jJWOjgikzQFpjjbQlB5+YdCpdUHZ9pYrsXm23I03yv7JRpqC0DS1UxoF
d85F9xgh2UvazoTwC7DLKDS1QTPeyUC/zsY0x+FsqmTO9f05gGN3vXbmI5uTUOB3
k5mDRwWU64F7wTlyIzdJ4cEPeeSfbDMVGuKmVfcjFAg=
`protect END_PROTECTED

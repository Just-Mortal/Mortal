`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zj0ROMjXpYBjxrVuR+HeCkHeDwI/vulUN5xpMcGEraVIKr2M6YIwoDPDFiYwQ0K7
Lg7ov6G8AfmnEPGodrtYkd6TT2l1YBkRLDneyHjv3R/I/VLBOcximLEybCsf4gue
eQdPpP3hVDMz4aj1TdfpS3BnV+gdGbKSqZx8XTIVHg1peG9bO6ek2KnYAkB2zjp5
hO8ErkQoTPrtqaMf3Fj62ITxPe7MEN4l5WVFjDKNhhVcYn0G3Noj7zSUMRJg4kZs
d5EaSJGYWgd14hrmyBdI8CEdJMIw5qtGtwNH0a5mhNL7DeAforyOoFeP9XNaG6ee
28nBLrGd2yTsiKTuAcoGXD9wiyZ1D1OogMFjILaY2YGxDmAj7K9Vs4+cenStdvYA
7YSYTYLPyOiroacCg2N7YsAjh2K/BSKzqgtmQe7/N/lCVxh20JrMjHVhf1+FC/fY
HGvuexzO+IW+PpV0/oUhcO4AIBtxIYXG9+9yQ7526BhALYJwAtT7IrQ4ySgfbqQs
gFz1lxXdEuqhm+ZHpwmh2Mes0iTdUb88cxK5l2SvWwI/t/xBCGS9Y2FABgIFw7wz
mecwW27Kupg6gA5SxhT2EqFcIdM4422+w61dP1dBjgQVrDHzLh1bS9OLpdkgW/Zt
jWkHkN5R89DIs5xtrj1Qs12SFMKdpi4lr4FLk1mTWDN4t1ggfY6n3MvJmJODIq7j
IRThqd3kKHn3Bk38F4OatRVSXGddP2g0ef71Ls8PfFSy4Fn7S9B+ZC4esboPiK1M
E7VhKX8PdFQ6KiL9OoeH0BwM/176CmjUHpRr2hTb5n+IyIHPMCVqVoEEIFxeHgUp
uu/IigQKQSTslbTsedMm93eoUEijz5qtAZ1TXsTCgZxOGwfSWqFcyCM48Sd+GNFx
zPDqX2piRuWozDxiQmfZ4cah2AiU+pijv8qnD5aQlsUbrYRgCXT9AL6dSaKoKCCJ
u0xxwRuxSZf8wcqgBMfs79IZ2NVdGT5ORRhh0mAlWqPxlHpebCa28HIfp/7msSYU
FWN69VDrOMnKMI6k4+yU6QRJTmHCAvDcDc89ATE49rv2smUjYPg/WltOljWyAez6
gkb9HIjUllEPbodlq9wplkhlJIRZyJAuSdFjcIabfFga1EVaVIfFgarVwxCG3zFS
HOzcuxIi2S70Ak3stG+ke4NDdeXV4H6eq2nx0LiJbhGQ/2Xy1HOrbmU+Hte8OeHu
BZ/dzldTN7nK3GaAWXm6uWTgmgfOPEYRReQ+QcIzITAq5cH3z/zijzSALsosXrWT
b4ZozvGIoQk1NYP99PNiAj3VpISdsZMe2HmQGFtw4KOD+fYOasABFfNF3Yb0unit
Ub5YNzRzBqSCj9TWwE2CA3dAO6j7dEFwl/ESeZmM8Kk9jFZQibNwSQ+uF6Wj+J0F
BncWlWP/cGDBXTJ8K+QBxBgSV7gqsjJSOANd2CFoQAkvORYi63ckIlRCBSHMOE4J
iIYaFL1r3KGbaVNi346U60zq0QBzPo82z8g1hfygT6R19LBWgXLfn2AgmvvsTkky
mPAJkhPD5ceu2G9JU9egenbQbmwG+5+ZNv/ulS1gwRZlW9SX2yLmM0vu5fyNKHTx
ARQ8Tsn0uhK7VmYZJ8rdz2Iz0W2e1sW6ftrmK7Wx78mQn46UCq9fEi4Xa/C2/vvz
V9QtQlLMpdprkWokkVlChIACi/3ceNcifjO56PcGHOF+IiO9C7XuAF0UUFsnJoAy
IyGGgsUR6v6uf67vyEfqA1nUg75BqUgV89rqTeFI8q/pnxNcxa5biHNRa6q+2m/r
Yb4G4MGUDvYKJVREqpV/r9V5fZS1lrXrlGvpdGKBmpC1eClve9DIWrwY9riwk/Sz
t2r/dBRcXXonwAvvf9Txm0AE+ucm7e9Lbe+t2EU6Tm0HlSMvNDYKGtABJUZ3iKoh
gNEaIA6H5RXtd6F8BtQuyLcHP79r3knumFZqf3UaE7mVAesBRlD3xRsZJReGG2Lb
3cKEFjQdzAwuZNDMgftVJqx+myVMIOANoQTW3AIZv8bRbzg2tvICHdbpocwckbOi
NF3sDTtov21hdfnjpMCEOxLC/Zx6m5sTUWZyXO8NfwoDRCkzfuHbOBbe4SULl/7h
BCG6f2D8F/KvTTaP/lpsqufcKEvvVOdIiDR8V01GkutNhsRGxKjV5F2qcLKhJ4oG
Ill4aK5QzQx+yvLha0uQGBqw5vaZD3G+xQaS0g4KnkYcrCAJjUlgY645ub1Il+0r
hw9csyEVZRadU5zFQAF/i5D+sz8jTsdt3UsdMgCgRQEx5Jn3L/CmHH32XXQxJjHg
M9nJ4dSQhaNo8gjH27hQdoUyZ/GU0l6hvCUGpOTCmS+70Mw1KwQUvp5BG+KZC8RE
rEOs1C9km3JCkeONLwPAFQO77Em5U9Z3VkAqYiGnlHmyQmAwo2tflJSMG7I8wI4j
UlhN5kN1kb5ewShvD2dEZO+dW3UY88jXGt5rjoWyyFkxdSSUt2Emmrh4k6gHcFhQ
cGBaOdYobKbYrLgILl4ndsjhN9KISq7n/S3Q08saaDLq1B0ZakNk89AuUgc00vu5
dwJX4XfqkDLYqx5rCQTkjIlXUfr5pQ92PUb/QML+DVQKE6Ktb13PiIRyInLWczOU
V8N5vKrolkJ5irCHMqItrKNJ+Y0RDdXNn3NxVQ9UYwaslhnWUaDFiBCgFUpH9J9V
UfsMUHjBCBEKp8uIoGIIgfmSVd2le0JUdtll/WVmdBEIZHOfgs/EA6RbHl+rYTs7
hmYf+qTYbEV0Q25IzifNU5W9l9sreBq/kzizme9ByzMyiQB6D54ooKn63Fawt+A+
P1xuj+/mb5P2k6Omln4H7AOqtpt4yYvujwT2TNjRBAOnwRzUQbUjtuhjabVtKgY7
56Nn6lzMAoqblg74mLTSD5cGU4KuqLwkWA4sSv2etPeATfzYAd++9PvTSgkyLv9G
Mh4T4KvtLY7hsc5Sa2F5c+b81k62fpT/JPNRPZ7KeTK8A/vNDLVMiT2Sqg4XRrm/
ktZGx5sJ/dT1Fa83ep55y3cA6VQ8ncaqfqG4SWwoKu03N7dtgoNpOFulgpMIMXJM
XKsdu4cns6+qWVWR3eL3HdZl88nkfrUu8S5rEcB4JF2Z1+75rFEJoMl8LghLkVud
6nIQGa4IeZIv50ocegjPgITLZCiGSJJIsV2IodbIfJmhUzpXerS29hMQ6FpEs65a
RsG/Co88/kbv3sPMUlqqtiCPCmJxkmPkJAHlL4LaVbzXpb2UssYV9Dbi5BhCSGoI
936jSAPX2F4JvDJMctPix3Cr69aPMUqf/StQV4de5NU7rBNuRg15o9uJDsumLMxo
N4o7FHW/lAvfQ143vYXhA3R+sHHfLI3IexlSsctzZagSWUIHgG2Nfr0vel7hxCh0
MfS7Vub9HFVJo+QK6j3tjU3CV/I9dz6X8SS398lLI8LmbjZ6ozyKpJLQi03lonut
Kq5gBdmf3hN7VwJsfyyhB8lSBQiMD0yotYPUGVgLM50prcgQzQeLrE+bKlyfX31n
AcvQBDEkCoORWxgosWCz27Orm7T3Pf8SkXEWG6Cqk4LdMexYjfs2HuGoTKvH8AfP
jtGVJHLzq8OVWJzRNsbK2WV1fgsv42JRxswJAoHEWHXyPBCpYeY5kw0bdgPxidRt
mDuzQMVYtjB1bqEai/oJiA3ex6u9jo4A2adTx4sX4QcFQtkwkJ4lChR2fnMn7iaZ
NfmcYsx3yfii45tkGBIc94iy5DVmjGSqjSh9cxbODON9Bm/7XGa6WrpZH+oyjEcF
y8tB8Y5yrFkHBz/hxCje+H06qrWbbez+V+Ejqq1cu1bBUOEOm2UPBMwfIuksT5PT
6691eEfYgvGx26gZejI0iRqbzCYUCZQDrs01G2Mot7Fybq44g7z4SsQQkSMKLncC
HPUu+MqC0pF9UltXj+Xgo0o+/RpbOs6ResgP4A+G5asMp87ktbFTzwnuxg/hs6OD
US0zaPwaUN6Cqlyni1c801puEWvnpIlsddJ9Tf7zmPKtmh4VK8sjY39DzQoZRnok
vcS0SSev+M5m/wPKpl7v5E60ocaHas1BfUsKnvkIfF5DB7nK2dzfxdg9uqSF48Oi
i5+AILAMMY05lhDM2jjmg/DlhjUcrhQnl74TlXFp53xOFPk+VMsHnJfpES3GZQk3
yDA9iAvn5lBP6Ej1E4cOyK5UCdW7aTTM2eqq8KJ+BWaTO+B0llUr+j8/aTVYPvPm
ias2zJwOuIytPyf0SZmQX8hJs6eOJhOJqnrXwDbtWb1xZc/iA5lfvo9O+7D/IdvJ
zgS2ACvnhVqNwcwmiVX/0D0UOJhYvNwN5CwFYJKIbqK/vSfxnk0+Z/6ojriiPMlT
JClrs3ouMEUz4p5b+HtqaG83i4D++KLfL4im+6UkMWSDoWw3RCJnaJCO7al+ITu+
Fv9xp6Hz3pjZbxHKxwZhYX2/IcG8TsPNR39JQNYCyV9HP7IHCDIQv/2Z4u+dY/kc
oJPDMVAUhlpRzPmKUz0N1zeQnKmv04imvpWaveDMrqggt/aEMTDxJRzb5jbNS15x
+VCMstRxaM3PFV2Ao5IGxh5XmrWQ3QpU7+AJLD3nA3Iei4aM0TVbdGrKrsk/0EqU
/80s11bOw/HBnpdEY4HMDprqFRCzeqYIF/5NoeB/SU0IOIvE6bTnRivmehRlMbcW
wM2KKWIItyAMNhLdOY3VlIj+YN7QR9pIJMPWYFyzhnw6T3RntUn0pexbFWsZFAG+
2yDFMKUlCgDM6krpbwyxeMTkdRC09D0VEGQMKDZ9rIIUUPDkX2lPRCoxOtPvC2iE
N3uiRHENDnOLZWbA7Pd7LB/5WQPMsD7Ea4/44N7+bXcuiF+VSSI3gMeTha/kb1jP
Ac5QgAMcmPAZ/IDLXzcFDqdCeW94Upqy1wEnWXXX8dkCZCwZA33ywEGvrdye3JYQ
NVIE4AVIzYC+Z6i78ZljBSNtwv8QnYLj8+qs6YnAj9wohHGQQpPvNebpQAN8ZGw5
v4B9A/hBnU+LgaCZlIxW16oVjF+giRF1nnwTGj+Z6pKobOOR2vlKsTHSSh09aR9n
RwQM1yzYVImfPG5c3LJL8FluYhXX5kVZ94zpyiYt5esspyGuqyzpffJ7PixDO3nG
8PDWyxshTYyN7Ko6ChyDevY0SKqb8GAvFg6t5nLp6Wgxk44qkiWi7PTw8aM2f7T2
QiAlxnbqUAfEhxxX7QcJB0Dm6h3jbHI2pH7tt54k2kL5zf392EYhTiimq8lS/qej
ZTWYHSswN1MkTPqZ3Ua/u48RZVN5GBZtBcSciJtS/BTEKcwR4cZ1MOBk0LB86U5r
7I6K6lWZR+i8GQUZ2OboP9o7faP99pl5S3xmMVJgimFkyWbwWKQRVS+r7euJQ4+n
i3ajKrqzE9nXS1hTvjxKu278bWFr+tkSm7U2cWPbzqzYr4cgnq6SYkxrHvGLm+gi
N0823cmZat8NHRuA4mJbNiI7PsfJKpOeqAAHHZa0rSXGe0wZ34wbDwO/fEZ1/4p1
Ypy4r7+Jn+mqloSyEIdzjHSsqZGGxHgUcB9yJcfvVDfkxGOGUXX/V2zGtQg81XE+
Desn03whsBujDYaoauryBg+LzobAO71MeD766Sm9nU7+CYz8onDl+aa8RAIncd/A
jE8sfViR2PNSDLojNnCFeIgpXDwY/ekpdMbuetkiXoIMWpbZn+si6lSdmjKkTJH9
cDPUKzfr4/QZXPoyQ7ZyRpuxZtJnT6GqLkTlQbp0598KH4Ad00kiKNA1feTBobYl
i60iXjpmfLB7gtwQO0fcQwkZurK+Y9pupK8LBZ+f1j1AGjS0noWClOKMss+HKuRX
4TJKGiUmIsIqmDf41cAaRbume4VLMKN2Wk3bvg39jgfI50LqHecGBOG4/mUMIo+5
fk+64qXnejFXgtqcqe9OL1iICeKslqKdGLPn09KE9TqXTGaXWCt9Edoq5dsTke5A
mSKc6JXjaAkbazpHZqVJbUxB+D4SemG23FDF5R+Oe7CjGsuoTcwHC/JyWVNJXvt9
x3byoxdT42jBhzviNla9HfUlnn6bs43fOjiSEHknUqcqEyalOpCmTU2sKLZCYJUk
qHavw+XsSxHLTD8hxp8bk2sq6z1IURjkkwY0HgpfEryLtzWmVTfqtaZQ/PI5EP17
UdX1toBO8F4Vr2nwJ4msffQTwonQOjDXG49BkganGv64W4aD4WazAzCYD/GdHb9u
KunOxGGheK3K3j9t0uAlo+tQ9JCt5xvcIemA4Gj/Qcueu+eHzMNAGnBRtnwmDb1y
IvRnhKwVbqDLvxgL5M3T5V9umcqjrXYDd4ZjVjLMTV3eSbIQJPMfWrPVtmIsyNPk
wxYcSFzaMx2DNGP5OenJx9kDHtj4jD4p/E5g1LkIlrNfsHtd+K7jZeTYh3cRLcIQ
UKMfaB6QB+2eIAuzG7RP9DkOsLWal76ly1uVqbxcBmVbFnI4tU7qbytaNADNg6EE
Uu5oasoIoqRqY4VEXnIGHK/aZfLdlYlZuEAKrzovrepHTJKAm8KQXSXeWTq5i74+
nwt2xf0fyYjXiAAbklbQrrT5FJ4rTaEBblLhJS4VTEMdOmlIj/dQeejGMT9R+D7p
W/JKm9BtPBiM46r+JbF1dgO86YlHWbdPGC3KP500m8DVgiOic+rknCc4yqRY6E8K
kRXk3gKrcs+VeX5lFZ9WdnrW5rDbc1Xn+K3oS16bATY8Rz5djuJZHjQi6M23zi3w
iHACGj14Xg5SNkDp2Wu7S0TyknpM5jibbyIpdB8Qn9CVAv/5PZ60pxA7Ra+nphna
LJPFEKQvi3BxKoCD19Wz/Q/xAhCfAmBEDfuuJah5Zx0DYhGmIlAN90V2iUcrslEF
BO2QEYKVOeZOnfuHhh3aWleqOOFdRQ/RJ3sffslxRjWRAHXIKRWI9+NuqSCfnt/I
VoFBobwErE56z3033vYfRtSEQr7dX4wOh47EXEoXGWXeRcZr70XAs8kIkpe/6BgI
4YNUR30eKvJB8DVWjZqPwt8Q23jXIR2b3YgJG0Z6Lv7J+HQVvLcL96d4MHrUH/6T
e9JCES07QlFInj56ZH3CwEc6B14vJSb+Ap9NHrbesexJUz9PVbQQCR3ghdxAtqT4
wLGhOv6A338Jo8fcVPWmyM7pLPeChm/O7WrYQutbKddRPNRW1AT4q6XhIiODPAgZ
TQfvGurYM4FBebJglTQsjExxsyAVdxCxBULd1TqXpMKAhb2d5v+d6y9lAsgEaXpI
unsfWz1SG1LhlqqrG/lu9YXq/ZsZtifTdlKDpVKn8Bx1L1tUFxqsWBPNBBkAIWIZ
MR6fP//Lisx/MGgMgK4y61Cox8W6Bi/agj/CzviuqAZAxukNcH3TzjNDu1nQpLjX
TdZA10fbKQspYIlnljRg/re4DJoWqN3xFHehwqZ2A/s2FmUD9XlcctX5I6rxyQz1
W3RjZRR5PkQX+m6cwd6WJcU9rwvhAxds+wnI7oLNi2a4a1sV3ldlupvOZ5vGxOXp
oa3zVjcVUXzIi1/PejfUCknSiWoTKxYR0c7mQ/6o1dtH3UDHvgqH20e/2VAbiYGY
hs5njA5KBDvz6lrGP25cqtuqWrnTEq7X7irHKtUNp1zXg+m9h4wEhh/FrQiJJhEo
EYtGXjvkuLyKXFX4s14xzk3d/wXAtOtqtyYOkE5j3O6H6GU4cAFxu26HJ7gu36iW
pGhNG2y35rKhlOBFCy1gWeoNcaR5gHQ/lu9/TQpGfApTwHaVNbLxTEOzGLtsvNyp
fI6lgXz78pUgs2fYXN7NdxtQ+Un/DUyPrdaQcER+d2EsD/3XsWAI992NFAbW+499
PkkYNPyA3MPa6Cp4uETuDoJrzma5RynBhNlxFLQ425lH0mwhrQCi8IUBO7dtlFsY
W0wxDm9IP1/BDVLOATQLLDcc8GblHyQqrW0qDY7TxV4ipeM3m47ZxK3JVI8jadlZ
tObYN6ohxRZzBygkCIXq15WCgfoLY3unJi8JsfcpUIiQKYrdElKVCOdwTEm36a9o
1vGHpMgyCqY/ZrJZmmvvdXJASFAzzERUWoRn5bgFw6x3a+NgBpk3RRfcJj2R4TEX
zYwTXeolvDavULutlT2ftnie0vebGC1vG9bKtyNIrCzNqGJJp6QNTed7rV26iw2O
anY+HwjGQPFbJJuQDGLU1eMO3Xtnv57i+tysaT1FqYQIX4QvH0sDjPOBqRrJBBxi
ipd9Xd6qS2edajPJ3sz5Z3WHG69HiEuA50j386uShpn/KowbSfol4ifW6C7Pliov
/lJ3Hfsoj3PHWkWpN1ljY6gkVQGXf6KhJSW7rTz0uVqfJl8gwA+HM5l2rBePC+1i
+ny1KNe4OLrIvykX25DB77TT/0lqmS6GOKy7dnAvuJdJUruTc0IcvO1VP0obS9yx
kmYGtXfaPq2m3VqUq5aJbJmQCiR9bUDihUBsLqnvRWaCwH6qulZPvyQXHKvHUegs
up3EyxzNeOB7XSTcfSzfSYy1ifwV3bTeIQE3RVNB0ntWe2f0DE2bwMlqryBcvwpC
TLSb+F3QfHjUe4hyKYUynvBEV62BoRtYzzutN5wHQidAvZdCC5SujvBvy9XyQfUC
kJYl4IsdLeXguI569M6bh3jXWnNVafCDfgWdiS1/8OO/TMN7sdYIh6jLYdECMNHj
4dJiD+3Gev0dXVtAJZ+YXDFaDEX6H4CtgWPWtSBIXgDoBD5ximnaVCkUfJemp386
7IJt80q1SmFU+iKolxxtzB7SR69e2aE8oGeJUgIUy4Ku60/0CKoA83S3cFGbCYlH
pGSOkpH63JJ0k6Y6N42cP4UH7LtZQKhUwzWOBHmWpHVJT6djwKMKSARhvwu69rHc
SwYXZz+Hb/NfpIXNgz3mTa/i2XgeEAQ8rv2XinDgG+Uet6y5ItQ6b9sUZBqnYNFJ
bjnO3U+bQPCmkTEeh3pT3niIJdy8Ow/oSY8aXWq+C7WCzY9qZhL3LqbOIHPzhYrP
qyggjjRcBnfEzMnFX4RF8QiMVm1EjPsdqchs4ezi46O0guVt1Uy0a+h4wB+tHs0q
MGDmpitL1LSHA0TyVi6JfISy1vtmPFTJCSUDoi/JLNyAf6OHrDsNSR1zE180tMG/
DUHwqha2JJPsaauMMkOYOTxGzpA6lj5aNix8Wlr16CsN91oHa5MYN3pmsBV65zlV
Yq8kUb8ZL76/c8Qi4PVAZA9eOD7p3W46rw23Rqo+Mb9zVYjxDxVNXQW+aTOBKXXH
vr4FbNjXbPLbwU8BIls9yfHEhcwiDlR8kYdbVtcqvhgmhIho+BkS+8EkRD6EekpX
BgvcDBNbJbxla7UtJVtgQR5mW6+vSJsnymuy9rm/1Anh2SjO7DCH/HHEEDI462Lu
tZEZ59PU8vLR+9gKm7kyreTF3ghk5qxAHyLKHeFlA9DvlTi3LQUJimc6HpKhUSYy
VV8bZ000lTOhf9J3vmZ3I97N63VkU6jhPK+o6h0WUqnqhTrNf+QmXGOFuhqtiy+0
zew+ZOL+Fys/46Tff0Nt5lDXfUDrd+vEir1uzMe4xC6A/Nzy+NOxezTm+Xvp6XhV
zzXf1D7bxgJXBO/2EX0bxN2DsslyB1AeJg5jjg1tZ1K3JLhv2JPrj4f7ot/Q++ny
+YKi5toYKbGi++iIyi2vXbXn32Y29XHPbOpzpyLOd65Q0jX4b8867sbJe4gVj9S3
ygq/vpyikOfsOPrOvgZVCwjYbwEu0xXIXVoZgg5etxNx1vGM/qbU1pDD27IaGpIm
qbifmEw6MZbG5Fk+NBQ15XfjxaWVVAaoKrgRVSgX9eRJqXU8SBENpIldWa4JWT/H
5w4L1IACtvWDnjjSHxU3ddq8F8rlQLpyWTcHsDU9/owLx7JZiOc7cdAZlvq7kjZD
DPpol8EzWWALgw6ob+dQLEabMuwydIbqpyn69uKXITzGpeZbgPqdQJPEC1bnzTGd
YboOa4zEf/ZiSnX/po1V8jaXFnFcMDVqg42BNBTC/385dMR/JfFOSfCRTiCkvpaD
bNQ9E8knN2NUvwMNAhmch1FAIuQLpPhaZzjc1JaTAdAQfDL898y87xxFLOUJwEwI
P58Ofa5TFGEeTDDurMaXMH2tbLyVnXd4MvINzIh4RdGPGN4zicM58qwD/yp4J2ji
7kTihccwurgdBpk+0vi3kSSN38L2ivCfgbXoe+7G46EbaoqzhAHPOwpwE2x6weD1
AbU2W6wTztgQuQ0uUo6RAKctnZdZmM7JFVd0CdhialeRTj5mkyKYQ/cvxdxPQK/f
/LlsFOMqMMqFqCOZxuXiuadwncNYudJ5WYGe5WBfEkiIfGgLbQc7zQAfuH8gZnmn
f4sbdKhnQ3CbojU6p2G2f4zafVtMWfaH9nqUV9ZKSW48xd06r03SB8qVVyDpihtO
fxPj+B/O13ACIOVmaFhcPk2qO7yAQ4o58aFmT3Bfrd4fjI/EksLQfzLUbEsbM5AR
Ev3oxSWEA99Xc9o3dbntTXIcpbBTVqlU5UWExoxljQoTQd6pBanyduKlu2ICCFR2
h3EBKIH8GBzlWe9MF041gk14vky09sKuKF0dlDSvbmjwTigN7S9BzEzPxPV8NiwX
Q4a2XNkUiA6GXLefCFHYddMeWITg91KfKyR7lbphS5jSroiVWdNxmrcfJaDpSunL
l5/BZruTeNwDt5jsKZd/d/a4WgGpP18LMxnbDb8P3WZeCbO7cUXYdpBVXw4aFaAt
S2HYdGYFHyIj96cXKo4TWgVR9MWUNT+Jo+L2I1WSTCWynLh0VYTjW4SM9EgM6asP
Qs7RMYUSRs65WzI1sqFYizD1j+PLUK65GeU767NyebAad9crM9CFPfNNaSdm5J2H
QN+9JgTo7fHBvRp2nwbsuDHhmerhCt9Qwkzekr3nDIWNxwyAjDt15aSZ9EP3pBqP
XlsgCclZLn28xeLIfa3xpyKpFgTXc4J3Kw3zahoqYobEUBojeUZLTXmZ9Z2LM8Uz
6pXVRSsPnVvpeYfRFeppzxoeudNd1/aEW6qXP4V/hAtxhefzMA+MkDsVfckZuk6w
YAP4ed01CK/16Nbb7+MAnttpxpHb3BvTqlyxo8ru020cl1r4VTZQMkBa5gs1SzV4
LXNI+MXmaMcJQ7PL7gD3KhUmYMINQl7QEa84R9wqIfoVRW5OunfmfO5UIzixts/f
VVz0hOiabbOgp5pLmU1ypnfseHhrgAdSt0znn/ugCLP+uBRlHpaxzrhtXz93dGX6
/+1PyiCUyhrGT0EiN/+K5e80IpEngCx/NM3eEiw8PYRj/DJ1577zrGQ7JA5v0N2W
ilXEBkOIjqlaX9tX865EA/43Pmcd/gbiAhi9yO/vU52oZnk/wasM1wRYQ4rWYfUQ
6AXcJSaToWy7O2bETYdrIWdw0pzWg8/VpIXQwr3NMni9yadsu72Azvjn+uyj6N2D
1zB4/0t1zOgQq4j2EeeEl0qYqlMsTzLbeBGGBjRYw990xL7G+X9ltHcbJpTwoglY
F2vhMNL9P6J/GHU4T7LEe397XM16GqtQ4aL3LtusFaZX1Y9hIUNp7Bz9SfkSRQHH
d/jrcaCg8vyC98CC0eSkGOeRgrseEn2ZrDQAHw6f/lxFgSdQYrIU269AStFB+qYs
YET5YtFqUAF5bcj2zTOrn5mdSkMxqeHKDiG5u+r+bU2LfZ3eqC0/QNEYUSWYqciQ
oISIycu+f8VChqA9gYz5qGEXxe+/+B7Mel2GnALTG+ltAJ4cAPDb4mvapCdmpMis
tYv2AcaFdeUlGDggw8aM0jJdOcHKeyZ1INwHt6WChWtsrgf9MleJElBq/4yIpCFc
Hzh3Cq3x2zZw9WefmU63lMhqolhNQ2WEHXiPMTsuvYPOXPPNrg7Uhsg+//xW1HxQ
0RES4sohI68gfkS1bcLr6a8jVXq7T3m03PwI2RoUgqLIUhnKKH8O2JhkHTdHvaxO
NaNFb+OVAXLhhPjiqR2k6kWt/2VDNaGg9U2PPw4GWdUgxKRDClvkOoFyYht7hm9N
4+6Ba/4pYGr6n9y5qzGflXiCktUvsi3vd0ubOmFBS1vg3Lkc2ceTqYjR4WCKZ3jJ
FPp8wAE2fIJd5XjhDMzwNVelFZaPVf5+sSUhcmuBnA6Q5A4agmeg3i2+T1WewLs1
NUJMBn4MREH0yej3UzV/eSUf9JXN0eE0crk2nM+0vQeiQnyn6li9MYg58zeW71qQ
+XyO0Lin6GJ0zB1mT3JE81oHgfMONIWYslqAwFw4KtHBuVWR2bIkXfGnJ7THE7QI
Z6Ct2I5C1V54kvWkYESuQ/lvjzPSyA661lnINWBw37acY2eWXprcFNdkBxP4glMl
IYRs94vqNdvE5uRnt4PDo/xvQ/UMeJQ+9O0obMdopCggzdfffhPaVvkAcfGJ/qBw
4hGy2PYPvdb/A5VTsECAoc+5UVSuNkq8VkQxgJi12PCJ80Xf4OX4nrr6yWigm+3V
YRlGhtGUOG0mTBkITMZuoKRTq7tKrnlOGBW3m/eoNMQk3oTAStejbShbtALt9KCd
NzWWsnXtb9ZHjIuDD51BbKSpAdlcBaHrNDkg2UKcRXn0jPXRyiNFq+8oS2tfIpn+
ojzOEhaaJEToIo1QjKa59SM381MPC4QGqDTBLt1ETix09BbPs2DnE7/hslFfPBbV
WDSO5vasY7EFyKpxPTvIb7kcWzKwqz6hFZK0DBUGo4NkZtAGiITQXGZwkqHdtxQJ
E1zkx5rbmDxAMu8M9It6cWOmtazlUUOarocChocnJQUelQosy393d76O8KDnJUw9
K7Uqok6vxkQQduTA+7+oWxXR20GC2atQdbaC3xFry3rwbh0kypqNCoGFd7ZeBGQm
OqezWywQwRMi9PGxCR38Sdh9UMdFNux5lzT7dTKT/9gT9mA+5MbKWyIOjOF+znoB
SfMLI7PJQRQ+c+vbVV4D8ETE+YceiyQnKbMn8KBC9gKlPfER0KF+WRTflEdiEh97
mUnKKSE/NHcx4I/mT98K2XJyVZ9/j0N757RiY+s4ZgkKkNzZDrdyuVIEPU9DPyU+
LvBB+3B+sHzVPw1NEHFJPug0h243E7ORliNVv0hbWmjOxwY3ZUsM4dlxvs2/yEYJ
9VUcwok4UIjt1VEXdHUARQ5/cW//UnsYXjn7We1zN2cozkYf6ERngUJNDDcx0yw0
JuZlFf0dtU5wYb0iJlNHeKL0F/n83/u5NhJVnrw7LJYiBYNFKKqU2+SHsOyXNFIz
a1S8Itbr0XyPp270z8YannA8hswjpRb7gFwWQAcDM22DZ41C2SxOcPaDgB5fRPob
uJmwa+FQBl9V/Un5Z2XfCjU0SlVjy67/m5iVFSgcZPPy+8oNc62t3OH38T5+o30I
zTcKkC1DrM8kxf3Y3H9Kt22R7XR63RXo7DcBGwOqYlUGh8nZdxw3wKyL+6CHv87L
aFMEVl/kJCN2dzaekoGXFig//m2Sh/xlwMqjUhqe0WEZqc8hvEl2RINV5pdgHfO7
IV5CUpPqItbHh38X3krlk7i6oNSeWDVmTeLKc+wZopZ9CNkTc5oMqWeN+cEOCRAr
qHGjlBETzE/UaTp8w8XmvWoL7nDK0VZ41OxYAHnCff754bOi5rZKSzMITBvUdOCk
dwnYUwBBfO1IIlN3UKchdOsrQW2OPro70Hv19FWNrEx24wcXAFMGU8AaSi6BZm3C
zREWEgbeRgalOTmB5w8AhcHjCB9qJxcBwFylN0vkm8wQRNHzvHI3XgZipAePBl0P
ciacxx2VUGr9KSHvZivvWluY5Op27+9MPhcM14rai2sAYHeu++zEt8FWzX7Jc3GJ
V6uLDCGcyajDf9+xIHw91B6TjWMR9XuQOLAbXvhfF6wj1LdT9Cc32iDx3UjLbt4H
PgME+KL9Kz7YldDKrn6qgw==
`protect END_PROTECTED

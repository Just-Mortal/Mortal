`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjFolo6OdgyRbO1DPs1nt/2v/MnhNCgIMwT1RTTDMLcGDBlSsw0QGriegGlbwYcO
IFPRWg/IhYnkLsSTrX/HVt87MDVXytviAr5TgGbj+ZSmkjicfuPSDPqyvdjFLmDm
QrDOwLItF/9q4KSW3e9elpNpOYB00wP5mVcpb72Gna9uAPU6yWbfLLUpmpRutbl3
6GriM4RkFhE5FvjC3KGgb50swx+KfWaOgpNCpMKRqWgVltA7ejfJMp8NISvpPK/p
j0C+xf517ztNC649sCTDUKRgSodaBWKpuu7KhGwL+GziTYdCLS/uSpKUqw0viQ4K
d1nyO1h2/4YX/j5QXbq8QluZ97rDoYAeIIUSO4rpxB8jlD1+raJiIKHUBt7ioPSX
v2HsUX6KMFfkMk91J/yhZcOrSMWb1rySDs3JDh3b7fIvh23jRiYoC/d8fVR+Zf8Y
Fqg0BlL0EqDh9qHzl0SSgf1xRycols5YVNpCi3avRxCbq6PPAuKCf2iLmisKPDOB
jcHHBHPcOc1YN0XYYTWpQDAPmJOc/Sk9ndPW0/nVUyRki8C0aHc3saqlBnaXhEpg
+NHFCbC53ShAeTd00HBdxmseDZAbIsvAbw1+azrq364jwTDc2JD2crFne6NoabSz
NyZX9x6qcBJ3YKDQX5ohoCZql//tk57hbJ68VnAdmGA7KJEk9sZRm6e5woDJZ0hp
RisvLBqBjk94TP2rk5AnKC9sXuNVLiH3Bc33CYnKsvHg1rnGfRmSBC1NnJ0k9rj6
XBP+upNyjzat3QOKJ60pTChAQYW15mvVgf6EJUKlnBeXTQJeZEfDqsJOv8AaWGY0
XtajUE80LqDarhjZx29v+Ro7xXdA6dE6dxqbvvAUxdcMqaEuo/5EwPQe1WtlfyDI
QedUQV0VPsT7Z2qPAOr3E/CdfIQJYkLdClze7RmQBnd6cUF4zWxNyqfr8NpRWgrr
WdOBWQvTsKzA2BHxOo4LQ7ov4Gry3uRaIHum5teLDJqylLcvvr8HAfADbX7YW2Lk
nCwJvJlPY2RYj6fn576eATrfvBGzk3Bnu0hDTa7lJXdiGigetv715685XUmlP8g6
ZIR3lHf04JGBO1gS1FY1JmjWwRiXSN1syrMgJNq1xNVauTg09XA7jfR9zHjjiAEh
osKHBxC9GHXNxSUOr6P8cy//mxRolwj+8sfpoezLPxZHRgh0hY8cngvqN02RXiaO
YFlRSwPptWY5EEefAdqerEpLbZrg7TW6MqRac/Gxp7xvVdMs/KNQXqkuBybiYiTQ
1YV6xU02AI9xx4dN2doKBKWMii5uxNrYKrYO6QKv7u9EW6+xepia32yy/foCKkac
ytGOWkT+hkNzBFcfdmOPNujZ2f7LOGWyo3sE/yBCGOUL4DQGaRLjeETxfuN/srtz
gNWIR5xLuGQPwNT8/8hT4OORnBJgO+e/lwPwOYO7r1OaySaf3tLvIjSOvQL7VPTx
BhfQJ43zhnxEFMaR9IDebLozprtanh9zjUJk4Av45zqOLc2pnzYlNftr0ORSQe8q
5x+Y7JZ9MnejWJVAr9uTlRqPnISSGVxGvusktcFvaLjK2vk9RPU99aJn36Tc9lzn
ZfzTPp7QkAH5+EaKkR8ixRiArijHO8/lhDzQqu/Lczop0gbg2imNQSkLhEHBFCkj
RY3lIdexchots00JcoMlqZ7QYkpKAWFwO+BTD7OYKkaZjPEcUfp/+lz4WG9q+JK8
0in7C3AMKMMChx9j1iuHm3T9zT38D0QL3t/ZU12QcydSCdsC4K3GqTtN4areQWRd
hGUE2noeOUEirHeYSxOyGCtz5jpwhp45CKekbgiErjcS0oSEmh19834ZMHxvF54a
yG0aeI7cTSjFsM7EiNj7ZQmZzvPwSWciGkJr0r/8ny/QhfsRP3cV+BjG7Ty/kOi8
p5z3MltbBPcwPd8wLJQmnmZJM6PxNkKAxcYEJ9qIeQvBIDuQ6IX0GBl3IXOTAY91
ZAE6dJrxmpZ8ji3sl8Uw9/F/fK0WiSrtmzQvKkXTWTWU+dwENvKs4NmdAB8uuK0T
JFSm4lUKwzgu6uqouw8KUoP2DiUOLX3+It9WFMB3Vr4KhlXr5Xrdk6hlr1LBhzNY
cZnpNHs2u2GLQtQjWdJ6fURg/Q7iBt0rQio+eZVqLt0zFnujUTaRRQAujD0wZsWI
NAV2wR+w84f9Uzy8hrJRRf2wtbSo0RJIBBRXmLLk+PdUj+EOZWxWSSCz4XJaE7Xu
tNqvQq3xVEFBDYX8LJcMdHac245iLirsqajuPfDH+JttQrxp9KhefwjtzsBEa0AV
S2O6eNBIYB94j8eAVxj9aNEx+niWKHDCJoN7RAMYcpqI+TIH8xK9cZYf3znoZbkO
FsvPnDfNfEH1HRh9uBoqvml5YU5WZKo+AvghM7f31AdhJNy8QG3CFm4uBZD4mg6q
SGJftmrwW6gNn7fyoffM6EaLriMdZtD13jgUnVJmwEqwnRtSe/4nulM9+FsRbzju
aMKXsha8fBDexIwrE1BfUj6dNCYfDPXXdDPTUtK16xTNxgJcYT2xJFnI6Conn219
zbn7p537zEwKBNu4QYmzEgPs4hBrWadEbq/2FpD1XxC9dRWhJD8y70EVqa3HTn6j
BspVdbLgEqY6cxdM16kMqU6wF+PCG+ZSzqdAHZFB6L5TZTJphNSBSKoqImSeaUyy
tc4tvTrZPmMN+haP0j4BiaNAlCW4mlH3/EOoM15JkU0tNMX0L6skPB1VXSuoJ6ok
0DQaAG3yQdZWvbX3kOgB6+UPOiIwXlpFY395fDm92mCbEJJVc6+wEmM880ifXZUq
GTSnXvhQbq0haFTzXAwXZDrhFzZZYRAcf90RJjzlmsm8J0jEdwqiC3XcNvzxbGJ9
VbBPHcEiXtqk3ohvxgb+QQgQJYEckVFZ9nrRu0lS9Oas5+2ISaXg7W2m3WuyWmKT
KE9rC6NOroynjtOnpd8CY1bPFPeHLUB8Zl+lHptszjEdDenFGPYWFmhAmcN2iVst
rd3285iNrTORoOjPmMwEdHzBVqU7HEwGgrtQSQy1r+6Nn6hSehxXbyF1/eh6187d
euh5YESV0SXeSEt4v2scJRHPjrAFiU9+DVs0Tl1fiJXsMOK6kGR96fjMT0vgeBKy
LEsk2+GpZLKOAnizsxEX2G5ZATVE+6P6l8BjMynGcjrd0PLJleNLVyx8mwMRTIQB
dyezgoqiqk2Ynz3ZFYuQqiiw0j6BSBsRrdl7Wf+LOIYDoDxs9nRPF6vNIEnBNq52
Rl2GMQaij1ABIeYUBVREV3tbfYLlx0wEnTlquJ9Vb9AIKdzpWJK79fk/Ps1M6GT8
J6fxAjGbe5rCliMuYb396Xdx9KAAtTknGz4hLse079v2ES4PFcuEqphB43t3X/mc
H/Fe4Yf5iyW7LkqLJgee2swPb5Sqf4oT/r/Vwb0kOrGDwMnA+lplftwSVRu+aVn7
n2qIPHQEbPnvUYhYSN3d5FKzdd8YTBeMUY68LGQJ3BD6Aw4ZKjbmFBKtgz23+vaD
KAMqdl/etfCMeOCFPFiPyMAuACwtjyoDXLC90wqB+IFWK+ehG4CaweXo/e7K4KQC
qy4Zpjfa1wLTSkHnenW3w3Zj/cCfZFRB+PCKOG5fyWNw70mAsqLyHhjYENbBmXt5
dbRBGax26y9BfPdqMAJjCYtlGednuRaZnQIwtr85jPUw+SLxggVnYSdtmQJkH6EG
wzGIziNI2G6w/aI+NGBtEC3Luw6T0XLNlPBKBOvWbuL/cqxehDibaT1nhf/UzmCq
iyLgmWKS5irBQpD2f8JjZVW6ockGE+hjS9veVsDihmiDyCo6WTan780OustQVxMq
Wlq7khVlwcgS5KFwVkR1b/ZWTYsO0itTIVYHjPypad5Sdw1lHKQC5fseHqVP3Rkn
+oFMPaBciCfdVLQGOQgS2MHcavBaFZExpCP1F5ZaQaIwnO/NdP7zLZQXr0VFaRhr
lN32gHOUf3GhSXg99JSqjAEjx5SvbwYF1vUzNIYndUg0Qph5q/fheYBdLythh3A/
nvCqcmRK1c6NoNmGybEXeSLkhsWl8P6Qk1dM64f9/y06YLz9zzN3SXnuBK1O4q6Q
Y5QV+PsV/RA+ChpWXjd4BV7LvVVvJ5Zx4kNgvzoT1rZUUpXtMcCuSYoaI8XYRdC0
ZN6DjUAhBPwlLGvS01M0AtFQPlopkzZu904YjDEuE/cpPLsIStjillvuXuIrzRws
YweMxAj7Mvprii3gUyTDRnE51pBCvtXcqu4JA0vMmT+VHlv+kts8ShU243kkfV51
R9TVj8WR8av4+ZNMAipLDG9scGnkqGolTcoB2wqAJH4b19RA3ewsLsKvE4R6NZT7
imtYFsDjej+FyndQcM0+paK+Og5bZ71EODRmFx6hduajdPw2Kd2FinQwlHfeMSfj
KLW9ii5DQkgVObGuXMdGwbUCIFp7oBwflTmM6THmw8D+ENyXxAh3SUx/nbPWHuyH
QBzUe1PsMtUBkJcNR2iOmLfuLbOzDewY34T+Fs6Ayvzy4PY3buJYlGo0F//F4K3T
h71uWrONh7y8heiG3xA/MDjuhiXrAJ8F984sRv307N/onniCjSYzcFExr2W7NqYF
a1A2q/C+b7QwvYCR2o9cdS3ma4gjq/dY5sWOom2gj7Zdf0pC3StHG/6QAd0X7dDs
nCtcH3so3+Gssi9hGvcnPDA0Z9ZFdvvj8EegoI2MIc2D+QJArTnsD0nnGmd/Pvpe
5rqXgCD7g0jQLRMlCOvKOQ0l1MmZfubnxsADyRC/TpLSqAgXJOrsm80mQWvB7n7Z
u54fgByBsC2hq8992SBchsOBQEA9jjodc+hSsosayliUpJ8CQWkVdhrC9TAcL+WL
j+dAyMGsqQpMYIZb6gX1yG0Lgi1f89ItuzwbO/6FHV0TJsnmovSVHas2GcDC3p38
kI+MKqnr3O+yNq1EN5843mqLe1EnsWRz8tv6P3I22T8hPEUr6rmp8mApu+9DXoVA
0ebc1balzKS74uRjwaxNw4WfuVX2v0ECJ8OPQNQqtRFccYDL649U3TANWekwVJH2
4odAQ9i+BJhx8pHiLFGtZsfSQ7o8ztqXHb5IAL2sPxo3e1NXkHYDNklckUTDdstT
UKGVqdON7KRccdbIDGVWIumdoqVmqFmhqamoTgVTj+10uFRkEf4uJ8l5PSxxcyAP
px6EkBKZV/a/NKc8L/jTWYRQBbeIEsrjV25ThwyzJUaF6dX6tCF7xGuXp+9ez9g2
wM0wUEK7i82tZH4U5hcuS0m5i6pAXKCmvDBpeuCXxrmYoVPhqCAI7JHPuvb5W7Bl
xF6PWHaOe4Iw9cRYS1T5ntMZ4rjLOwU+pF0EdBpXklWgEKLmNdM0c6Y9jNae4KD4
7t8YEeQ8ENRi1q26+y/6kEsk+e7dcb81jw7kH8AyW8Isql6pQulMTpR8YcHveMfo
EiEbFg/zr3tB2msaoN1Aou8OIQAbU2QCFlGqk68i/H2KIYJQwkEJG/Wnb5T/veTq
ctDyuyPbdaAMu0wlZUhO93Cr79CsFsP7QlvNOcdrYU2hSGZdOCtah5fJMzkxTAJk
cZ2EGzXEYby5qpX+S+snlJk5ctKbc+A1wmObzCPt4pXmJpD8rf6JJPmrzMYgmCjh
2QEijpfg1UUzBh6hka+H0CljWWRYJo+RZDbBYn5TQsJU8Qs1CsXOPyj94ESiqgmr
3UCIbRqi/mSwgxWhermFA7HsskL2pRYEOnSi0mOTxVDGbKoXC/Q5ttjwZ9rqezuY
JtV85yuhhbi/t26EwRjuaH7TeeAv6eH79twUR4yU/nfoQF7ioW9BZfeYLJU6JMVR
ofL8pOAC6L40xfKXEQoNgwhTUkE7MIQgEaGs+4F+j2G7Y65rWDCezo3jC6L/5h8u
Hc6hIZXJMXcZRZtbPhju8Vs53rN5V/8plHSo6VjqTmyrPg4Tbdfn55RBEpqLjUcn
L9TTKODtxEKLBjBrI+6Kc0CCIJiwX0V75Vt136GQLuzevc1GETHFW83kuNbkOf+u
SBubH0XEaUpm5LH5eFnI8CQ4CkBWFgglhwSQLYwDWNkozZxQ1okK+Jed8mYKVzT6
B68XnXpyfg0rgyWPAo+NjHYj+rl9Zept+58tsTYUuj/bXTNP2mDzdtMgsDXAlyL3
kQIB6g4lX018on0zCmWNBEnj+4jZbHqrtfR7IYYisTiwUPDpIaW1LTYiWjkKv6an
u+paVz5Binm5zUGwbO0cWMB7ul2z33ll3ILZfRe9HDk2G2fkVV6e0qKYtN0FfHKR
7JXNb37KAUEyMpokKgetW/dTpv3Zg2O97bZi3Ak66KB26k8IxeWkO0H+ccQz4p+d
AFbiD/oIFLRurqvbND/mMyt1LNFaNh2TG9yhiP1ebJb/dUkQYMOAe2i388PGSeow
asIT9SK7fmIBQ7SA4/Th6L8RTBlrKkMz/fxYIK6aG9+mHUXqxFP8VskopfdAL7He
xxjKlhrvePN4ySWsaaDJK4B6mDHJFpX9/R8Q1+G5Tofpgk3NxY0tAhY0OMnkO9Tt
Eh91hOv8xKIGX8y+fUI09+Vbsw88bC5Wq2+UJN5AjYpqkbIwq0UplyLMc+Zhjvys
mBNPpNwtem0r2McgwmqHqOV7I46YOV1g/cKWzR5fSDlpoo234X5GD9vrd/uj9PQa
qpze6QlmCJHu+02dYTFQHYArpocNtmRl/XlRDN9W9Z8nQYWgYp5idIxfO3Unj+cK
llU3gabzbh4sdL2iYEce1RgVr4ai+cxg2wnhN4wQlnuIIDPD24TNQmVt5ii+IZ1i
1YcGpMLvQ7ii8HYXUIx9kJ2Y1cUAOApenqsTLW455sJ/CrfJGjdU1EHQFcVDqpPl
JnMkH3mmhdk+qNLOifR6+yb1JN78qvzWVUCraaran4QEPvIR1zmv37VrY+5cra0f
OARkUhUKpK9gkiUIOphjsBvrKE9sJ1katFANwUMUKuqKSwSu7DgTD/IjRmZNQGul
adRpmoksteWNe2Me6JwnXomZJCIbF2URnfgcUO9YSKBIKLFZ3lksg31C/iohYFH5
5vh/v5CMQ0Z6/5CZ9KzPtDx/X3z2YrKYjnaMzEt6+1oNaY/fy+9PVpkiHgRkv1ff
7sYbBz/vmZGGEn3120sQcTuh2Qj9rZ//LgrlEYbx4waDs4lHgFHJqU0d8PxeGzD+
7Vj98uybnhPy2jIJcgvMVDvdXSiwXW3OyshfUufM9GdFYw2uTsnRsTiBhJYj4EO1
gOMN0Tz6+rhf4PxkpTjCmfDF3BVf7QdJMgPyLlFhRp2kfbE3S5UZhsziktl2oahq
6AGunGgZwssXLaaTtcX8ArtFXjcnzHOM8Nyxy9/vWOD9oEoAR/0k8GDAJI6I477B
8GMBWVkpe9hx7Y29n+WQ04DCHHGahBagauT/IY0Mf6D3py5UA+hdjZMgigbbsVWz
XwyUGdQN3avRX3YADriBjCTr7g6hEDN+0DJOKOH+OWSxHB6l8GJ5/HDSpemP1DN4
A1gXWfeWQxV4j+CW8qSVpkluUeF8Q9Ypk5YPktWr3OzBh8MvL4UKyhvNmD+ORpbB
QODdjucxCm+0R0PSuQaCJ1oWoIuUV5SylGqeIz5AbT02F3Lm3ETDphG1lvJHX/3s
a/ki/TCDtwzY5WpugB7LDEnJ+Oxe2HCbLwPiPhj6jAkYXa+TYSQqMSsuSPjnbW6S
OYkr4VC94T3Ixlks+4GPRZDTitN5xW+r7pGQgb49qrgw3d3O2xYW7sUQuvz5htp2
A53EexkssoS6dvxzn6EvT8wQkLlW9qEHI2ANn2pJrjckroZC7+QVxt/gnJ2aOXhG
KG6DqxJJiHRELkAAmbsDK8PEpqexPdEoyOyjmsgcMtxVBL5wJSl0OVt/baGsYuOq
SXgXFDIjrwj9zcTzqiAKVi9L00XusDLujSrhWmqeAe7UUz3XpbTf4bvbOMCK3R62
ZVeE4KYeMvLTDP2UsYQDBUscEuU364j6H+esaoL6FwbqI2uG6uUCpxItxYpJKEMG
1mxNA4Hid6/IAJtp2V4PHSAND4cxpQY4k+kVSLZQDRdRqLStUhsI5VVWnmO/al5Y
EF0YpGbKDF/W5QytHKpy6OXUTbi6VM63o+7tb5nJEnbFxLQxCbhYfMK7cjGg2ZI2
Nfa4oWBVB5NkLdDJqU2/DJQYn7YRxW4qOhow3/Ac0XxM/u2RHVn6z7MKN0bvSpM0
5ONN/P3OFVUY6oH6D3Aom3aaWI8mP6uh7lDzCKLQDS5aPuHYXit9Y+Ek4PRgudb+
2TZZ+PYX6aHFkKLlXYkqlUCTRCtl9+Ca+tBSiz/ybZNhK+r2yKGiM1ZSSE6GQ+B+
q9b6dvBuuuCmmNK+bAMHAzlm9xiO5p61ReEBMzItM0xs2ThmlV+5abh0C2nZxWUi
OGgD+k/oQFaKBHDFFrxonaE+6Uivo1KFtJHi4zcu/cpEPuUIz6nQFi9r5Ji5r8a2
dK8tRzGiOE0N1mRpZ1QSb/FFVBpe7vXKawx65UAPfetvMqCznsr8onSn3t4DjOZG
e+P2rBZaSVx4AdraNtPBjbBe5ogmTjXWVEnlNCDRftc0z+JzUOm+l9C2o44zo4tb
PqGKaKRMp0vH/wrTgkyjCiQ9/IS8yaM/k4jYHIKzSGgJ6hZQ6RglfhHjuVHqvx0S
SIi2URkiqJszRhNGDxVDuH+wekAJPFqFejENS6N6OACqIMUaRqhZKb/TzXQqWaAg
049Pcp1NTGgaHutEO3VJ0bFjanN8Of5e8XOj5zra9Bhu8y9NHxng5ShgEH/NIxrA
/TzzwyLVFum0a6eb0npsxIblMqBqdmPj4Cj9sa3dadYM+pp6dBf0B/4VW+tZxLcm
Db+GENHBeR35iCC54fRTjXjHS/bDUm3CAW8d35CwiggZXmFqw/QvXzSXfiIi86iy
67PJWoZ7za/+y/Rkf6XQiE4rVJ6pIJoyCg4AqFtTDqjTQV2lxqG35rhjkbCZnr/P
tyK1syiw6t4Amtc34H8hc3PalqbVvMXQaXezMDSOC63sleUuImDE/vIYu5VBgL1z
yHW2LNPABz2Bobm0V2rhyt88wNFeaLaLn9gBBXPvPu80P6rePNbzlspaW79Td/H6
s0NmJ+I+YmVtQtPn26QEiOZStembfP+xLkN1T69E9u7p1xbCKbJsgf3vQV9HVsNl
x9rRwKhwak7Q/gcdn3R8DqoXuGNrHOlkZNdiWUfAMvZKid3+wUvANAbT6eQMOFly
af21BevI0Z7HdNwl8uQbv4vQBOuilpwjYBz/dnzV7s9tho40w7hGjUe8aNvjc6dT
Kw/Tqiad1BYR4vCRpWJhsnVwd+l3NAXZLVRN1AIw4xa4/nD1cCDmNOmSrlrwiLyV
YmX5fdUI2tMUXDrTa7EkoQl7Z2nHUxKepUdNV/NEgyHw+GLAn2cHaGpN6s/4tSi9
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eljkTAf8J1zksC8HstDz4f67ak/Ihftp0OoC8eApyvbFv68q40fijkv4hf8C000G
9ckeCNhq9JGsEFV3DjlGkOhZ0hop1GNBiEa/gggjfQY06n0eeH9pasIzzQ6+i5F/
xbejORemi4I2olW9yS/98Bp40KgyQeXnvL9yG/xGnITZuT2SSzKz+nQtFegW6KAE
wnJOQAKx3pPeii0mEvn0qZVNzWVuSVK3Q5+lua0BllStk+LTxL1VtR8q2XyJ1z04
WIek4Vzf1K9TtcXJgeyDXelVFbsvZnjxwNjwepcsfbdxgzOrZUFXD9eO4ARAyj+a
kZt4N04rRxW3oB6e2wM5+y+h5r1443yP7+Ahb5w7NADWY/HaXhLuE4yZ36XGukeZ
nNNVwa5mKyKjSxsEYWQbZCGmQdKmJS/askx/yaQDsBI9gX9IvUaiEHxYgOefRuIG
XL11iAcVs47Lo0cTnFPUZzJXMXk0J6LDSgFYEsN/AJ9VIDm2H4NuWt4phNecf6ie
nEOYoNpUkWUAGSYcUaV6S6KofwScI6BEdWfHXeeZxjxlJZPtX2/n8IGnIENjttmr
BE7WAo8YnhwgcTOgbUwjVAownEmv84N8ggxmXtAreBE/jUEtL48SHdMeXiqqR6Dw
h1oWywORe3nGSi1SsglDY1RPLlGw6+2Cp27LTNPIa5uyFFH7FRDiF+q0SJf5Rm0c
J3p1JF6gLqy+B5RzdoLrk0Ta7O8G+XE+Zktuyx01S0TuFug47KLKB0ys3IAx8RIq
xdAcEVfdcyoBb3UIASOO3QMmJrwWDbu+gWI0agSIGa2n1j5IcQ7x77eKqhuhAt0Z
eTp2GYzhQdAcZ7MFRkqqlwnPeBhOG6ewD52u6xTBp7mA2JNTwrc7KdqrGPxonkg9
86yW7bQ12to0bXFKp8s5cZuMm2oi1jWzMfJ4h/kFNCYIOWd4spn6RraGZFPBWk/6
VADMzMmCZyU1Mtt5VbFo9fw6PCOxfbk7ljAHYEsgGm0Bji+gI1JIiCRZ5b5bnc7e
5VYc+t30X29CfdaPdafmz21lMTCkAI7z5STb9F6whlSBzx4yKCnXz9tvMFzzMeSy
KTouZrwBwOVw6GoGDSDcGik5EUEmd2mgSEg7VIV8xWM/C+aM9LjjbpXYo6Ki6JKj
yR3MjSboNbP/LT9tTgp0zQQhCKlYSFJ/Emi9ecpf37rG2ZlnzxgsdKQoZ4fpXNxb
4unTiBkgAPgODl5gk+x+pXaQinkncBvkamDzJ/qFLypPFpj07ai+dCIYYYqzrsWA
WPzlhrlO6n1VoXBOl2CZJSmltWXFN1hsf4LNiWWuWzV8BsZZ+b0Ym8jqwLxOdHFl
jQYL6uEMekdGhRxXhAWSI7XROAjb/LzSMxElwO47kSguPj2cPrK0SkLXvJoXK5Ga
myfHVK8pcXs4ZOX+xqkk1fX3IDhCuCSudpD0kk4iZyxNBxlfF6+hejdGVZYINiWE
hhEN30VyarK8GcjeAPlsJbODvI7tX+AUDsoNrBknKbs=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
On7gw+3JxASakZJPB6zxBiAF2Wu65iuBB77Mtz+sglMc/bYew4EiOVLedf+cEhdV
tzKqyTRz5xslG6n/h2NxS+pDwqATm5bA5HY5AEkyBG5X0R+oY1cw41YFSv5JY6ZO
jRTBgxrvONPsgSYvP9yhpwN/mgCxU8hN/YtKwwzFLo5ol/KuzPz75io4YpETl1v4
YIqgds7SvWXSfEoZD0bLcdz/URB8vC7+oA+Ukr/XMotoL/6JXfUrruulIURI8o4x
NwpN2EhMxf93UHps2jQOF3aj7JT+01GvUQ5UgaS+OpSjuKyno7JniBysDMSfGCN4
NkRQurkBrKjT1BJfYA5bzuUNNZDjMDceCOem7nyzOpfl7PDHwwfntsxIyMuIym/8
RxC5vty5YeGQ2iLDVq5mObHA/3srHSpaQRYmwpxsSkQIuo5eP4gRl3/8ElBpmX0l
Buat+GJBPfvkzQIOoctTkKa8UaRfkEb97NJBRCcaZ2F8W3xglS4GHMFounBX4tvT
bTkEV1+dX9JZEwQZmWtOXkpxj/UUZQIt0UBvp+aJ3LmJP2Q8nFAaht+fIpdQEP74
A+h1um6rgTtNVXAAzx50TvytRnM6b2Dpfva+lIvealmxdWis0yADdPhbWqapJYPf
xERHK3PlLE1VIRoGAOxwKSknsKZoXcAooOncP239m/+YdDNDLe1JjFSrVc5FTyP4
dd/7c7nyRuSehtJ/do8J9n4XfI2Pcp1FfeJXE4ptuNtRL6ukaWLNSQfcGSFImMSt
eF6A4r1BuDu2hJ5i6B+okgUFDF2dY5T0irGwPIsySyrmiDPEOoJUnQpjPX0uhRVI
CI75qkBm5LSZWWpoVfmIAoc/euJ9Oi0idpA9DDnlhqFmoM9b/BZc9lFQ9N7CMC58
8l6P6V3FP9wCdQRCGt9dK48vBefPcPUyQ900TXOkHao=
`protect END_PROTECTED

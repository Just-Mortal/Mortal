`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xIzhSOaPmOktHMt8JTaBdXiWkvhRDE7Q7caOIMbK88G/JBBN/PjaC+KJ31VcoBY
y1XFzJRFKbbBZI+nMyEURX7DenV03OoEEV1uwYZm9vv2cvY9Bc9FXtbhSYWoBKv7
DS4StNzweSHwxL3VVmxc7JSQN8L2niXNYVcM0H6EQsQVmFUu3Qjq0rBor6J8EwS3
eJZL/vh/1bIomT2JQG3btUSzfPBlhEi0+J5vYiK1zNvjkRD2OKkJgBebZkymWPwW
h5XTO8Nudz09cSkS0l58FBpyCA7o/m2e9RUt7yzG/N2eELPmIIPCDO48fINQpGgM
/NxbiAqSXRHAGXvc+Uufi2IW6XzbkR/8kmDmDHYEQrwl00TK/XfH2/EXt2g1ynT8
8/bBVkAQ+OIIbUnqiiRpQ0lwMYmEB5plGQVjDlmYEG64tfLD0D6UyZv0DNt5I6/9
lGIcDIGjQRzhoPYiWTQBPaifGlTvBVnyTEI3Jmbi49wlKoQn0dK/BFMw1wHjXW/0
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yb7vlmeCkY3u48FWS0XkhlGDPEiAZ3c9qxB1cWbUJin69kxYqCS6amKoPaRKVBcM
/5b1NK1EyceHI3NsYSMWNrK0Xt+Cdoq+GXS4niZT6GfriPkjsqY5gpodbmgei5wW
pRAAscv6c/1mJtB9Tzs/+xOeBW0TZcvHNHr/VmGbaWSwH1Du6A9pCov8Mz1LYLw0
hNrqM10IzNGeI70ydIF8BSN/KJVzxdMxjCsT2/PxAE6wMR1kMJatxy4sMLp+SBzN
RImf7Uvw6tPzIpaDOoRhIliuFsR8jaBXIxekgyBfxV3dV3O78aEIdhc3XAJjmWCv
iXUHo62rtKZKxuvm1CO6WDRemtk865Ef1Dc8z0LJwgsZbtmM1/IwLFGBzZIL0pMP
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXotvsR8xuySqyVTXkiK6t4CGD0T3mkK7tIGXsF0tREYNeWrObaM5TIaaHgxQeZ5
Ujj8P/o7pGhuW5QkOLK28WJLmSdirJksdu0NiCbdW+C/pNCeEekLpGI1fYxjvWaP
U6Ukbm3AX4DXFcznBOqd1zzn8qhuf2Lms2OQCC13lkLUd430FCNP/Vh55xTvrXP4
7RA/1YbB4Px2x9bbs7quKmj8zJhEsY9eibMbwMRpXJIOX/TbMmtwQoplduUJjbSL
aEP0W57M/ma65+aUCPPOIPTQbN6xHQLYhxTB7yO3OLIYdLtP16d+BIo5cP3mt7F/
QkYQy0Os9ftLc7Af5k3o/+C64WhdFSto6e+6DPdxcqFl4MhgJpKjJJegx7PFiYAn
vkTFZWPkCflUBPUJVXR+72B9P7qYDkrjMJBQK+6QpAXFbgHeXhkHkie+ZF6Nqf49
p/7rkMx3SHG2icbDBA9zGJv9A9rjbpuYbfSv5dtjiizvoDPF4ZSv1zcljCTEOx/9
Tq76uRtLznSn7RnyygvhJg==
`protect END_PROTECTED

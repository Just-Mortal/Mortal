`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnhAe+suuDpsqsfxyf4jSW/z7sl81r3gzZVRopIbPI+/YKvksqD8EnPKYzlab/gO
VCZl6wh9dJlD/85Ok5hohof4ReVtY1WAT/YbtqvuOIXkE4GovsoQur9cdEsJQFd8
WP5V6SMqoLlUIJCqqt9J9IpQM/6AOLwL5+frDLask1o5SRtiOIyyvYBcGaziNpEi
vJyxXhh2gmplsCIKFBEnsj7sXTxXnhqi9EBgECscAaC+jNvgi9nqSSvmK6lxtnOJ
t2Okg3p8C0HnwsRhJfIXLxHC4sGHCYtpt6TEl3S3cN+gUScsGNQs7+oTOTVKK98C
RIQACEsXUmRge6mIinGw37CgUODbF7nV1QCAQkztU9TtyT9t5eKxx3YEAjpKN1rx
8hSnIYGGg70SYzFbE82CiYzrIGEyuEi167PsH7nnMlOmQCBW6c5j3wLNw45Ydbmy
E2HnF24YjVTW/7rJAcmpg7OTaApsxYr7QJkg7SaEuGPBEu1i5mayZX8VRedr3f24
flR0QfZuFHSBG5/Hi39DGUjskJVL2pIIGiPPwm8A9Zd6/M8KrCMOy/8OFFMQ/Ml1
hTWjneduEG76i5n2BC7+aw==
`protect END_PROTECTED

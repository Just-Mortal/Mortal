`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Ts+g3PZkFV3U21s4FNIV3nODDBwArjVXy6xAoSYi1X6AqYefJID7Wson3nixW9d
eYdTlcFEnxjUI2jjgrwzptgMD+N9eKWQm5vSvJ1fejQA46Yk3yiXVktNuQ7daSYD
GK94FDYyeLl3DqdmYpo0kYR7vXb+rNRsV+Ua0KJYg+z/a4h6HkFONp3V24FG1rWK
0lbmjrVxIaY4SPZiRlKkRLfV94iaxMzjTme2pIn3h3x6lV5S8t4xx288TyrQeBMY
Ql+WgeULtnvBtnQKowK8gXfUgBkFgVYyh5rE3tXxTxe48Grk2KoMpCnw83iVCKeq
PvGTtrQEf9bXp/rZJZYrGJeJs02eDYOMH8x94vMCdWQS520hViVrs7v5yDeK0CV6
gNqT2s+y8GbnPNab27p5hzhsjdaWiwcl5meJgyFl52zvET+EOmXIAZZ3OimvBII7
uDRNMh154HkFVkiuLoaXiCYGTap62tHxzmvF8VU0lhM=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C+CuKi4aXvZ1H9GZQrgzlHDKrOJ2gdtmIUeE2EAo8wfAWF2l/I9KhpEvtATUo67g
YgMmSm4IDjYkn3b9mPheG7VBOZ2w6wlyFsPe4INRk1sllpLEYI7LNncL34wiuRUW
hADqT6tdtn2Mupr7du18E4Ih7HkublFpDAaFvnOyqD1+XQF28bBS9iu0QS4US8jW
fykHP3HQ5Adp2QPjL0lDtRtjLZKDYIse3TeU+M5VzZti+PCTFI3gzBJi9XC8US9G
XgPe5qyNhcHX7ee38o6KcI3LxCtHCrCQG47lprlpxfySz2Yf3FmnGgpPD8OdJVBz
Wqr0nk8F2zO49j7QleLqfyxyb3f5a0Sx+0hBJ/43R2qLOex9iwGnBR+pmnROqxtI
P7m6SlXsuq0CWC3GXa3x7ZRERwHG22HlyIqEkkmWMAzgUwKXt/iAoTXD7T8eGbPT
pGGB6a4HIDQDc9lP5R2Xc+FnvHN8Favvy9XWpi6/zfPSy5pYVyP+SCiN6CxZgDLE
Y/gnIEX3L5fyFglgD17qHMo5Z676iGhFEtDhF1AuyZ44KN3qSNSe7+dEY65QLmMv
InNPxaZ+afUsd0yu9iIcZa7wfbW8dQyijaTD+Klw3lmRia6xwaLHqsI3mjPqs9pz
aU/sQ3eIEjqOQlzQ1HLB5I+48nVo5NGAZXcj73ir35v79XbMgIq0OlAnl6Mo/Rnq
mGRl4vskPW6pAZGZRlIdR/7ugl/S29uQvOMQl99oPJjJwtUw+6u+gPBTPQAKZY4N
8C6WoESx1pkM7sHiPmb9edVBTtkRH458LCx6qCRVe3wfXqjY3G4HP9k+5DOzDmqq
M09s1cs3815/7W0vAIP9byNON3jZNwLb6f8xOPV4XNVz35yy0SZwO3xkKfozDTzf
b1HTyb0jTLfZn9UJPEi8tNwzzNkxHgzFHbTaQEaZgq2c4veHrNO4HntswcVk/Le1
/+RbX606bko9gcYS6Spc05GF4oTyuWz/EthUDZOYyRsQKKAiqe/On7IOJH5mONPe
aKBTDet2IXRWw4CjMliKH6XmogM1LDkymhj8CqxURbHaerjMF26J6L93JQCIr69X
pWWauCZmz2flli2lsuFLiaTT0lEgnw5X5atcXNN12LiTG677WiQc4j2pqUWSwqxd
y3Rpr89qeysgOi0feoJrRhm4w13Lcr92EaZabrPLN39+dxWm4Jf17EBFTvLngPCm
LP7qSwajQmj27lazwGNpaIYN+O6mjHMNlbZYZOoG+N2Roefug13JGKMrSNVpGJJO
aZCJD9dQgTaS+jNR7qGJIeEe5boKlSjLQy2TKGpABe6PuWUEY5a6+9kWlrnWqY+I
+7q3MpqhzAIL7366zXlnVuHFwPwrHrgXK5PccNlpnYqrs0D06D9zaiWWCF1Rsmm3
hqJTyQvHmTNuU9zI/fanR7xzsZ5T+VziglY5nWsURYpTReWzBtWTIph8uvQq5ruL
VjkFtre3KGEQHY7u1aYVuB+xCI4BbTVA7jxb02MUCI8ervpdZY4VVzJVV7uRC7Cz
8/qqC+JZP1EKsibJgVUMvozzLI75mKMhZ9zHUwLfe/15H6k9I6C3t+GAgs92yuLZ
q40hNuNO76sjS6LpXKFhmtXiKLDYINsAPxkTLI5/HMOd3+Lti4A7Zm8JthmciAFC
B+kSQeKufRZ2hOeQ/iMhSdugFKE6s7NI0HAsNSWNLzVRqtJhC8MR2sBN7uwxaFh3
kOpvixkbpc7z6nmAhsS77VXl5VagI/mzds/oeGxE2ZGtoubtxBOmG7B/EgcAlm5/
8TzT3cg55lUlQP3x/2oQhG6wXzzRSmrtsMi9O0wjZzQmmyij3V9cS6FjUvJ8NXOa
UmyEBcAdk8Rm2AhvD2gDf6yCBw7m5GgGRyOjGkAs1gKoy51MFcoTwl0PLUd4vp0a
8Dbn1IvsGpeJcOEkxP6x53HfQ02S5+xaZ1kyzkFxZxFK07rbM4C6HICbCZ4MOqz+
5X5Q5tOX+mOMmJYCIOH27+lfk0cHWMCTGZKBfuwXQG2JZNZn8teym0bW0Xc680Lo
74gFG/h2XZ979WMQxMC7iwJBytCPNDRN7q06YTVYqPC6uTQrIXpAJuckC9NjWaHj
/CB7geEoZjU8dcpM1o+Uit6dv3c3cGEjjXSnGe8CGNx8z8REdM+PH6S2N8mDLFGN
i3CjfZAEQtav9Z9jwCsp8o47dG9vffC0loGoSkgnptj6pWYTsECDemgH7xbLohBn
ki381RdfVuVI1dB9f3n3ANMChsNCJBUyv2GHtp7bQcH8fyJ4hlNsxQtxg4pPngMN
Kgh6N76JNDvYI7TyTZpGOInNZWcV70xqOHADtFh4GB6viRKw2cKdcMHSWt0GFT66
aLwcpc53Nb4ROMgDnYjVoMEyaGTHiTBmhbUQu6fJ6ynler0b5CdIqY+bICDcwMfp
xmxtxCZcHBNfANEhh2GMfbfHZbLx7d9sjmRV0CPAE++0pu579WZUQgqCv/4gYgQR
VXBcMary01t3HRJMjHTLf5UwjTtxWfCrMcaD4HIt5L77PArqFxWx9WUvswIhhzR+
szOdRv2RJno34N46OPul/1aKuarRQHneQAx6+97c8PLO/6tYakpj8bieuJrC0FlZ
Qf6MRIT8T1GDyvTEF36QbbzGlbLY1p70VdW9vze80JenE9ZH56tldDlCsJPeZrCQ
oZquQ/KGiyNCd0afPJQES3SYzYfVNvGhf+3zYj0iXdoD6Vut6TIBTqafazD6qQOg
0MilH5NFY3dmW+lkCZXYRMmY97WUyJ4xk/7fdCPRFD0zj2qHtCUBylemhTvL+yEW
4sl2iN1YXWRCzIuDwjVEdYZgpazoqdALi/qgO2bslu1J7hxWA/vAjJMwWR+pLaKg
ZCcBLSklEwCQtX2yrNuaZkTNbo5/zKQ/7Sj3wGuKbExsj/1bVDZJyVwlD+c2zIhW
QXPj968J98hglie8h7UmEbtYLKt4zNIsF30b410/qjjIYVnPpuh6sC3/xQOlC+in
BAQ3otvUIE+yrW/3H/7g0NzyUSGBgkARi5WyUAmtD8jOZdZZIx4FoF9+3RedDzJQ
gLnLzcHPNeNz5dV1SB43Xx/pJbbbCSf5BKzxqQTOp0LZMDKvsso9sXUq9th0OYv8
iwhTMKpbHUi31eKGqkDNoLf+8HXOwISIacyxWGTufljjCke/r3q3pRfqMxEXEfpN
ZoQNXPBhFpE8PC+VfFw0GtjdQtyYHimdXjxbvWmolHpzckJMK4V0ahShYzxsYddf
ANJPu+CBc/eJuz3urGXrHP8ZJMR0z1aIkYCswLZAcA9XEfOQCaRqj1bEqjXKjW4+
rH5V+TFHGZG5WwWcEUdvIazd3VINzY4liWH+qfTWveGBJ5eHEc+7wLoeiac+Tpu2
JT4xlE1DChYOTY3TsJPzosXSc4JQdtR742muiE0OqsMeAbUO5w8oHnQYPQfLCVj6
tqK0TI/wmS8ajz9/Kwn48xVeVQIOVNBLG1euPAEzfCfwIMX4V2Y1s8Q7CdJmydyx
VlCZBOk6ZjiKhgmyXbubM4wtMr627L/qYr5NKJ8OZrMBn5rvcdTMcU2dn9roVpDe
U8b+cZlD1E4nKJZRjd3L36fcXpFkUPMHBefgr1WMeAfQJ3e6dcI4nFAPdXDgKBEM
ipzZAqqmCQfaBoLYPL+9YeuZQoxAhXzjSgKjPvLvJxlr1txUiBV4Zr6tS2wBj2gK
CWGyKyP2uurNVopjgfwWsl7mQDN2fs86u4YyzraTuIifdTOpN1ENkzU9tscipXNT
VXkzXobFAGvIF3W7sz4j588cTZTA9DxVwzVUPoUjIYh//2ElhMXvs/SOZ1z4he6v
gTSa6tVPH4JnIukH1waP1kB7/U/DPgbeJmORby40MbFhJt4hhqxlvHn6Yhe+x1gI
sMyzM0d3nMBlEt65btGBMtUwegX5z6Vgk0mno/X/iQVsKlNzaLnfU7bAOXYbGAWo
ZORMIsBu7XzTEiRgPxeFh83BcP7mbxegU34KepbIaQunFO1+xe/zLOMrTNqaTwA5
2/Xu/wz4OucMVe1L7GOaA0vOymM0kjCEJIGuGjovoMEm1AjRooJBR5XJzcGbP/Qu
fe8bQv3azpMsqyOL58c1bFLTkNWHQNmcJqixLu2KoJ+JWosNpq0cka4YNcEopqEI
xkHrqYFiW+gFiv24upHJYG1DnBmn5/wDx4JLpjSY2B4I7KjwUogVHy5POXd2wU8X
5hdD+pS32ehjcQTHuANv8xOxdSHarWnQEeYFwnb7Ye3F9lLIXt8Vm3+mAASqzg7V
85HPsKB6zfxNUTVVZCBb6Vqswz59D2sur4WDRMwvWQhuOoZOOXIrGPr5YXvZq7uT
WRObduZJ9J60H3Ta6M7KjBO2GksuwiZVQXAQ0KtiXVtgTpGH+g9t/BZ2BVVJADdQ
BbbTeA1lLvWzeOF/lO7FNeYcbqQ0X8g7iVs1KL7fts+sKj+yQzCG/e33UTNosZsy
QhE8F3AQhNvNjv672ukGGBOIqPx8QEueZUy9abSk9ZJjBhZ95HITeFmeKBeRmo5k
gd1FGNh6AFfpqO9wjev2E7IqLlSHcFRPQ/r9+oZjPNlZW+O/fN1/Vjx4EYE2BPPX
i4MmLAjED6qpAnMVbyPTAtQ6dG38D5sdlChbB6EI/PwL61LirFbYBjuj4qrs3zN+
dVOpnRbyVe+Nj/mFmDTsJn+f7tTspiDqCbRkPStwQQB8LezdCkhAnA8j8+nS6/Xr
u0SwBy4/+9HuPdGNF/5fVZH1PqyYt5PMVz3Wni+1bIdGJYLkGO+9jHc0l1fqRQPs
oMQ47OkLdQVSUV5pOspW0El2A/MB8E+2ljw3ro/gbNU0AaxonzX81HQOieRmeB0+
F6EYijzZkNzrcC1xeACwULwZXZcTDPwXSaAx6dHsnq0neKEI38qUpPPOm5Bdu7am
3ZgJqm847TGBNoquNgzmpKnquxEt/iGSY0j/F8IaVpp/Dya+JuikaM20ZJuUlR81
NPAbR7wfUNjpPDLDJb3Z+1SRC6bkDZ6Xdb3cj+4Mssut7ilnkzDabWZHwVCZ7gcu
DvNYVn37utKSYbIDOOnI0Q==
`protect END_PROTECTED

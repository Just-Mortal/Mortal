`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uklg88v9gQL/YPMm34qFUkPU/GEfO2KbErBYEimJMatIMuyJnN5sBA+j4j+9DQVx
Pb83T/3oE0EewBkWie9Qh1iC4KhCy98AReHhU+vqNK+qSkGsEb2agkh5vO/H0gIO
J6haxlF8j7sxE1l2IX8WxY+otldVs3bwNaRXJB8PSlcXo7KLWokhuuu10PJvTpl1
S5HITadPxeIQVRefdB8ugTfoTDBvuTXI0O5Q5ur4HDdTuRYYoEtIlR1/hgo+raVm
WzOp9WPlg8Bm1de33Gg1jqvHUjy3V0PQNc8oW1L+OVqurlO5X+qIIdICa3s9C9xp
PkZvjVee1gEct5SwVGChb3bEV6UvmhgVrnH8RKTATs5zGVBFAbT8uKPvYGSpr3i0
YyaSErQe4F3l0hu3SK2lYJD+9UFIH1lLwVGg+3A8kofgyGPw332i16znyhw5kgB1
IBToomX18eKxuAQu9aOZU7/1KL6FD+N7ZTVRIoe1qb0tOaAVt6uoI8DxDBTY+So2
1WSwRa4Tv5IDMQOPloACTc3VITClnlAwzBD2Qyr26Z9OfYH4skAlpKil1SJk8v6b
C0Xzb7oQ1rOCNH0kaZgeuDnUa/uSJonCIL/uld8vmg3ZioXWV7G3ZyJXd+h30+5v
aZbwRm+5UYXU9d8kR/epxmLBdZXaalTbEFIEO0/+1MHt5Tumx7v1ej2goFyBUKHG
Jyk6w+Lj5jQEI4xjQWWE6FQKaijvvF1seItCzbbaa1hh1mRIRDqvkB1Q7jPyqiWI
WGNi+rU6M7V8KjyZQKOgktGSzol3LRkGRmiIK1zHRgaKpTtYpmhrmKqmzXO9fUGF
HOMyscorJXHZJe9RegiD6BaJKtL732Sg0Udx3IZL2lcZmzG6fhA+ysl7JtpZ2xM5
fL7NfeB9eNo4szA/okIN6HGegmQ36PkMs0Fhb5QrJqoiQcTxyoFLBFsyksYMJri9
eQxMQDb/nI2K4kp3ZkL1H3IjZNn3SR93fMB25xLjRs46vo9lJ27Uurf7RWqXP/vR
WDd5jQC2YeBojfOvW13Vy02JGytIbLiwahZdnHf4ue3r4sxWeFsrAZhqa8mk0BsP
Z6mnJU/VMPDjrVge+MLAm+qXHdsc4p5C/mVoCxVKfT+W6BKvb63oA3bP/xVFYD/a
JhVUCza6wQiUrmV1WZ2WykkzyQqab6gv+MB3wC4a4KRnepeqlM6cIrKnrRc3AgdR
OW9osudRZaWF3FXD967JLyfYAZvghfoD0+Lm31/PcQV4F+GJb0zUml/M2SySR5Q0
ytDvLxWoWwfyXzjnX2LXstoLqnOf4Frf+jB6Q4n41HQAM9ptccMOBzzvZZNebtBt
5BGNyKUYZxOZ46/NUUZDthut4eU0dhxgmdVTtaRgn0K8nqhNZWCvqCkdfycRxZwn
l/uZtH0hDRnFq35p1VVBfV2uBozG5p802/PQPTTJgiy0GoPw6FmLcZJa9gbwo5Dn
okyIa8NROVfdMebLMZxK0iEpnVddtXg/wyX1VJ9maoVaQ99wbKTcohHFJFxfZ/HT
hJMq5BbbuhULmXKWPVxsw9NbfLSCc48OhDUb8hiOMdLZq1stYEmkVJ/PIjyVRnN3
52mAyPR9f0R0MdejogUqNzsnA+7hruNZ6zJizyOCGCfs4edMB7b/g7E1WM+UVJsC
A/4Bac4P/68RLDnWAHlrHVwT5IXehvNWIq2vkAk0c+Zmrowxy1T3ZhEaiHYY4cdF
MdpdsObDz8A+Y3jBIpT3/70cq0fTe8Tf9/4T3OSTplSOXoaPDac+6NUfNMsw+W2Y
71Umqjfr4dGbkkUTDHaORzk2YW+n8CIK+7t07DmVvP5kGfJ+9QpQQ1swwhd0Tewq
ZT8e/LHrXQBdbJn5d2ZVxBQn2eqE3hDFaAzv3Huw2saBMH7dcDpxAIFYeM/c9DvW
Ai7Hqlrn8PYwUdheupGafuVXuR0UwVdPOyB2fWi3c5yOPtZ+nxD8ohzIAzfgb2gO
InJ6mzk8iGSi1WhbJp63F0k064hJI3I64mZeHKemvwD5j0y5q9Sblqj8wuARSBgH
EBEob/UZTdoBNMbAOHTfnDwIMOaB6Cn8R2J0WqyaQOsTfWtTOVXh8gAtVHhN/Z0H
rQPo6NgwyGlZTjjdfp7mZ6MboB2SvibwZOKv8N2nmoCKQwIBK0PQhErNfr//1SgL
R5vmdzUkH8Yzn4wYvq3dWGGnUXfet5DcHkgRTtHllNHVKVTG1FxrwzjyE2HXdQHM
iqO99wbG3ywZouyc2GoEO3LpWdqj8qn4DMsOJkQRRoqX5u/ZcEltesARb0hlLvQe
+S4zll6eHhzwB5wumjGRByrLKo7AxO+zsNcn+cbkoo20JGGCTBFXYDr2+1oT2z0A
mu5GhAO1QgULTcn+4YkfOtgs54zpmiH3NNCXjR30yVZGLD+931SpKjuNxFJN1/yB
2Molb+7FoC480o0RopWjRZtgQ94o1dI/HNFTYEgjqD4cRxZ84cf0ucsm68omk/MK
sd3McVZzI2ATg5e6RryvELU5JOj6OXuXjxgDnQpLeD55d4HTaaeBJw9a16s0kcp2
A4Xl1Qxk1EF3c+NfFZCMVjIHkWzMFGqA+zE5hgC6k+ncd8spFTuaOmmu3Ut9X4+i
6ZuILyz0dCH1/4G4VqGdFIMM9LFmpjIOiK+ZcHeTeSaq0/bVfesFehSRNT/sKUoG
8lhdn+/1Yl8k0x74q9Aysw==
`protect END_PROTECTED

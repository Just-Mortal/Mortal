`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCpGPOZAcVC8I8BtkwnsU1ahzhTFNVyBvCAR0dlsMLgEEfaYiICc0kxDdHWJscG/
8xJt35QhQzSKeHgtar1pNtVTdMEW/Vc0HPyolsL9Nhy8dlf4iXOAo//3eMGR0OCu
WuaxCUHF7MTvwjVlD0Lhs4xeCO7Ph2MOysbjvCHNehAAjgjLMCEZ3ocS9+bKrbdi
Ircpqdnq+nwe9aTdR/t/znFo/JvDH5b95SAHnxXpUU4RBOrOcxrAXno167sYio4l
Rwug00goFmJZjO3OG88cuBuofudZ/GpS7pz/mD8iOPIuIDw5wXY44bZZROCJI68g
JPSKSr14AkjCLgLi3p1zDvHsCl9SDbHCvRjZo5ikCSNUN34lgSikUCpWekmuWO1l
Enxes1A1eW9cYfmunYRiRh+bSDGwghaYpx5Hs8yDm+XEfUymCcuy7vO2S1LaV0NP
FpZ82y49y+o1HcZBVQ7e3bz8ct/jnjfV9ibezm+vcItSwMR5+KzYtnAjvwNRnX5G
85ZQQenQbrGEIou2Uo1iTkQmPV23Kgj/shP409eZrdrSUnm37QgwRGD59U+Zijuz
aAg9P1HjvF2XuF8cxrvuac0TWPFRtXGEDE0bg8bCgm3DKa0F1OTdQ5xVP58bjt+1
/+MC4yD2e/l2a6L50qkCOczWSMzAtAl7MqJmsF/PbKFxhEjzvGrHPglgYCi/h+WT
YRuHENOXBxxicjVrgZeETi2Kl7L9oCYIQIozjzKAUX2KTEEsQPRLgQNg/hldIuK2
j26U0HVLFriVif0edjKP6HpJGxL8Zah6s2Q/8C2nWl8nD/hKeoT+Kqt2e4uhqzoh
PqJjjor8JflHKaFqtbbEf4YKWeiWCWypo2hsuhEnxIBWT3QhxH59EpFslVEOhDhX
hvSH79Oc2DKY7KamDem2p94lqDh5GiD6NcQEUrWCJAlgYBrCLm3WUxxw/ExvIoXH
rsvZbJuKhcpi4NWMjClYx62+GW/C62Zwjc1AVfPP8CGm+xTgFEdTrqLp/mhy8ccE
0FLXT2vn+2O+6bHeBULB8M+bW8t+jvVDmI5ABLvzXhNPJGp0UfN4GTCTK/Z2Rg9C
/1n9K9AGTZgtQuM3kNrbZVWBcYJNx4E2HUR1VIrMLnPO/r6D29y975oDoLZz4+83
i1qJGHWVAUcL4FhL0I8iiePMz43brzproEQjDy569eeMCTKA7X5070BDLPBIWpfS
rfqnXuFpOitsOWkJsVv/B04ljOH1UhToKOfYSJfL4fnq9OYqk7GPf20PY881UF+e
m3DFxRHbsprJaqBb9dcoC5u+MfQKLhOQWJxUZx5Aix9HN4+Vt/qvG4eUFXZ2/bID
vqOJWDAnG+KRaBO+sE8AakdEW27gM0xaRvfaPRYE3qS9NoWAD1ZGeNB/oto/PBfM
FtklPxENfkp4Hrz7QiOYINODSpENMXX6rJoY7M5FSH7I2qC9gh4sLjRLNM6E55UG
bj9Ir8tVOgoGuve73nnANDSM8Ttx7t5pAaKzL6WDjnv2CpL4DUDuWf0V0uzCGsh7
TZLD6yjaqBy3lgMCQ2V0EaN1KkYzFTayj2TG4K7V26856QKdsV0EhsScNoGbomx6
qY/Xq2w27++Yjg97WLug8pNoPeX6iTm4/7vGjiyvb88Rpaq3T+8lMP9b0vFJeI0f
3Zu+ZBT28w3aFabXan2ZBOJkb3NHB7eprHkSNC++k4i4QoKRjdqyfrgm8UuhO9YY
3oivDuvqax2iJxoxLNcMiDBM6krjn73mlthJUYwL63bm36v4u+cwBTdRnZbVxtUK
ulsuI2PzNJigvC2XKfrO/kd/mqoBeRKtqNLTK7UAjUb7hcz9w2Y8xKsQXzIltNdA
mtinOKS7RBWEQ6ns6S2cx7VDDx9LU/H/Wqx47rntIf8L7OPaFJjLu4tXAeUQILGD
6prrIjTbtvlMS75TCrn+vTieu57nn+UIC/Yyrwp5lxHjAZjACbn3eb6rLJNbVbl2
4Uyj5IqCt3G9fSE/doQid+ZjK1nwqAX60W3Rr02ZE2QEa+410Rf7EzGv6KUyahd9
+lltEU6/6c3jZQiDf0d8F8WkAKRxwC9doTWQfgKPkn+QisJ8ENphxYLAb89kZASn
Z2E0d/2d4UI4IrGluSZn+wchGCEqazLGz7YR+b07l9iuTKDX8eOkyPo6bDSdZi1L
Ncc/oWNPDt34Nf2Bl6pHhbJaxAYrtcW6g7t1NaH8nBk/6sFDFYBaNKFJ3q5UXIQ/
T0ssu+koerwDqw4zHmDo5G8bn43HpbvtDbDkQXecHgVjhLMlruk4iIRdJw9ustaK
6qFOsnZ7nRm+fwMFdysjp1Vijyc/rJQw4QaimqhwAB+6cn2ZF1UbJPYddiaP1RBf
tXPZY7Sdpk4v5E+n5Ns8ns3e1rM1lkThOVsAJ0MsPDP94pmsQhf87t0SRdQVYCXi
exUUvsq4E7Z9UXpCVd+we14+NtrHjtU3XwvUKJY5RmzqH+nR7BipFHEx+JkJUEuK
hMznSNQANYttmTVH7xM+bmIRMMZeLvf0yXPxxMVMjTLjzfpXsJuIVpSeMjOHtyhr
gj3ltU+wEPYOZBlH2ldf/HhSLk2EZj6H1TncX47FKDMeT8KbohuW3r9gqyG/9BVY
9wr6AGpIFHbr7i/OqmdjTfGGn9Ycq6RgaRB0KjzhXHi0MMliJjfoTYfmmqAy0gcK
kNIeX+FB4F90QQ61RKT/M4Ts8CUHxEQdbLdUAA9ue3eXNknA4a7fmlYlcA0R9aiK
lFoe6iBw91PCwlmGhPSWdH3wIugx9rFwDohDYnarjZSj3wQevl+UVo/8XkeQjU/+
suiRZoqh9n1tgreusyBu0ryl4MkMlIOy9KqH2X+Eheg=
`protect END_PROTECTED

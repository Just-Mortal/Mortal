`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ySXxd88+YOKKdnF/U2aikmysfeWD0/zzTYXhHS964NwXAQ1ZT67M+GvW+SWRp9p
c5lNRv5dveEUj1z81KNB9lxpsT8HOJ1Uo0KzbTRIAhsoi3ffkyeZlIVlz+vjOwPa
hb3Bwf1rImeOnb7eqzdiK9T/mEVkF8jQEyTaqDvWCg51/FwF3M16WIWkGQQsyJFg
pbFIZwgZNZ277nqNzBC6Jvq3T9xLr82tb/QNaLo0vDVTKZgjgfvHRQAwGHutsiMu
ry7luZjUmYVRyCU/9wINDXh9zti1/Sjuw0NG0h7GJvV7ZwYV+0eErRGysNqvLJ3G
hx5tGBNNjxB6B43rARzubWLQZ7a8A0/2hAcOnMZvmL9uXrhGdldvfmpWGD6iGKRI
ddDV/V5qDBd5fJXWphu0HgtBxwz34gj1Y3QeZxkwsk4gG0NGr1Xv+YAFJOPXVgJo
mPhJ1F1RbXaeT5reEpLMp1OVio92vikoRjbUSqULVBFVEDi/TnlGLauDUfskALIF
YmZpap8GR+f4oUUK1eSa2eIMp9ZQGwpePSMbyzhp1Oh+2Ng/MFZlx7JijuGMLZ0h
lASCqwLdPC75FQwZMxCQFG+ivlbocsnHiLAIdwU7ypDV/+dC+CupgwJ97UjY7LhN
YVi9Uf8ScgTwgBGUoZcaXj2Bdr/4kAuipWUrzIorrqVbIr2hr/YHm2t2TPsadEXi
F+qVr2gowvgPprm+cOgXf18lUCm419Puwwy1uz5/BbtJCvNFdLt/65v9gKIDdL9x
wRkYjdQSmqeF3ADVQzY/P83H4RjcLkrBiHXRpkUDoMVjY2EpukYXFqEM2QtKIudM
qdB+3NJoCz4/QXVilgKvGVeF7HWV6rze0vW39IWLD6QcOVY+pjIQskdIkJ/Q4cHX
Wjx5bHjdWU0ZuMWZJT7KxACCjZcxxeLeXOvDCkIhuVoKDF53yB/Q2a0QpJgjrUcL
ZK36sck2U/WY4xoxxX7aGCBVpoP08niM4PT55Un7E5jxhbfMuXJECy33QGJpyzK2
6E8j21M5clfkKLelfuUNvX4bFDF+rqgpONmzmWrPkwk9xrk2jYgPMixiD2f7vKGG
i2biAaJ1+60AfyrODCiBW3tawfd42B3REpMPmBncX1LwTTxEWv40SmBzHb5U2R8c
dDpywHAp3MBB0JG0bNNjUO2qELEijfC33yFIpOTGRRXrYr1Pg/5eNdY8AIzwqCuu
kOEcYRRRA6O76RXOJyqED2T6rZW1A3a2lKtrSV0Kg/VXTe8VHIt2dgs3jLLBX6eL
FU/D9BRrvztlkTkQJdsCOE2aTOUpIkZMFXfZOIXm+jOtEjUe7JZuTJVSC8Ki0Idk
5JPHTQDkL9QnYt6z2JYoMvc28IJ0ghPwAV5hHhATYYgwq3pfkYjqZEbGtfrr2Rvt
/uGzKoHgs2hcObXF/uAspT1hDaosgb9lLyyLK7sEDY9dPQey4bmL/cZDouGeFSBH
CztGVDhBloN5ZSL/N73erRnQmPtwCKpWoVu0qjg32e3F6u1KxcamJJHrwix10Fyv
qmOOTzdhba22Bf3IJvBGbE/o2ogzDW4f0qAwB4/y0EHEcGqefyoEEYtjjrtJY7+o
BiNQfvNRof5H9fzimfWwy0Mkftm8LF6sKQVRnMd2EHk=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+FcUeMt6Z8IKYg2KERIt/cD4yKnvmbRCcE6WwPznnaK3qbN9mcFkX5h/kmFS+E6
wJ5B9ACxXzil4ULcrGbmSvJx7BfCQ+xbIWgiTeUwXK8lsuEKXOeqJ+GnnANuyns7
GLKuBmE79H7hqZiP45BUoSwlWJiB9kxNlcLxeiUnu0jnoQQju3KmRgcVoRGCuV+x
ySUVmdfq23EOIJ+Dye0dgziSe21xpLUw9lRuC4XlRHmlIIpql15sE+HWDMLvRMbN
lMWMLSMI62p4YuLIzWom4c/QYNYz0c8dHFW1AOiNIH/oIe3fzqqTsSjwY1icOkyJ
j3pECYoljKH380m1Z00vrRrdg1mbWhutnfBbaNYq3+to7IU0yo+EKRLrCMdv6m64
oKaitqqEQeL6xJP48Ir0X+fwpmtOoFt8epFB0XDrByOLCRrOPEIYo0r+Oc7LoM+L
xoea9xPG9H9Kv2YsTQGKWQByJ4mgbcO6jmtpyXHgSqL/8SquvUDBO6zzSM75/NMP
dEnLs0V9W3/YRfOA6jnT/DpyFMzq4kqztgyRlmbSPnFw6AM3AFPVHDcNyEG/lao0
A6otTyhYFUhIuhLWc6Uzvq/LEBkJCwhtyrThEj+laX51FE2FvGDEl6+j/GZ9BbSN
MRkM8jlWM4JpUMCEsznxjLo8Ua3FGl6dYxf7lt+Uz7N80wWrOJ41sfo2m/UyBkLU
sltXAsQ9xTHPl2uoN9kMlPbULq6htzNwHJ+/blcKdQbyRKF92vf6ZkKdUCrZT8Tt
Wnt80DRX8GnhBg+ZG0UY/wL+q33gtoJ7yLSUF3irNY6KKyGPG6fFTbaRqStF3kZM
ZzpYxJyZ9QcO0Uxyz3iR0kPE55xA1CtD/amta7kPoisqnvQ5BzUc2WHKbOagq5rH
0/mjpFK8FXn/6cX+FxYspC7PCVYiGU1KjeGZgcSBPQBB2NfoVX1qIWFyQhYVuM62
Bgb11eviKSGzIUy4dfbellYtf1Y8kSXqqvoSITGqL/reR1HgGH4HUlIIw14k6l7/
hX5pgP57kubQ476PHHUgDE5UImiOpDl6CaQmE9Stmvq7Er6FHMGsmqOZzeng8/h+
pHACyLicfITX2YzMCJAFyHqUYYu2Snv6dUqUj/8v4IMkkrCcPrQNJYyKGERyoC91
m6uHttUUS0jeL1+vJhHjOAvb3RTrYHtICdJfVzksH4pk9u6a/LgPJf2e5T9uNOFG
hDEjJXdmeyXTd7SgOmRl7gn/9s59RZ//wyzym4dGNFmLYLTWb5hF70mTa+t4Xv8A
F0BcPNZq32GGc6fULiVZGN/P+5nQ1EXQfP61BClGvpkt0bczQC7+nBv+rs/F3Kqs
baYPdV4Q0qkiGU7RQif/S4c33/5hd8XprRmqitkPXudUuXJcS2LuxWjdwg+mmHjr
ZMhvJ+xV04fxPXQZA24hQxGUYzBgmA09wzZo14DCbSWE6WI9T4eRNDAdbk8OPBLd
lfG2Ox2Z4EleTsbJ91oZLg==
`protect END_PROTECTED

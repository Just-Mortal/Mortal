`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rU8skmNStLMCytL2Fj9hx9Bg08ajcQ+n7fr3HGp3HFlVmEiAdfi7XffQbTD1Nm5D
jO1JMaE+Zg6Izc1UQfTknygtjEQW63daSULr5DgTwXNL9w+NPmtxHWL0SdSdqkZd
hmd242zMUmqKoXrG3cfkLyndJb9jzB321nIr+YHDAN0/CdqznpZ4I+mVe7MIu6iB
UYvAnLcLDU/1F2hFND19iVcq3ngbhQVWe9sUYwqlVU/ZLoxeU0VHznE7ZRAo8Ubw
lDKqYsajugxfWkpRxq4IP2B+75A4Cjbv4O5Pw4Hwru9JaMNzCXLjiLl6/d5V0H7I
d12qWaaCPxY/0CsnmzwHqwAYwMmXX5TOiUX48H/1MBDpqyMyVBA/SY0blpQHBSkw
gP8wkMseudp0orWfPwLbSikgKGccskUcJG7nQCxfzwuGhNvvBMV68yVetFba2Rhi
myyaTkXhgaYKrZWV8ZH+pKXrQv1jJzz+j7k3NsycRK+PudDZCLaPj1M7QEK0y8ML
vZeAN8xeo1BF/MBRmpJKDwN9HEUvwv5i3ebWQguo9xqzcXFWGqWLwvO2lJzzmGmW
Xy9y/nflJlDeci/upqefFWpH9GVcFFekLCLcWHWugq2BkRY15wjz5dmVTgkf0/LW
KhOoQBliQnjQI1ExYlNB6XMsS8LEbXqPH+dVKE4I96QAmKm/s3QD7XaEERpcES9R
oEKzYTVl/fKa5CmYfbCU//iTfFLdS6ikZno/eZBb7fY8Mp3o5mA53A5tN7hpfvMA
ey8TtL4IUFG/JBwv6YA/V4NUcg4NwWCSY2A+5/Jjrylnnmo24ZamKxB4Iht12EY9
dk9cPlmoR/bfLNEfDIKk7xQ+YLDN+qNmJyBPMKffjqXY8MVmUIts/pSCfAitCGZG
GsOxK9/PcSNFWvcvCI/T5tmjr6q1phmRrwoDiQCdMno=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VRXdiC26/B/alVLo2B6QLczXBe9ti8Hg1sKdfmVIxc+gAjgo0bjuQOrs/LYrP3Lt
RWtMNofE0gruHgAhZkATrKlvvOsWEezz9ZAl5NBIxeCaibQQwLpb+c9oVPtu9RO6
S2uHcfz2VyWMXk7DuUlCH11zYoo0xjTcaSKcUy6J9czXY1efUyA/6+yi2dGZ5EYr
BHx9b2ZtOyPtD8ukkKqysBFBe7PqNXWxRSjsRtPS4/wjy0+NrZnjHeSLUbToOCjl
EmQeD4B3+PZ0jHZVtbfnrhDD/okJNCfZZLUO92tdwXSV7PhPCfdSi3pmw9Cw9L3s
FokVF/HO9xSo4Pt3DYc0W8IcCwZNgoMCZexGy64chMrdDl8PlaiAHU41S+7qGbZp
3seNtV2zVhCvYWhJht5+Qh0e6Zh+cRvgCUnX5gLwAFHRSIItQwvADH1a6f3+q5i5
mo7AFWkoluxTqPBi9nT5HXCHwx/5gOVWLFmhwtYcsklecrY07qagZoHRuKzvmh+A
HjMDh+C9OhskQ5iWk7/HsQkanuHnIf8qzo25RvQWI4prx14Z2m559XW5XHFeRVLl
a+xPl2o5YbXSH4B5r9brmmID4ke0w+0Ec45sssh8PUmSq4yAUFsFeam//33d3M1r
olb1dxCGUZGdrGXAw5q7v/ZlkUOnFqS15EUKhZP2D+X5X9+w/ExXj5CcmZ1RgIP+
B+sMafN6WW0CRrAWg6rtlADG3DEDOjs1eTuD5zJQJvD9/atpW0/2IgoHPCQQaZGu
/dKn9WF5MXreaYthLYIBBwG/ukeHIetcMmlrbPnzKKBJc9wHS1oKSmJwGlb8acHi
evqbsJaSduj4uOBnfSSHj4yKuM9nBWCQDNRGr4qIvgyAFetI/pBRI2WT984XaqXt
/pSaT/kNZFAzRXPRDkipx+krfsYNPgj1l08sBrHeQWCbstdAtS2fhy2hR054r6QW
5iu/jtThI9aw3Z9g+ckcuS7ququtMfuO1bzEj8dHGBvrsPf+KdtnPm78b8ktuqvw
b5jDyDUwPd3xkLUGRfn4TsL4OtDBQSuHNabJ0u4XpLKEgy9OF8HQpsaiJG/Zc1Ch
VDeN95SAHIkV79cDmkIZVMYcLg9SXEebv8uZICMXmdyD7wnxyFbw81Rz8FV4/1Hu
/Oz8aqNePWhKToU2VupQe91K6CPNDMkVKoviqB09wnOlSOLo/B20VVQAptvgARFH
0BI+FpM825yoHURmoMBS40/jsvdCa07kfPbRw5VyCv00MpZKsZ0rMS31rswhCeZy
XalMqxbgbTDmQDnKA0e816RB3DujCozMCIHx0oIKtM+9cMbjCJwhGP6q2uTYVKl/
ltuXTtLukvY6rKvjRkBvyeRJck02bzRN3+dzyZ9NDLiDutAhVs3jkG3Zlfb5AsKm
9Z/mmlu9aGOx3gIryuY7g/TS49qDc0LYleENDvqnVuUElT4o5kjkqec7r8GPe2bD
KOKBzeQKp4LRaDr4FP3HL2nZK1/8HIYVO0jPJeADA770/WdWQ1NRB00aBU5YnkMF
cP+3ErQEyGVbIg5FaOBQy0UtNI1A10PgX2ZFwyKuABJi94HtHFmSUeblHRDxNJwF
FD2J+PUMK6peRMR/e8YxZvFl2chqnUX5EeB2ygSuV6BqhbKUNjAE8Zo40MFqImS2
f5G3XZ49oft8U8HYY5kCFV6CD4m6Jp1mIQ3hZ/irlHp94s535hM+MXbGZ8ucn73W
9uDRr9njmd8K/36MoTUj5vnX1fT9sLfXZZVaOOMUeYkOtHTioe41CnKflgpP+GSg
RytMZvwFpZbpS0AikCQF/WgY8NWDvSXQWvrKwOIo8QeJ8VdRk6Ns/3pCuzJlGQnI
we37ja31c9UqBTm4unKscrISfqLWekUyZbritMYtnwwqsnk+XQxTiLI00tQbEnL+
GLngIu8pGZ5pI+Nv284BG67VgdrCJ1EExSjYi0xD8VYB7HXpps3PZqbmXSVt+zo4
sMNJAn+W9Nx7lB/KT7DCniFHtSaxwHSU+jFTzSHz/i1YbmGom2h571vBiDiY3yKt
EIzPfyVrtVwWilFr0x9M4eOtklwgddJRKaH1Kx8R3KwgOFiHvvZV5PJGfRxlSzZw
6xf5QJkiJxL7+/0Im992uHI/2T7zHrHCpm/5Aknbdv/OC5ugV0oh1lVlpsOCLeXQ
CjcHsM483BRDsaYRi/nWfXh4i/cX+9A1prlYWKKNYlAGmuDZbJFgI2yy/slN/9Ey
eq0IIl2qMefwABfoSzFJXMsHSx6JQi6WhYIYFfNWTyanixN2hkuyfUqy5LBI7fdd
XoUDkN892mtCGEhCGtSqpktIe8Y8PGUV2c92osVLVff7tPq9RaM6HWK1IFrp2aFY
HWXLlAhexm4nlipC95xJU9jOqKs3b8oQTQnaN75K8srEcqPIoZHmS7bfsj8FyCuG
tBddEDCCKlAfo9Tds+xghBoHHI05egiiizzC1vHVAwu4dJeEZrHAjCGwZwaARp5S
FZYXGFer9XMGikkPfLniZQ37aFOnOpzcfYEzr0eA8BYVH+/u0HkJz52S5rLxFnPD
972FPbRCSPBFw/nNWlUCRYhyiQOzjCI1AYSW9sc99Tvo2xvO4Ol5zl7DGBQHbB0D
5xJSS47Je7fhz2/FUp+V2iMD3N/7+vrNAIn1mHtwMIdcbDeCuXiHr5oHDuOicrWQ
1+VATda7mlKLUz1hDyrBELEo4QZ8QPvn/3dj8tOMav5bD30ulx5Pz6VpYPYVVvVm
Bq7mxAozxRgWpw0MYUx2BtAP/M4Nm2he6xusI75savhLYIA7eVLXvefSWjUC8bCt
PztOgzkibP5Z/j4/taAq3b0hPWn2RUFn9QuLthvpK8SH5H7tkK99VyYbqSpmfuE1
vT5c63awTNbiXwf1td9aQBdspJLOxzgxZZMTwvKp39dlozsvc0Ch77/Uv9UrO6P9
UYJIqT00ytD5yC1M+n4pBI2uD5rF6ZQ9gNXVhCASCOlIOA5qyywT+ZHbdgHmuKKS
F2ooKy2r1ru+O7UwdxDGUcqYAozemGqU1g2PcnOnIKputZeMgyiQ1nZ29CT6z+SI
tYMlYMhbKca7jRMu8D1BF8lqAkTc3XpglZt3VGK+bHkfNUUKdRbsRo+0tnnIhITL
XN591QohAT/7Ij0jcNh2OIA+0xzIl7YQ/26mwovm8BrXFSVKGAziHjWFCVszbGZZ
TekATJtt31CM+qEI7bdZHo75n2T7ZsQuakt5ur1sArFhtNcuqiuucW+iquBLZ71g
FAHBfz612hY0QSCc9j61FE6nx+KY+LNUyPEcaZgzeTeM1uI0Jt9HL5cVunrlhfHO
Sc0EnymYspO63nPLn6Qa0nuXJLOkE7kJbNjqlSW+4IfxbeG9E+O5rMsdjcSMxVin
yXO/0T56U1YpYPi+gT5EsT29vjJU0E30brdrWn0xcFDH4EOZ2QfY1MnrQapSCf7d
EpedxtFB6C/voVuqvVBVjxHos6YjaXylAyoGYL4TsY7SuQGhlm42fGxRQ4IQOFqK
tZ1bmGUO4AjlJT8d8bpytky12uaNVWA5BZ0XvD+VUuLOMcJb7EcT4Mqtu9mUkmW2
fnv1GLj1sPlSIyvqUR+aIl39C9csZNtKjYG2HFSogX//VZiKDUz6+dVQ3uWQhgyp
OVXIuIkVEWSDae0XznUAg3UUYu5LCFaRK+bapLjzQQB9ALQSoMNiIUZwioVWEn4O
2suk52MUSRlALJNmAOB1lv8M3Ml9JHaUuDmuwIpT7XQs8yjQn4Ug1q6RxfLkfFdj
+cMTd9Yu4fwh2P0kqswJgDMIGYcu1Shh7fTAUbYchLEMOdNuFsmjsVKfdCueWhnD
Hjy/UF6JSUO8w9WdldEgZh3N/M0DFW3dN34j3AeqKMSHxg+TCbOYh02ec602BWwb
n3Mive8ktwuoPZcUEjeWqdWR6+f9+cLllsCjZuuV2H3pWQYwIWcxeu8+UuPE6eae
C43i54B/sNR8tcuXNLU+APgTai7WlxNoLgXcJ4pRivhMuL1f/FWhRKj1yvc4kz+4
ThXrta/1r/4zrSpf4dekMiau7QxvTaruW9zBJSQrKCGHY2TzcrksZ3utl48oqz0a
71t7jomtx34kOScr+xPvzvR7ycGHWd7vaDLVy7M0tA1t4aW/4itshdOd1D9KmNoe
cA8B/3aWPk2ngY7y52n/9S7i1kybZ/gTK+q3HKPHQ7EHVkCguQ2ULFkCnptiCL0Y
PmLffoHfvRj7wThZQNRWVfz6CHzX0RrsIT6YrVfHXNStwuz0vPYIzLXOt8VB67Qi
UuaKUsXU7lvTgabwI8PtRaJiJyC1kTYvpcg8UB7S/Jc2ZXglxNp/sOrigyjZpy09
QqPIcgF6hBiNr2qffwHj2fjw7Kqh0sSmt2H7aTsWeVriQ21BKvu7BzAGVYj1OuNY
pTwB89c9wJMCg20dsTGrLQ9+Dl5Vhis3B3UR9uprsCHDZNNTU29iWskACU0lEbov
Z9i62GDfoHpH1EYvyD/Pb04QYCcblgq0mFZfPQTiK6kAnDJn5M7ut8TXboyPxGUW
Ji6EYNJFiiQLP3CoyAH9HOC9oAbYkeFfVL2CbaK7Xgc4oWXpUE1QL+6pGWXDPcIL
vlvH9ZvQuRI2g6Svf7uN5kBo4L9vM7865JKE8msUChDa2BAKP/bcZcu5pm+EyWE9
a/pwadpuPI43inxMDDzfPbygybqrO/5s18wOArwjeU4=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eKLAJh/40tlUtoQCmA8qw2l/jFj8rrg6iQ9nrVTZXiG8Lgy5C43SgBiEIIRbfqdX
cR5MqWCjDfUbn+vUHoVDkVyJzoza/3wAucxyBzbMm3CfLkG/s21gRZulK/A8akBR
FmwbEwETslBFncH4ELbphdBJqJS+rVCES/2Uph9ACk5FyrBUuLEdi8HTFTUH1YmJ
muBpfuHxtmaniAeBdRJKgmEZR20xIHkMrFPEEru3bJeQgq9sDen4wpBLjgxZYzq5
f9wzkHKeHmbjw1YgEl83YfCTzu2ctH3q/IHI5HqmZnD/Qt59atOc7wqFx7JFVwRw
xmItpIKOEivgoP8sysUqf1ILRTmzHsH5jep6BtZ1nCHMOOHP2w0z6/KiIUuKU4K6
Uo0Bt+zz6Hx5lOVVpjAk5sbvIPBSQWlbQTAVMQH4CluFdFrPi82He4GADMfwQnnC
G3PoA8JvWS/4FiF3Wpj45Ucu0ERPqyDWvuib/DI7Rt5Asm/d2dNfvnrh3oCz3CnZ
Bn0KrGmr3TieQhpCpUNMV5Nhf/fOeD2+c8oUmyf1uLvJL2byNu8vobHSOLEDOIOz
MT6QAh8sItt9AITRMRHfFApgO9tXkvfam5MO59r6jNziAFAIMtDmWdtX+1WUdHZd
Sr1WRrRWpC2wtqyrADt8eNYp17gCkuUShxF/3l8qngdkuOsCrPJvE4wRg3f1VTwv
a5NyTSXuSaPEA6cKPZX4380a/e4DiENr5IVRNiDPQXNAvhOmFMZHrC/jR1yD8MO7
YD9j7acYzozdAy7UoRI8h8rtaLqf+TU2OIr9dgCdmBXUoXP4FinQqLpXRbU4ZPbF
EqsRkkup9GUITrw9FOxf76NY3wRVKMtrg+hVb0+hWClMBw+X0WANFvzXhdlKEXEb
dom4pe4dUGjpq2mr778SNjLxC9tl8m1/CvGfjymO0USd47CECt21+SeYdrmOJDoZ
Mq1+5ojak/m5ru+NRMIj2olUw49zGOfNcJHOb2LRp79GF+8ldANy3wT127pzj0oi
YIOLBv7efBqKWHckImbeS0J7/7VoeYOnB3uN/cWPcbxGzUALrPEj4ok4ij6uJtJe
jPSSUf5Vq+egTHuusUyvkwYo62WCMgdSeO57MfXtC5ln2fjfiYEDmkVcTB+WI51Q
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H88rOIU4kTCdbjx3XttOEsrfFoMJ2PmjIxNPXgOHYAvJK4dciXPUBgEs8xnnNGlp
dTwjB5xGCFxLnlMLjDuP08jgUsZty5mrOWQCkVlHEKSURbB7ydO4EOi+ZTn8veHV
XQvXDKvmq0a9j6KeR9cnqv8FIDPx5fbbadeve5T5JOvwVKhLnFcNsK/d+7tkUADT
d+EO9Ko0bP/2x/aN3BzDLxJqw4n8tAKn9G2sUZxY5pKOKWckoInM2XNvnWIBTwlr
HHtXkdS58APsI4OMZhbSAAIa10Rd3Gd3MYRxaLyAyUa2sEXLVMQRVf/AmZdGAMfV
/j7WsRpv0yiU+sdFe4exjXwwMO9ReqU/kVQH1cUANsizz+6LJ4HsDJzQpZVGg0Bv
AaUK4OyxgXEzOH+L9kPQo3XBcTw0Rq0tfJqR8nvX+SqJYEioSXGhqacjNwUlRQ3b
GIzje2qy9aAvWnVW5Xs4OzUZmphx73kFM7C7zuCoW1nON9RZlOuCtg3qN+2M+m9x
uVGBkQ/eC1rmxOQOW3uS0+eKAoNMCKv5XYO2b7iYHEsfk79e5pODxbM9GJk3XBaH
gQUlhdGvDpYFepstwa38MQ8Sdhkjs0RPFtwGhxdbwfCK2n+KMLPVS+XLpQkkQWYK
h8RgNsOWd97JlZ7rKk8XcO6CBrx15RaNzKaVpJ47aqAiXahceiAmMeb2hsWh8dbR
L2z3UOJyeK5cfNuT5S2wKjwCXLroEc3rwTStdLHI50KWdtaHR64q+p/pEGGW/fLS
jmmNz695gd2Tdt+9yDMqYUVkIlyeBCFeswB7cmharF+hU72wb4nXSiGN2ZvVuQoO
FgwhG9I6DRlM1kebsv1dvzBBc2U7QC1m5sqAAo82lWJHfqnD4tQXJl4PppgliC3+
062Fv1Jf8bbecBRHUMStf6FP7d4uU64mFbVvxLZttosqEcZroghGoIro3zT2OL1B
747rjIuskax7jfcWFXfsXYsOx7Utk7/cc3HMOxzn5w8TFFtGscbEuBwVzgDtP2CJ
qC/gnbzhbPLg4tIig0j+dOa5TWP2RJNLIPRQIf2HbLyMCbUcAvlXPMfeNgbA3LyK
S5NvpzrMW7pwd/ALHvzQAKMbjhPWZud52eBtALOnt/um2lN7mHkxwweBODhcPyBo
YJMjuinhLf4gvIQZC3LB7sFhqvM9V6E3aHy8tZlKfCkUTlvC4FWOWEtsbMdYqjhz
0ROYoVOHRCg2ryYuQBzesxADVAKM1EsYqXDRgfm6RcxmKm0UMvhG30aERdPIDuvn
OBrPtasnX6oT2pW1f7ZLMUEmDIjv78Z2f702wjbPnK5YCPhJ4dajxgXJeiM46Z4Q
agNwVkebfvvVhkM5MxjI3XjCi53culeJYQ6VsaFW10UbiWfUhdtdfkOFL+nzoLoP
kDIfHT5oI+VXYwTBD4AfLTLs38579afOAzrLU2YPrt5GjOTphRTFGrzG3zMHB7Io
Eus5q0OHUnJHXwM2QVVnHWjAEORD+GLIDKUPqsxzNL0NYYwOCfu56STNoDQkVHCM
xfsNL4qMfAPJWoCBUU3a7Rojt3xpKkIrTC6iA/m+ydUG1QfYJh30YyX2S3051LBj
qNplVf3pQKQEas3ndQW+r6ReftPy5KwuLQy8VhHpdcntc6CpB+7xc2VXNqTu6bcy
AgdwirK3vAQr+/S7ISJqFdDRDfIwwjzbOxawKUoPq8bkQfkuwQ+KPOFva/RsTJps
4mqgK7gXA9KVvIK/Dl3+0TwCxhOCrDNJyYzLS02naZdRhZ4iADH0szPnxxdH6HDb
wy/KjtllGDjozNERii/8YHYWCrVryRJMcoNmvnAwe2U=
`protect END_PROTECTED

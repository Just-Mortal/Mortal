`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWGjYqvLbrW+DE2afQ6DcsViS/SIEmjlGKZ9ZkLbVCzjvEfFKNCWNRluBeaQwzWa
g/e1BXkR7odl+olZScYghU5waM0QK8N9DWvcmZ5OU63I6oik3uhAeyeX16erqWnv
9tEfB7Op57W//EqOvPS37dCEdHTzs9Kc5PQTYPXzRVk+Sw84oWnO6mFrjho1l04A
naZb9lAFJ60/9JfRB1nKhzNbcnqlZfk6iGmeSl4L2mDNaezXNfqCiEiRRiUK5P1p
mMefm1kmxS/o41xrtxi5DyqSl0OEWL3eXkbVtzDiyjl7uRUWjP/3zYypUJExGssp
LwcfUahJa1srzscDCciwRsKEqrh2DK3CDUNLKLsab9DejjSXsS6Ijy//xqplzp9n
xhHxA0/kEcFiT2yDgJstNNyOThNuXWJXyHkLSddTxg/GgsSKqsKjQXfYBjpxx+Zq
J/gJMyixhKU3RGD98wbKFbObngBAsqFbnRyPJbKDThSwysyPRpIHFL8vbtwEz8ik
KaY8R1mIr2dcSAZJLUyyNLzi451n7InKHHYJ05lXLvh5T63ylI+2wM207i4dx+3s
T+75+G/ZOaQBgjDa/yY+gGXSdomWIMjuzx5Wtz7Tcjcfl6AAfVpK6TIuptcXZIkQ
9VvOYeGX+0eirwOeSSXOFhhpZfnEkmhyT1OO7xQMWKMsl3pXty7EP39Ix8TZ+PPr
BbRwHb1V8tuIBeD0YOXnvYsKA6qsoYk+27gfezdChJaLICTFDpMsoN4WWceoZ96J
kdF2hJZ4RTsmXWxaps5qR4vGrYkI7rvrhV3GxQw2WlOHyse+ojEZQs500wA8UR12
G7Bq7Cr+FCPgCmDcpw/K2V+mUHVHFVy3ckI7eFWqJrPDv8VUe7jfWvK4Bi1cpa/z
+v4JenvWiRjK5uAlhDtFS81L7hZlPByGtTlJgOts7FqanS1rKM4sqolzGOJV+v5C
qm1BswH6hOCiQYqdmlY8XYbVqVmre1pKbSJ4tnTAzNF5P3D8gQ9QNhDAKFXRQi/R
yxSBceOaeP/dEVVCSvRM7MyXWgC85kisksftPT0UNZKSUtIJAVsWsMchLw0vyWBD
VdIYaCRfvNwBSzSV8U/xRZhciK1PUtFL95ZdeRtw5VytvqcVHVpIhRN0zyK9s2lC
OwKa1KS2b2aq1g8zCh/FaznHwghHrgQkgDqzNVo8Uu/h+zeBEv3oUjTwxcQXvpc2
Beaw1UWO5d/SAWJdNMfOBZIp9/S5CODbza2ly7oSNvTzkd9p5IyFeAvunUqIUY97
w0MQHVfHuWKArLgytdpGsODc1f0BPYL+Q6R1wSPWdS3ZNVJbYs/VGe8TzY3RrT9E
cVck0Kn3k4JKCRKv7cm53EbwJdUv8v0pQucpjEIjMEHPbF4rWy1FBB84FyAioZVC
xONy+U6xbyfgtMRMdFWiqVKDVK2f8ojk6ZQqlNUjmd9fp9pDXG4ptXhfCHUQ3n1A
DqnplFFKp0pG5kjVqReBzSAVEgw3Q5WSPe6WyqRQMnQl9dMrpRVwNk/95cPrE/GE
mzEkT/JagOHURBICtms5QxHoUU3soZxXs1Or6mPnGOnsUgcHmo2RNgKJhkw0TTB9
Z73v6SpbWiylgev3vQS1JdvRhlDmnRK1XuV9reeMw13tdAwRfqshbSRk94FBrEcd
DiRKNJlhGn/yuB5IDecPt/0c5yOzCZ/eEdnJD8QDu4372bke+oQ1WFmbLkqOLwpk
eWUvipnSTUCJGGg0D7mcLeZfYrDJmPzHWkSZcj7eamEuKjAnkNTV3yiesbpaB7R9
JRrw8KLfYWRcfjvSJ6CKwDeddM+birrRKmoI7RcA4kkxc7aFLO8WvyXAzL1a6SJ8
2AkTRJ8/eqDYAQz1RIqH5dz6ZFrGIpXIBKTQ75mt/OaVT8FWMMfOvzfP0YHp9vYJ
nvqt0JCdZY27g6xndPUx1vZ0NqySfblbhq6di+M2wW7XH1PmrR1KVyvTnbi0nNga
4rv/DkxFcYfQeHEuZx7jHZTelIzRE/MGqa8YHHYnF8dRIIMTkdWpt1IXOceRuJBb
fSOpUVoyPDjdu9NhqXXHsTME8bc01sm4Go/xZzEuMDGlC4mOTLaVEa/cLID5I5Z0
8cyeqTTKmTgaorF3r6r5UVM5RCrHLXXA2BsCPpLczfu0mieyruJ6dVBSZPlAI0KN
IpLLVRxQRInUrV2i3vNF//TrcfeF34VpFRzrOPzXq+4P8jFxFYAe9AcVU6geivym
taahBVLD47ZGAVZECHRri2GvqTwCnaTfC/0nt72tjHSERH5RhjpDRaMDHzCLg6/k
HYzNqOlIJQMLyoDdD4KDGuIBQtMUtiX+TLQaQ6YnONE8rebOSJar1LS3Qvc9j1Yj
AZRpyWTu0J9XsiQMtfENvfFHyc4sCkQF/1SJSwmizb0Ijf2VySfYfUdrvE7a8znQ
HKo0455FofukhdctFtRhefq60ujdyk/mje9AIIw2c6yRCnJ5cjFjRrNUnw65Y6mY
vYuGv3jESgeIFdgLmHcLkhx25w5TjAf3UlLdu5gt3VEyKvXeLbthMNzX4tWP95g1
v7Awqc6d/4Jw9Ln6fHqnlPy2GFMc2k2BEcV4PSHMsPlX77pRUsw1guiOP3ubn+Pm
uWdLaCoUVIaizFcZY+wgPGk/DBIjHcGENeiXD5T8IY7J6hSFaYDIDGedlUTjgo+Q
WNeJ7AouOOsxu1/Z60PhMhSJJ06C0MIw+u3CaQACDmoQiwAzn5w5T4nMWbfSoIpE
taspbF1CH7qfQNqKneJNhQRTrhoCyo8eDpfpzkNeemyiLMB5iF3AWFDl4pjFzko+
099QVToBcxnI1cnT4vuyjJCHRkBBwTcjUzcbxFQsunATO+XXdlNTnqVnhmdxNuow
xeNK0WE2+3UcM9za7/rEWE9S4eVUHEMZIcjKbzTJH1vyLrn3/Rx+d4clXtSBa8Iq
WnkQ+vJgH62hiaT242yzSKFiSw60ryHe6IP919moFd6NdGGfSwXodyS58HrhWRRX
QTHPj9XsUvy2Fxc4I1BAEgwDPikFyIp83KY6HJc+qE1J40dKY0y/jPx5sNrWwEOW
wqDOygfsIahkFEGXu1CiQco6q+4byY/8/BRaGt1oeapQ8OpxomhmdoAC/Yd9dvWM
c4Vk9IkBZmvmupKgrTLaX3Lqj+1eikLkvdwCs4QSEle6l3g7xLHEeQ5dM2FwCtql
m3SCIwUl+BythMz0PyVNaO4fvBW4G9ZzH0cXxW/+XW+iXY/IVK+f3/MkJ8/1Y/Xz
JdCRKf62r0Gir2BEHDY058W68YPYMFnfG+0I0EJHlu9HZfSC4UBefjlyibVC5b5F
U2Q0JZ0IoMkBqIcdO7bTJDVWWMnJfz+/QlsI4cUxWYFaFakqSUHaj6/qTowSgS3C
eDNIxsPj64fxIOo+jEvC9iRWylfPjPs27OZiqgA00t2KGirnh8OeB9x9LdZfrPlO
MKC+F61zMjFPV0df0cyCkWdhgplRbnLzP6/EUT36AmjNRROwQ3/XzoLmZq94gJMh
6SA0FQh/ww8+jYmKmN5BJmRTw2/j1cRNYVx0w+qauBvh5ZtInrk86iH2nIqdei/9
ZNssXrLQpxEJH+0tAVuxPvKOMHwLf4gNwUxn9eUD4udhOQCWi79f58KcYX/EVfCJ
kYjj8vIJrx+gpiRzvAyBzZGXIz+Dre5JCB2WxScw5G6ipbcjJtQy/Kli8NrJjU3R
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qZzZfzNTso8RM6SlT8PBg7CeeAmscO48F9A5bQROvbzomHN/4UJ4TBGE0G4kg1r7
ifAXvcZrrkVf7U6FhZkL3zfcAPZX05ABsBTwb1aHUwd+JZA74QDUjzd9yv9NSCnF
whhWuLu/SL76fVRktYZbILT990w6GvcYsd7nJpoL2+mCjj1sekKALpFpZWeF4Me4
Ye1Dxluc8L8Nqy6tdiQvvs8QpCi2qyLEMz8Kgu0x1wt831NCVikv7SH/oJzVWO7j
ZErWPqV/eM4Bir1S0X6lsp1bp6Tt9hOH4dPgKtYRpvBRjpkz4D9l7rVDlXPcLaEZ
rBJ4ufbirB6y0pYLvuDtoetdTBzVOZ5CXDJJKV2TN/nr8pLyO2wXTiEs53WF7NQe
6wwxLPOtC2NZSFND9tkUl+Gu0c7RZhjByScX9JjbJf5meMWWCKLuG5GeLKDJrJ38
g0W9Z/FAdd4NcsVdCglBNGjqOVG4VF+5ia9lQMNyWWkyRG7chsluOKDeKZ8mg5zn
FdVmqQMI+gmTd5zvwgCqVpdoR9+cWPd5oWmSyqSY3wBlLsXBdw0fCWNTMNv60hXM
/0zK30m6cOFQYpIUdhk2JOgHWKUTHbXRv9Hl983dil3U9tqUTH07EZ+kzVv6PfQX
pPL2CKwUANI+lFBYBhLRFHGtdtmDjDoJavuSHucSLhtNOZvtl/N+P+VdN4qIc8PD
noPtCQGQAuS+j2SnHJbZoIvSKXDE7g/WG3CR5lj3SVgEoe1Ph2h2oROlb2sw3tvE
2lYq7s1GoEYzfG3ViAHxRLiOf3lD76hwsX7Y7jZ8uvi5FR42qoRqpauErIAuc3r7
9kY1sD5v6FnDMLfJ27yVbm1tbyoA8h73YYjhrBzQBqjZQS8jO9EYeBUm46FQfLcf
LwWTCOCbLKHMtf6vZV6vorXEhNyhfSDGciTydvlTycfa657hUeQ6igk/E5NXMPxb
yaVkvNaNf+sAU2KwAuqUWKgb4yNU7v7GObqm6MHczfU65IZ2L8U7/SsYwjK3zxoF
gb6Ka6Tph9RIz1feK2XrmaW7AzaNv8kAys/A+Kx7h/FsR3bNdTL3qIt/XTduv8Vg
EvCQYG+7scQXpE/MVjEMWAvoPAuFQMYpCYzPhzaUWgX4nMsvcW4n6Aq7qEka2QOt
HvyRmAvcbHxnQeNm4OuYrcaCtjXec4U/4mBQG46KHTLRUkepSFG8NX7BH3YfD4jl
4SJetBWEpcVNQH1Kw4dlD8InboX5flRFO0jGpFnTiUJbLyatekGpN+i0NcNXj4bw
xOVe/4Vu07ux3hKQ/XAauiU/MqJghe5Kn3ybSZAqoT1IS/ISQNB9JN9Jl2kS9ftr
E/4arrDktALMTEk9FsrFh3f4lzoeh/Z0+3TUBCqPqlQPNZrxPLPbV8I4GA/pVvot
it+3xnq4H2fbhfTl3/e1Y40MbjuQi0JZftZ4Ttd6MKXfeH1mpKP+g4vGgeScuHHp
wN69oWd79PI1yZncWY2KLj6WS3Bnu58Go9CAj1eebJfuxaEYzIfsnA8/gbT4Yq8d
IwLoW61eSuz0Kwe4y1hMjZmYi8C6iW1mAJn68GOAnsyor5JOQHpWykdC71GsZowB
79OgFefvhPIL7qP4LwDkFQxeAZiw5SSfWWXT5d9/IpY/Q0te0yBBSLN2SsT0s4QK
I/QG3v6f3hjLwQZcPRaOocdnpuhgjlKap16AWPxIqHSozksQZRG+JqHQxO5PToyL
7bT6RSh43Z92CDt6hvbMGXJ4LZErqEikgkfbQtpARR+lPoZ1dMNcN14DdeGRGiZV
Nuxjrj8UmlKpuUG4FaUzF0GXOdA27lwyKiIp2hD8iuu/leDtsy+tbnffiBN5bJ9V
ll86LuQ5ywSDQwy84closdRWnSv+9YwKqzdUyGjdi2LgTEPbdFbCspuVi67QscXb
h53LxMDVbWAD7tESGyXmofd6BaQcJSnqPq/YxAQn8Z4JdIVR+3QX+wtPjAvj/Yxe
E76LKU19Q7drjRWHGeP3HdZHV7O5DJRLUxlax3LWcFH8gl9kMN3ruoAXllaxs8V5
e5H+heM4mlCqfQz3YCm74oaUJD97G6DVaPLzI4GDpGDWh1Aih/E0iaLmwCupqlN/
19WXdWWvzYcEcBV4AJ4W4fp0Uw+gBabYuSo6lxUe7J2QBsJlBuodqiySqOnWz28x
T1p3cyikqZ2Je9mP8YftlzXxC1u+DHFd+7Nsp65iX9o1jf4lmCWmBBZYbteaiPWO
+EaSNQ1+cncfXxMYICdIvFaBf4fERv+nc2C71rlngvkrVXj1EJOb14sneUcjA4Xj
NHxP0AwcoWGaVUJmOa9zyFAlJYpJtxLNhEINedlWm836qm+2RLhQEUIM17/I1Rnf
lenZwczxJFbdTONX7iSF0pfWcWR8Scy5ETjgspJ7T8D1rlA6oCye9FhbsIM/VFkm
Ccv1OBqzzq7+nUlkq4+868HQEiI6XYbEVB/3lnnou9Civrzfd79xvfsERa4KP8qQ
8/SwRR6KpUnIqlAk08IkLOePItNlW76gBb+TydYwopeFQI2WIQU1LIXSdCsJu9Vm
t8D9OgSvxOHMpiTnMGntlEvDI7+JkezEjJ56tfSIAy3IPM8Q5//sqn3N5CP+EIzc
k7p//O6M77DrFcIjR6hEarxpIXVwobY8NfzQVtUgq/Veip3xiyAD/uv2DnJryJgn
o0SF7kibpcsCl+3aCRWb9TDf8KSa7Hdnoruqh5zvpjPztzBeifaOBiUxUdWlxtTz
kB2pU2lVFgNycguzKS2CYJRVrO+I3G7NO/7uNzKlEtXOMpodURmWotc7tV2MSygo
7q6cMYvaVPHhdVyUtNT2drrzKLRTwCtDDCN/ZoLI5XfGAE3oyVzw7A60HaghOsA6
KmyS2jmb1Agcos2efq/gBHFpJS3ZicoUNIoUtnt/9xsaRUDsCi8DJ84JSQgjQpv+
nXI0M6Od9pQU5/B9sA7oxojtiv5NmKQ8hhkoLAydMCjQloPAqNt5YbRp8+/yl8Jw
JLTE+jwCeKrQzAd/sv59SyVhFQ7HjKG7cxSGQRXKbu8=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xnq/FnahBY38hTFaR1VIgpiKM2HQb6oNe1xSimhwCcyaqhMWbIlsBPjySu8QQRTJ
n7ZqVj5CDaJ0EA6vrQGRh+6+lheFKK7H/Ri+o8dO4r+8Su4Iu9FYSYuzMnU6ni13
zrGqdpFVCrcu7Ig1oz+0PcbTvbKJw/c1WSEMZbdGTfmy4rG5AjhMXhkQ5bVwcPy1
ONOiDytEEtgaeMqQEeXA+DAvNZSdMv+q/JhKboP1BSc9JTT+iW1td9tZsdkma2f4
SQFoLABIos0e79xErpLOA34J3QkymDcILWO9iyhdC0Mxoim9FKispSMB7pfTaI25
hWGK5ZaMVpRhQFDu9TJ4igBt202pJ/TmEEYfuwm15C6jv8T6cbXuMjgoIpDNKin5
dR0/JcCnTYhRxIqFzPAjYBUXlHU1BQfyThwTmoFa8siHspg8XKZfySKXbzg6XbDo
8gC/i7pRy2oDXXnMdmYvTAttuzDpJnFJHoxuKjO/VsMeRy8QbUUn1XJ2SVTJVv5n
tknzNRdhZ9EB4Pdt91JYBaZ6Qmto/qhqlPMocnu/ysSsav75CUaZd6XIhioJnIiL
9RO76O9a6qRG2pNishB3JTXCeZZnMAKyGYumx9fJkqwewyTy0DX6yZp495oSfe4K
3ZezWidifNRrwWWK/9M6lPjW0MeEsxDwe+kxWwLkmXd9yXbWhdEwUyyI7kfg45nX
AUDMQZWSgm8c/ea8RrDWY6TACpqf+IT3w/37k1n3atxWoHhKaVpdtYwRSWMGIbmS
KRVDJluKiAFrfRZWPtfd5bfYs+6nb2JjrCoy3KATdZp9xW14KfIGao7Bk8Tz+2HA
PZ7h9gIJ31+D7uXaF82U3ORG1OEXLAVoGW3nJa3nfdfOHa3mn+FUzzzCwd19wNqb
Zc/PrHm8fokAYYX2JlUyphaIqal4Mr8oEqERghqBzBThSDnWiod4oy5CAda0IL2O
`protect END_PROTECTED

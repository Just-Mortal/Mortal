`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7oNHTNJFsLeT7RNrMPZjD2rYQec4juUn6MCrf6i6Gw5HLEdl3yNEN4bivFpxf8/
6+x5jLZJ9wTHKdjWprMchnz8ByiCd7MGJxjH0glsUzZk01cHWiUUdncBMwn8aosY
4zeqIQF71gusP2gG4tGmnkwK+cyqvlgks9N0RvT75ySvB60HXSslHnue592XLo1t
8aasR89sJ1BhzSm54zGQwXXxgXDat9Lk7z3CvuKUe3qUwCLDYJxtQ2vJMuZUXoY0
6lcFS3Q2jFtx9RS6RBxRnx8jICRafN3C7HkxpIAV1ATzFM9D21uGzKexKkB002M6
JcLqq8aEEB6mzI5+tEIwdmp0QCtFUzhiOTCwYzKT+TN35QpxONYKVoUiuCj4oJ6D
YZboKIM0B3jTatXailQgeCngS0fre9HUjjFZ82mjxzXPvT8mGxu2uAhMrb35aYDX
QyEhh7JrJosMnM3a/poN6yjlyEKAQLqnwRG5iIpUcGQ6MNijmqQdufSMW/Za2JxM
INOvQbGx8exXinjACRmcuz1nHmwfSyMXQ1hP3Cg5C/dKSDzku1AhxH1qVZdeOZ4m
/4q+OCV9OtUcLvL0OwmIa3LhbJBP40B1fXmuWTw9Eqat3j8wKKjk4noitcyjg99E
jXqylDmzd3F+CP7HFNBKmV7zGD+PWxR+eoPe0SqbuzOkC5l1LY6RjzWI9OtsV+gG
PZEcbg5DnPSq3qgz4W2se20SILLakAk0rmP02lBdUB4MBqIb/Kh5dNjlM/MYClEI
FKJZIBeFgJ4Je1irhOHRk6gk20zU2O+aLeEj5aEqa1sOS2P2mWH+KN3QhIDbqkXW
MjQP/R/RLq8WHUjTWfkfOnn3bMKkOymxvdO44nVRWqRHAEzEB2RJYSOFN/mmRgmh
231fEyv8rTf79MwYfAZPzrRdV6c6h6Au02hWiUoO9mfg3rRpBKn66A6ySDiGEP89
WfjNriUr1X+8MfaU3VROukOjlzUe1wVSncIbnuBRrEG/3cPcPl28Di5TBbDTUVcT
lCkvTNACIyNDj6GFXeCA6bRFvxmY1ESNhnd2fgLNugB+OyZ4IKlExqmqB6aSpTlI
IHjnJIhUs0q2c0oZO9k+hCxSFDCePyK+nCyHa+0rZ0zWZfbm1Qv2aRRqx3rviHbL
3QDft2hNtVx4bMkcaCVAOalMx7IR30OwvUNTebJk7EV8Fbk8HuBkt3GRG/W+DK5i
syTeTZJlx92Vo9mByXx1nkCYwQj5Tk8u1Oxk2NmFS0slTeoHhmg976ZqrMzpLfTl
bbrE+yvG+mi2m8g4gdRfKApj4qW66uhtiUx83uuX4F3u9sPUV3KpwSivuAzZxcd5
ri3oUnevuPjQJohrueALmXiDdhvCBo4OVVa6L4foo1FQmn7xOBaHXaZhm1O4PZh4
6xHBFvo9yDtuyGgmQf6dnOR0CEZ3cwbANrHyUY8SbxbhqN/f1mOqGz75nZntRUhk
sYJJ/SGUdmpbvKa3FSpbVvVYUWLXafq7RyLJ3qujEnn6hKInsSbGfCJW7qg96Svz
VZlgfDPYlu0raIEa/NWhwHQoD3UWIoVaslxqpI/+KJySXvcThablSLO8HZ+imRGj
Lrqp3uYws+8Lj3jP65WBtJ3KBuaxQ6teE2bUOA7Rta3ORZGSa9ufvTkhr/ddEipG
j7Q1hKuuBJJcY/CXtOS4j3ycGxsOx7NWrh0KYIm+COv5bqT7/d87cU+V70csdAp3
IFLDDE5q/WevdFVX+Bm2IpssBT1rNhPrKBSZWJPdxLyVMKoaUefNFsnDrFanKKIe
4uLue+dj4qmSNC7tn7g2uWPLHAm7BQ2OanfMjEuXp4nM1Vef9xXh1KZB6FQ9kopu
EB/CEqVh8JU5TXTNcDBuOzz5RmQ75p9JMyz8hs2hyCmELjTqnnIeUGWmAJgR4MdU
/faVkANGaitMWNXOSiNR5FngNSTamXqVEm4r/wPXeSt1nL8YCw++cF48rK9lgrdA
WkslWOjltMB1+dEjVP5vrNbCHThn4fBr8a73WgjtyhzXkXF+nKX7FCk6FZ96JlMc
eTDgARg3TU20m/QXBQf9XL+Ivj74VJ1yGpRfsMZ7e+RPQfv5J0bGJqQgCRDoxP+w
CryJXu6CmpTi8LFs2dF2HXPvlLbPJcGEnSfNibPeJMbs1KsSObQW9bp/xt3lUml5
cxn2iiuqBJsQ26xg5MzafMbzz0qQ/clUfgifGgqhhiAi9pxF6P8o74fCvpWSjl+A
fQqYtVbYFSjc+02xFcL8ez6xUkUsfRuuMuk/d05QyzDKwitmHLRPpjZ6hyv9kvLx
avm2g08s83dFhhxgWhV4mLvxYV/XMeqiChKDYfHcjKi9MHXEHXsMNcU2isICX8r+
SjfoS7iMH5WNJlhOLGZEW2S7XhIhlf3ZG9ELLeEFrL1AHjefSovCHwYX1NfD+f2y
bj4dFQlUS50VglkpOh4TOQWn6M4kNqq4jpbAQFbZxo6lcD/2gwQ5HK7jpr4MFUmg
t/fEuMBBMf3pDc7Rl5eTt/WzwJc44Ihbg71wAm8LBVyR1EEuaI8iDMKPKysn4YqQ
+YmVdZi8GcU/xLva8vuavGNUCCRc0m/oEaBpEg8+m9qjeYMQdKUqjyZatOw+5Gsi
PuGtzjdgz4xxu7nhtTwu0OPS7ahQ+EWDiynw2QxwXA8NZSkpG+Isybr29wUeK6yc
oj6Z3eNEjIbjJDefdidjcFOEcDN9M+WUTxFzyqGxF0kgEOT5OC1YG3oq1hm9NWMM
y0vj8t+dS04PQB1l48NOZEFzITU385qM+uMnM3PQl13EYyne9dIUCdDXDc5S0qtm
poDhvXFX3niAEfG9nuBW2vYniI3m0WiCyDucDosRjbwAV+n7ommg83Moh72UNinp
kOe4zc+sXsqbz1ZeCK9Ig0jxtyRtBDD2Wg0ygXVFdLEGc/q0aNTTVCDWsHWaFUfs
shyit4lDGUFs5X5oMkkeXIdZZSMn4bkvYKjMZBDURA9XW6+vJMNYHskdAeEQgjoZ
Hyoo5ylT+k62J0XGS33BVhnf8tw7r3TN4iJJXLRs3tg/al0i6727UrbSIHqHGo1t
d0C6MBZ8rLczcjut1TZs8n+Mc4cc/8oYTdvsGW4ijXh9SMILlOUfVCcinORUC4+L
urCBppwwzOr/T1eMbFIuPkVxlLuSC/zERNSB3BVCK/JjoqbMBSv3Q99pJJtD8haC
qIzpZDVrO9Dm9AK4QMR7B6evSKoRV2rSYa8J5L4hf8sVEQQHQRoY7LXEsnekKzLj
yyXoUn+pRqx2ZdxbgUPkFyftMAKNxVToblo1ckdB6oQs16YFwjczAoSkBE6LyBb5
P2LNHKMsT30ZoGpAtHTuu3gHL69hS4aLmXuUl67qHstKguyiKC1ICI1XexFmjV5/
VtmIgnI/1mnkBc/NJTz+Yq40ZM6aS3p77pFpQXv7lGW2D3gMk7dw77y2e9V4Uyiz
4EbA3FVF4EyKvyKRGt/enKy6JtVu6LwJc0JPsJjQo7E54CB1t/NnfORFZKk+FVEK
NccJeo9x+K/bBrwXRAFdWCFgYy7YIt0pukJWrZ9QnXIqH9lAjHijYH03C6KHdaeZ
HwatYyKpbIrd2ot2Q6WmieZb32hghuqzh114V7YiU63gpRb20gcqI3KZ6PIPqewq
MaQuRtP4kqrx8+d3en8C5BFITJo6BV7h3Slj6gsikdL1KFScnViLp/WOOzflDdXg
qwC7b+MpFxdTWqAevvWnfF5ucznIwte4f3KZw+qzbbO7NetBAh1aRp9apCoA5v39
WLu96uS9yGFp3tEOP7QUHKqAZ9dt2enqYK/73c/cChI8PojfpaT2xeho8F6aEp3m
WJLeWQ9kyVULuIiM/QElWZhvxC5U9o6QIZkHA+FxaMhSzYSc26jaxaAstHjFZbME
J7JPR9vmNuP9DmWOFLDCOpwrCyy0SPtXXLYssH1tZt/6WoAfZuRl73UjxzUunTYF
PnBJ8e2JQy6wAMCm745tO2Uppzh6cCSwzD7Zv6uT9aZW6EnpRV1xUov2caQLYaVa
hME1CqfehLynXaQSwCCg16QQkWtc7fwYTKqBLZDIDgBwBhG22jY1L1Ztsuj7LJWg
7IcczAcFJBJuTI7BWxk0xMXmXQNPtBueKu2YJ+5ucqTeDfM3xzEPcJ6k2S0gnsc3
6+FIZvbo9MVkidhHZ/ngKLYadAyV4kKp4KfWfWzmWBIjBG05I8BcKsJvsDfQInxM
x4PPrlY73BtkxPMbAY11NR4vHJe6ZpLbuxUMlosDf5aw2Co4S8rsDCHR2GZgetGL
B7DZZk4WXf3GeNoFtdCiHfN3aIF+VoSiLdqFvXyr5RtZYTVkpBrsgyKQv3EYBgRc
UD31+DBxT7sVbLoaT25hM2xHLA7ysMifAos1TxU515mMoKuypt4OCtAsPjRaqulJ
X9j+FPfsJZeqNWRn2zUnUun5nVaClIxLnUxJPeAztfOmOcX1DuIeLAMXWsF3a0v6
p//NGTEZnFNWK/4npnITIMUJBAWvqNa1Hpl/eEjXBQ7btxqH962uhQkGV0h/zzy5
f5wI42dBJh7aykWgikV8MtFiKGuoY5XB1O6u11xZUyUUe0hRdBs1HzLD3Vnu5Xad
MmNMtUQ0dtAMMEv/H7lP0wMLzTiMWMWtnjtx2sxO5Oepk15SypR7hqX3Qi7HrFQe
Xq0G2uguBdca3rSCuIBQNLqbI07Pis2+4LuDI+sQ+OCsL3wPEXKMKsIvwrtQ9SaW
RYknDE3wzZw6BASuyfKrYMFWAjAfN2e5+0nnek2/DeoAjxEp3GL/JcjzIxeCdejL
ea/yiBwPPXF6Ynb7uism0h5lsi5EEsAiMVuPt87U7QRo9vvxZPK3TInlQBk3A40R
0/9Qe4Z4XHwJXZctXDzXZ424GtBzy/1wRh+cd/yHuX9WLgsReViNBaQwjL/YDb/F
CX4gfgLneBnVJhTn2IzajOSzyziDpeFvmEDKGIe0KoZCihN2sdmkkK97W1uTJVvD
hmBfIVcCVjuWG30tx1xUCrsQz+3XXiRp42h7xxTC9G+yzvCT0Fy4ytBYIwmQOPr+
uL/UeZ0Un7UsLixyIZiBqA9oZkF0P2OTIlmlwHO1DsaNdyuukviiFyXZLVnVQTrE
5RwtmmP+uEdBMmuYZLrbHv0CfnpLVkbejz4uAD7P1dEyCbyOBYtA8TQqrTskdh2z
I7CMe3/Sy+LGCl6gLlG0tey3OAcEjwYUnxMn9SyotYFvDwsOA4+TDKc4Nz+sjKDS
QKmTOjnTAqK2GVX2+XhWaZWI9ZadVQkTV9bBkfSZH8IJT8jyHsP6OJqPXoytavc5
VrqLJwG/iAdzN9N4z3eXT0ls4CdiD0DppjGA6nXeRNg9h6T9nohpIXkHrw9m4lgS
7zbQz1x19PCHt9yKgQA6rdq45cenzH/ztTYz8uLTfSpCemsIii9gY3blR5Ug57bW
l3xAskbu6zKcI5iFvol43tivVejsYhpTqSV7dIDgKeS4EPBG2UidZ/QJ2XFfv3pH
0E97sR96udPShElfi6KXaegb1g8IDfu1l8dIGlT9RyCpMnOMcEqGN7azOhkA4v3o
qWLisxD3Usl7IwuqyUre8HhFVGwHeKsXJ1aSEiEJZmhvbggDZrZ6+84bWlyjFTV/
3XiVuBTRuYF5MPMHit0fyPEm8CJY7BkUh44Ab7970E5Ct7A6GxMaP7KD2rDXMI3s
8/xam2RKo7vVNQ3egB1NHuxa8pNm5+1eNPITDnW8ll76qDRmPNQ2DHWccnnl5lm8
coVrPXtWfjgagdC3QJlCzbHzTF1Mq85UJtoX4pN8g7iEuqGsqNiwsLGnyrXmuztw
tzSAxRNNTGNEEc258W4g9lfarh6Ae0WsE/QcUU7cHGL2u4kaTRjKJpomPFSzF3SB
T6XML9mgZzUkb5BuirKTQ9lifARBs1lgPSFUvhol0+WO7a02W4PYvqCmA3Pf+Vt/
KBjugUhnr/OJjEwSUWeNq4sigxjcw/SX4vL64ZFO4ULB7D0g0guu1RWy53hYlJbe
gf9I5xod9lP5yeTV1doQKmu5ZOW5u468EUy5PUWIUb6kwygKmtvv+yOSM9ZCATsJ
c83DMaah+1xtq3IY2tGFqOixgRFJALC+ZlBpupZVROqNwR5bluqULV0hvQ2z6qfq
Q60V5x87uVyu/as5fSk8ZxDRrrUcu7SD5hDYXGpfciC+CidYQDlOG3w1Cz7v7fmn
XdysuobgCHPBK3JG85IOWG+8BKQ5ahW+Hu3wIqHv1uXBx82xngDlHJHy5NGvOeEs
mB6V8GcdMneqzIktllKAHQh8BPwk2sSK2D0jgs1PwyAued8h+N1OcY8jPWfZVaB0
JXQGRtR73kkW4PpC29fR2eS0f4E0lGrgZV6RBS9v0kA50A6ghUD02CY9sOTibAzd
NAJFeRYF55RIrBgPi7jStv2GU7LJEZPZwFAGyNXbQ34IaZdFdxSScsxV+oLYGOqS
QlnSewCfEXsuFA7ZBPl1uMhmO77SHLAx0+WW0Zh6DPepsQSJTw7Rmcp95YPnt4Xt
9zhMSZcCQ1Iz+4DFxiPqDL3sCAFlM64telDcE6pucPQN/qoW48GtMmw2MWsSOxNe
Qzu8ZwEg9j6OI7+Geqh+oTr0K3A1VC/YKlhd/ne+Rl3FByFh+WSjhjO2AGQcKA99
j+tMHC1PqjR11mlzy8Jzfywv3HQeQqjaLBhA2MtjNh1V803ez2/yO89kL6tbIhmz
fKJQmj9HfU+2q5nQbDdxrLohLL/4xqO/9QtM2Mcs6fxPUGNVgFFbbqh0Dv4b/nut
skf3yCRKrYiqPFFEULx4PSKDTr88AJe0FQ9JvxyblB1xP/yxMzgLPZF59W4yXW6+
A6G6vHsCFkYgS+vCjQLHH5Cm3ubKUeLiewzVUwD42UIgl5TEyGLPPUtpsIzLPXqF
99c6L9ls54vti3EBfxhw3nvgZZ61PIKqKxnPrtY8YHsMkg8J3Xi8FzReuR5bn2Uk
mpeBt6xRRg1QTcy+/Mjh5sE8O/nOMsvGF3m5UxbJfH7rxpJS5zZlqrGNpxzPCFQL
ckQj8q69P8Gm2urSbgJa/bKdLR9a9OqGH9IimTKoM6v1lVMOU/tYYVjUuXPrLaiM
/TT0jFrVdWCfaE4/JEzFhKL2t0wj68mzUEx6otW58dY4R0IwAl/+fyn7B1iWmPwJ
iIbfF1wcVHLCT37CSdUUMk+OqBtWJPgzoq4sQYqAi1PS9aqpw+uuZ5qFucq73FNc
ntU3ovGH/RC+pYSTgNgMEmXiUSej0Cyz9w9fCasu/kPNDsH/XNW6hnf9kGn8246m
0NQoGf/0NEpryoVnaMTmeXQyGoFk0b9iLwA2eXXoIx7qFo5ljKi6fxqHZn4XtOtm
A07Fw+PNi3Td6lYTf8/HhkowiXkxnzZHljjjVFtbEk8PfSbUbOeGQgIRjoWkZjnV
+GGea4xHrklUat6EbNyOxFiF74EPyYLTKI1slmOrTm5WuGexXxm9gaBQOZ9bkpq/
z9BnXZtmYRAsKd0vMOqlWUPzxn7opF6HWY9PhjMZZ9g1uNV6X2eN6MejTafkSiA2
QJ6KSwXg830631zrHt5Bw3oSVZR5ycT79H0Jpf58ARLZ8pEGwsVB/+IOF63w7ZYG
fJ5XjsUULgyWSe8LhstpEWQyaKv7IWFE/yf0z3oseAnWlyGk9A7fQuAh8KOb8UJ6
V5GO475iUZTvjiI++pSRQmfrt+wTmnhMwu0jhwe8btIBTA2jHqMB4Q0/zSARqpc8
06ep/6chhkilWyuTf9wEUsXhOu6GH6lE/yWgWV5L1DycrKgh1No24r8LzBn0tKbe
ZUhQd2luJSQuIf4l6Ya/K3h2GRJxkQPsaviYOx9GoXma3vTHAOlbNuP7GzfRvsWJ
e40oWzVx3YKCvZ1ciR8BIO+nz9ZYMhVh6Enp8beGGMaaQJ9dMtrFhTUN8bhQLsbM
hqQ76RWURYig6YctSP+6E4YeEu0k9SLr7u2D92exsVRu6c2NqR6utIpPHHDBlVKw
glnCw8hAz2UQT+j8T+rHOc8wW+UMPw5XeHBEsvKnICI3I/hUme6ynKSyLtBT5IDw
UzVYpgiDou00lA1XGZdRMHYPiF0gfak8tDtaW6wdmbr1k0mV8w3GIxdn/VRdS3ge
lW6VF++XkeoBSiw6wiLYSm6X7wH/A80PXk9OgpgOEJKU0w9l/a42WoWEq8IKnoRl
2TLdOjTO1c3j2SA4KxcmV4kM55mZ01qrVy5VcrNymGyRaBnHdjj178Is5pRJZHqu
CJgO5XIUPv6ETUVbOcKRRAsrhDe1VJO8tvePhO2lYg+Hh+tgs6q9cVTjVziFYFIl
1mI3Wp1Ss6ZtZEkC5Kj/XUeLKXIqQwLDA9JAioc5rKXBEDjhCNJFYuGnAYu/yH0p
3mfmBH613+rkJhoeSSdRO6eHdW1BFUyHrQPvdFRLZ5RZMB+/BEem07NIV4DzlDXz
6FgHSYrPqeUt690cziMPlV4L7+orJHTTOkFXqS+UPI3yeCveSowHsuy6a8K8pfsC
DFc8d8dzz0AgYmj1RE+umeDSwsEEcMEqBw1DcOLEj0GMBoXUENAYZX5/3zSlbsFK
ithQet1CnMd19TJ0QkCAR7I88//bPluv6gjkfM9nxSp0PaaBlS/A7ElU98UZ+VCR
IDdGDp3NKoI7EU+ByqgCetGvdkrd1Mw1rOjiPnreGNdzx56VgPYeQvlWA+6k/yHX
k0j+csoLW6/r2XvkH37gXlbQDXkMEuBC9p0qYp56qy2Wlq0OMR05VzWmfZf6JelC
q2cf+5gLqAKtpn3lkY6U442X7/fSK5c6sV+c6bXGSl663XSDoijQ7WgtBA8RzfNK
S49+FepQr/qX0QwUa3fbmP8sIxaN6W4Lnrv+1N6IMfJNPTHhvRqcpl3S95VT3ORs
V1FhFIZKV8fJ15Vs3QHsHt4CH7InNcXlNx5Z//A9vzLHlqM+RVFAaTRum3arn2nq
m2JEHmshpo9b6OkrH+Ej10/zsT23GqXKhFE3CUZCLcTU3A2/NAKgeDTEjqRTJwVw
6rUcMgf2N/1tg/VI+7lMT7YybGrPHEhtmJ/1YyXKF50KNzjUzXUcTMirr5yM7GmO
UV4sHDxjxIlkbi6yTUpjDouFGt7KsEWqMQnMXSYAO6NWUKKfFARytDE6JiR+YkYo
bbv7AEV+bKqEuG0aibWrUEYs0A1YEf3EUAWoO+YwpX1N7QwTEom1IKrkUmCcOn9R
GCU10gczevvM7ZKn5H1lJS3HILI4ccBDs6obn9YEkOi9ulwQgUobXWfWXpCV+s7Y
Xu9gjanuyMSQYNZgflFZeWTYFanN3jWf/pEQkdX/ogmqKNuIqLRls2N2o6tDkSaP
LQqpWVW0X0apUAAxWI5OtFHNy8e9im9jdH+7lImFL+4KFy25oqe6kv/r/JW8A3u9
tjef2+/TCw4g13n7g/mX5r38UpDNj7jK302B+jSFEUfzETMN2TGAzn+gAQSjx1Tu
T1OjiAP1x3cqb7kmuNrzyMcf0FkO41BXRpHL8gEl65GIb/KhsL5mG8BWa9DZQxk8
OQPNvHH3aJ+p7FZYgg/gge2NTvZm78bWm/FWqk2Jhh68FfH1kjUOT4wo0kFWP4RK
4O4rS4n1AIdSzo6vm0L06xfJfGbmp4gd/kMhEGZIIfElEwaD8KeUBrakWngPhdXK
d+88PlM0toDiyM/eCkKjjR5/EJNXtdhtaIrjAPuV03EE7L5BfmSQnlL/CLPR0WSv
HMkSDfEheiU2ujb9bFpuiRGI62aBL/OGj8dbuwrBFRAUulRKRr7iycjmpoQnoJlH
cieuJsBjaDs7+b4lLIr31KZh8ezkC6NDAgeP6KUStG3baBgcG/L9QkrlElEWDFIE
80vufdrCn3zeyJTy7e5s74XWKSD5Q6X/FL5y1oAiYETAkhk9pJiZx3igm5Jlqd33
sM+xQFzggLHTR5+PU5mT+Gl0Fg+mf7Nx5Bx7umqFovvvhxEPRShsrJMIdnOgaNR3
6+HFJntcIeLYbHyahy7Osk8ddKqBJYouiOCCp/3E1FjhDhBYp+31zYSfB3hvP40C
5uXu9I7Li4aBin94juqsEXehnBqRT8360IlfU8B3xZpo6CR3MQenUzvG/ZUDBM3k
woITXTYUKGMZPH+Re/stqymh9ZPZHpz9Pa4gogL8v/C1T4DoaI7x9CLe0rXaGA6K
2aMYETKqdPbC6ncz0ItjLhokjECx1UL+phcnwyX6nZLixQRyvNiY43pnmBTWhKQo
vfU4gla5YNs/NXHfNHlf8uffAffMfCIMa6NgevOa9oVyCZKpf560Ho/aVCHLPoxE
6GSabxM6yhRK64QxBT6HjkI7eQ6FkAAZEHZ12+HnC6Uaqy5R7RVv0MJaN5mVU6MO
malX7rW+sa3lWQxTstbXTL31fk4i9n8kyHuW1Sll8wJNBPDmLjCaDqIKxOGQKbbt
yRjkFGV8ZKP7aKV5rp7pA2Ogoev+tTQWo8gQPbCI4cZ7aKlG4wbIJPOeASLx08ok
QZnoVF8y6xB1ugACw6a4Mio9Pf72WY9qXcZ1tKP8yygca7QGYuazTSQAKASvU+Tg
yI/cmJL6HG1TjEYoDAOx8RRFPWvWR0Q9eYKuX3emHuUNn/j6AiSq+l/MM4/8VzLK
Zmb+58pvtVzySaz1aRY8pF34OMo9nioVFDZCW8jnM71xUXv6EBGApphkcd9b+wAG
HHdLUKKVP3uLu8koZTh5yER+hutiiRucBahRypmK9a86A4ie4UWsM3ila2hZkFT9
NxUyP4WcgqkAOgVOHp/76lJXaJpGRem6PFyeYEMpjpBfXNq5N62lBg/qh+7B2B67
5fUs0xfkXSN+et3Fj6aK1gtID3ktOAaLekuy/8ynGZtt9p79boQSMf+vSqKaXOGX
HmABS/X5o48D3E79MifLG+MdnPn2Le0NBFTv8gQOA86wxwxCq/NiCqLoa1O84PoK
nUGSTpJ0NruY8VQ69rJQZ+EEVuBXXHu48amm33i4kk0YQ8TtW9lL2oa9huQbt//J
GBz8B9iTPyln3/2iEIul4JYEjZfBdPAnP1yHxZC4fO5piMys9BwHibtF/3CSkqls
LBj7xYmgPpusxbjXjEhmMmWRjbwdubl62Mw+TxzStZEOiSE5mLCerQR1fXMPmbvg
AhMDBwJONZOWjqOYLDsrGzt2jjgYOqPyBUa3mA1TmQ1Bc7NcEIkDKyinsP31CHSM
vRlf4fw+IYcGuiZSl39t1UrBM50w9C8zOHmy3qIlNYCNlCL8NOWuJ1gOjYTG0c9K
OFpM9oAl+S+MXXrNbaCaclbZDkMzceXUYpBTo3IhrET2kd6BETAn9K+Mu7x6WI2R
/ejGaBFySRTdC9k1GwZ4pTySUh5xoMKRrEcA1tbjASCVyj1TxZk9qRAN7ZHm96FA
4uhFBWP1XFiFZFdQxDE7g5xks95kqU/67JVi+Q2IMZSdnJI2P5c5VByqz7tElGca
/wdNGvxS4D8jyUpFPnRrd1OYNkgscImBczVR5otbUxPS0ckAQ67MmZ+rZsx8ervT
Brgnc/KECANcGxfO/L/mQ45tJmmABk1lR3aT6BAEJQvkq/wOabwbgvJD1X8uuxG5
82O0RVCyXDITHqUL7d3SHQwMVtqy7y+2OVAvU5Un896ysRYx68Erg7E2Eit1bRpD
WcpM/Vd0uT+DgvlYFlKulYr11jVs7MPQl0Cf4UmeI6TZ8E4ITmGGKKyaZM+9OAAV
ioq0l5IVcYMcHvNZXYEWZDMlIfiZvHG7pJ8eBvVoVNVYbLNS9OQFFlxdSwjRVzBn
dxhGVIM9QjvM9E932I+OfowT5n05AgrSrXmvccESJeQM+Yam46z7NqGj0wc1kicj
sn9AAJv1/pmx73XYM9lEBD8OnQQIYxz1hG7fclZvavtxKxPldDg1T79RHM061wZ/
Jmb7Z7U5I2RukLHimpUdrFC7HObxC6FIjVdZ8fJq6/G1n8RISqzGVP8pJGEaJYRD
be7S2aXghibpb3uVQoMQkKKNLysU1zGhy41lpJT/XFE4LwkpRaPcIw97xxrY/UPe
xbDwhCUgevuStKgJwkLiSwxbPD7+tN1seWEyI5IBhlghkhhSSbsp63He75pLacNy
G4p0imip7s7H8UR7aVE6XCv80oYqi7KXFAgeYnZlxWNf+9EKd5foHED3sRh2XTBH
Q7eDwriFDjxtYC3bm2ExGaJtcTCDgqxlYShkV2AAtvLtjEyLOx82kww7RgqqO6cq
YQBS1SLXIKqyWT+E8TOGOyxLMhuq6cU9h/snhLHeRFjdY0MfGVMxJCrnxjwdkwx+
TMf8PzO5WIShvsZdiVycqP/LvKNiR02lrzA7/MInO3a5FFnePaPAi5AVmXgVOVi9
XsN7UISawFkDfF/yfE1C0F2qM51Sn8x0PZv3qmRTh0KopWcRFUU3SZMxICBwugfh
EmU5GxXeTfdw2AYCl5SB8Bftdl70yFK87ijtrrjH5JNZ9UUuUb054w7vKtKUWgri
PQBUczOU655QaFiIKAUiXA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qe9fjCRev7NXAvsKu5ERRMzhwkpXUawQMum0GHK7mOgIBzDCWmTgbw5k9iYX01gr
DvaK1Jt3QRyK3cfitym5tWNFjEl+dGVsYpW6KWK2mLE/XoPoLgVIRlUmIaibtMFg
wpAhZHBSfKU2twpjswTGbfAUwwVLtFn1VABAQY3vyGVXKzp9J5MP581ZjNoxXpQ7
alfo4XV6H6lIHOL6lqNEATAn7eq7i4RbUxJDZpf5u5DPbtclN0hwAIcydnh4Ffr3
2WOnSKmRkCD6bR1EMJ7fOHILXzaSyZ4VpLkO4Jf+SghpEzykyTozH3dgrSO+TKzd
Bjq/73ujYYG4XnRzZm6ai33c0OlSvfoosJdef2H8LEIbSPi+S4OwbjisrW7UvrWX
mBJQa8G5Hd/AE3YgDy01v+ruoQh2nP9VRZRm20BZlPQWEISPCTW1CIb3NKpGuCyu
fsc9l9KmgZ1xeZkETfoa1qeorjCaZdRqbJ0j6wufQDwMeNdNiq7X0SjwXG8wBeaq
dW6xhu+7mHnmaj2kMxw4QuRktGXJ6biGlSRd9X5wx3AqQ7MYaKe9n/QPdk4B1dei
W8dkuopKl3MeqXJ9iyqYH9HukDtYDok+svpy7ztTfooZdWfExQr1xkXWt2GSxS48
CWRrKJ7Ot+v5GJZtKzBhLwx73PIdWJTvt+wmDGiQ2jVn2dGF7d5b4vMTn+rfuYRR
oErSm+jIxioy9vSH+N0xwcIAyzOBamUarQZVHq7cpjq7vYCJDQx45jKeQ3L/15Eg
TvqVlFB2PaDuKhV7FOxzv68z7j/JLAPrhIX46BN7Oll+K+pt7nl5uyuYCOgRG9oz
2SP//viq8RCmOSZs6jfI5HmG78L3GjBzft2rPvHJYR9BL7m/YJC6T752u03sWdwc
NlGDQrTp+cNhSRTka6nFdyR6u/T5sTsZ8qw7m9gBwEeOOWzUo/mg4lp16d56EtMm
0G7oj4GAHyRry5o+ONgGD4hIx0oSQgaJwrWe17eFVVCYsWy9o4E+1ukzQW6oTKl9
ed8yTyKhbOWXK42GwFpjtKyNCEGpnettVT8f1wktxuDoSKlTgW8ng5Xh9WyGqfr4
9Nln5X6F8Aiy6R56qqN45+7kX3vXzymMhOEtDv3wlrKWtahGMbbGEwVfBoQfT9tL
a2JgLeByEV5umEL7A1z+Kh8RG8yt9vbp9JvBdEJUg46W7azjvhfDGt7H/DMTADNE
rE/7RevOuJa82RCeVQnzmcZQlnSMUM1R1WfigbXYTjk7e4n0q/hCs9rHxymk4s/Z
EOK4Y8sU9qnAosv+MccY7xZ2C5CRXu6lesD8r9aTE2MspZGukLh+Zd9Kx9DPoggX
AsoBMo8aWYtRwTm15ako7OD+na7gp4BW36CZARU5BUVDW9eV14z7zJNPPuoULofJ
XTHaY0SqWg9TWzlSCFsJw8BQr/5ssEbIspRMtC4qTjE7tV/CmakHWx4oZuNTcT5t
Ir1UUA1PDtv8yRKo/Qpv4JoAN69JvVnx6d4Z5U4wcMhL9AOPQa6HEoZLO5yG0BhE
6DzOyxGvKwRw3nSWEgTDrGjj6LE65iRJKKEaA5q8aIligKVkzscMRMV4mzofEKtD
RBscB/tqYPdUm14MBbcIEk2fP9EqOlQ8nmdJen6iGUkZj1JMwMwMncNzLhre2Ypg
1Qv04OYoPUIFrwM03TQHXtEd9+lRGmRdrCLqU1yAYqd1ot7ymuIO09UAXwC1QGw4
EscmPEGIZyV1PuwvFBC1OZ8ZEl8GaJz1TWjL8AS2gyuG9wkkA6TiHIazq/z2iltK
fNpfYknsrWQyECHZTsxJMLSfGgXOnmKVBeObG6EkzJSGcyyO048u8tP0rqaAHZon
Wk9IWKkipHLHTzlAVUp6ZRfrdsn2GgLQhNWT7sCnVKnVjw/ZyNoHNyQedVvGNhB2
yoVUn8xfI66YcRb1DVfnRne/pcugUEhuSBLJ8c5mPhpKVbokL6i+2y/mrxhnTOJP
bJ3kbQoTcBx5ZIUbomv4OMhaSEmsp+xEWDNA7W4wvgy6H3DLDTEZq2wlmhIWUV86
gXEr5yN4PjqUWi3k/DXdmNxuYcW3XvgnufHbkd8SRvFSAUAY9qDiMDTsGdmzmqnN
PUc657a2629M++pW5cNMTAfyEqXBP+N5V9SBoaydBE6CWU5cABfWU3rNE+YlGFZl
6UG1NES30B8bL+h3X83GGmMg3JI4WcVt61/rUGcUhVpC1gkiHhIqXp/rDfx+fOW4
eOe0Xb6+xmvBprcNa8ZtZZfXYlUxvSusdv/LRZUwoDq1Z2Cr2qDuf7s9VP0fCWWm
immHaCYcTBlGdB3lENqR7t0bI5YYgTpsj0FF1vEdHYftpAIDko3TgAbIHi8vtzie
jY3rUIdgstAfOYQKDl+d6cRipNQ9SC7Qu/iZ5ZJeEB1hjwFG2BxEi8hjWiHXWpmY
oMEChiejiXplLnzA44Zv4Qb/Gnwxl1gkFrWaEM7lxp88rxlTpB5LDdBj/bm02SUf
6gqM0D94JBdwewE/mI0GEwchjp2lnEvL6tHbTH7dB60zFqYi/U5X74bZYtc8vVdd
yZZjcSE9hFwmPvIMij/jRXe/gNx/AmuDbS0uS1gqECge2f37sUhCv50T1De3OvGf
ztn4OsheOK0a0v5y3t5L8J0GyKwGqh4HNf8MoNrLd4uRmykVmb7vk8Db6WS+O4s4
/ccQAIudlPzafkfoUxIToxYkzyiDDeoLnvLB6vXYNETb+wbU4lBGG1gZrH0YBD4o
L+7xp4U1T5mOQ8fwdhnMu0SQCpqw5RkFNKuTugMI4XiWLuztKeq75v7zutFwYeZL
+L0HQx+JKVJ2Pzo990rhKoZSeUqMcFKQpk85nai1c4K0i+WgvuyQgSvJVufa95y4
pOaKF+MJEVFmXpvMbcCHaFFDSQreHn7LBJ/WcRQo7Ks4ka4IXhURgpkzmXIpu8J0
8Acz3yyGVufFvVvfud/GKtBzUCDRx3mPZmNOBZSImEIs7KaxrHJTuPZIgD552rpb
bQUlBKqdH/m1rKY6z/nOlPVm0eOZrzlQb3VVTANamu5+mV4/bxdnoZAKX9Q+QmOk
HrHOZ8v9Vjv/pIW9UR87Xwc2AUoaX7KzmXvl42V0xoFG6U3eoaoNM75qJ7fcf0Xv
YRoWSDD2k7EpmyS7nST25eLd0IMPJFd+o/3Jsuw0H3Smm+ghQ/1yDbHbXgwLf3P6
BK5hynUUhR7Qs0rp5JLTCtVrW8Vdw2ITast8gE82dCZzOnOmxl7jgSJecg1SLjPn
5RN4Sjc+fs0VbkND6wYr1IzlZEVANBJ+kyCdDucy5JRv9fo9KmYEBg35362IixAs
stgmWbyFB+dyYo9u5j+3CXPnusL5n7pUlnE/TVMMPIRrudh4UUOau6V7PxqanZ7z
sX48s1dc/m1GKS8NikazrC7b8NhyBiorwqIHwO7hn37jTKMhLTj9pNWH1+22UlE3
xqAkowSVmwd4oEvcyu69stXEHbEJw7IvegjgNkiYbuBnWZADI33WEUTXpOEc2ZRD
01B6WHSyHyZLYktIAcKAWW570Dgikp0GuAgI+u1FYKDaN9rIbq67BnJ3AvDmU82n
wIl9EXjSOZ3BWby3wLMzA8yxFa0H/Ro0iXoBi/5OqlyeewIzFnGvIY3yo3BcOY+B
YHCtujzugpYvxiVPsh5V7grvCA8tMaWdsxSDrw4021DpzCqXwPcTCkJuxUg53VRn
FgQwoY3O86MbmMddnHAafXaLJqkYBzvFHBpKLi5FPkcWBlsHKyb13fIdika2g5Hf
QtBD04C4f+Zhfiq3//B3TnPuoHw5ZijOWzV2dpvH4YP1oFe9hJtxwWT+pOUONGge
SVaWGGEhwSfbckt3GYETLQoAZUhB5Ad+TTpWA9GCW/ApRddkGEmh0ee5KAMCG3rq
8ZJ0GeVbfb9Me1tuGrAQtpHZfIxOmaEWsYUStGWO8ex3oRS1na5wl4AysraUo47m
Y1V1+PPmFucd9LicmONTO7dCBh6pIfQMTljWNkjr+goS8iCQJyPjrV5c0Zv9ZT9C
1z0EToD9G7o+CjCYhhn4s7Vm0y4ySW1jnzbskAfMyu6LDfwiOdUocHhImNrq42dQ
kgAlXDDOJzGx5d7P16dgGk186DnVbvIj3+wUyqRTKVzDN1VpPB0pagwiyl5McmR+
+eSybvIlKLMGf4GrBkjT93nGpGROBIMklHmdOtpMappQLOn8HIEI149nx8PjgBK0
huSlqir/peCZXYJgE86cfCYb6kNzBTWFfz0gyoyAOjXq5tH5apVXKVLBjxHypIua
mzPT/1BkkyCynGtx+bTRVKt3nWiI/fNbKpzdZpEUyVZJCtXfySLcH8WmZhYbVv9G
morlOUkhx74L3/Mkq58qAZZsCBulUXIwmEbQUliyGGtagm4K3nhgmCRQNZd0n/K5
hNNaDNyXkQQVQbeXNcDtZA6V+laNrNKIgNjk71iNug75dcbvvGyY8bwcr0TSFEkm
18TWSRNJpKpb+YClVJseJplTskvSJ1xZhKru8NIdwWDInsyXH3Ppbvgee0tHHX3d
QWU0ECfdCgCtc5gg8g+/B5dqHEbhAZP7Uj67KYupvsHgg0qx9HZ4GUOQ/kk86EmL
I1Yk5dBsVTKPlUmt53vvDP9Ru/6aLGDoXZx+omo5mObpr6cOxxXAu8qsxOe8aNbY
OZJ4c8BRYPdL92LIf+Zbw7UsTu08D3l/JKyzi//BFiEJZxLLi0GWaL1LA93a3J2p
OtCfHnzB598g2sDhtNGTlnczS3oY1S6/2ijFXmLSRwzsCPkQqGtO7ANM+2xR6Ox9
9+M9YGJh7Fv91jsaCjuxFCdcOym6UgWeow7IF111FsghHh8GifSRTDCshiJ/Tp6b
KaqCvgBWR2No4UW6rDj5zSg/wZVXFc/k+uUDcBytzjz31gRS+MrIimkz+nUQdNdE
aw/9UeWkHivUKpYjmq6IeyCLnRhkhV2H7d0Muz6pT7042CtPfrBywqQ9Y36VG3Yk
KuDZzO92CbxmBpcrUGqjqlQnNFvghwkbZ4zdlV2wI556N5xwB+ZFyRb8qcBKYAm8
BLLV7SwdztYrUEWp7JhzWYsj7eU/zVqhPKZnkq8S/C0jxR+jUM4+Urzn7o+1LFQZ
qfKdmGQwAv+TM006nY5o5rMl3pZSKH1iqr6DiHNj49CuLVa6TgjXlCYpeUL2Pqqo
mJD+1K4gfKieKszlwKOgBG5H2IwlQ93D/2G02p6wa8u0mO3u2/X5fSjF6Wli9cIj
7n+T6EjeZB+dkqYA91h6SO6ttGrnhyGIvv+DiMlRJwKnuOwiRT2X06zj3pUBXtq5
p4Iy7/yXCdhS5p0ZboGt2YPzTDxYX9W+FzVO788ngaI/dJVDgxaz1qq+wFi5z5in
Ip/8kH8n04rtMjO39yHSfmYu9AcsTCl1auFoSJgSF57XCdyeFLVPnFhTjhcbgOut
HIKYTbXZx8lV/XP0fZp5IAG+Yf57NCTfk0XUzvWs0VFwcG2+14GPH/4m7seq+jY+
or1luuUwTauknEeAEfBqT99iMLF0oPDutpZCay/5WzMacg17k0u//i4szKf7SHCX
JUz3srwyKsS3EO3u/fV9KApH/DRNvsnMhDgWSvJh3tA3RmFvkYRAGj1p0sXmFbGk
lE9MqPjs0R/zTdpcKVFe5zoTcAH5ZxurD85iQ5pKCX1hDRIyPcLmkV6TDhpxGTZ6
f5zI4YQLgzn920gU0mwofVPhZAf6kd0GXrjfAQACW//2NUXHjZ4udJlyjXgoW+XR
AaX91Vfw9mYPcZbip8lRq7Y3cBfEO476MUVd1rhxF0SmF0tjZZ+kpbRzimNCGV51
4tZCp8iH15wjdjkY11G109M8wPV/BEXnAOc2xS9MD+F7L2hFS6redXLg0d3EJofp
LNOfIf+VTjOKSmxV/RJsadiEALotnvdJo3B01rldvDbwfJxNPLKEf4+HV1xXd+w8
D1vByWnaqFfI3yWHGCbiNfBJ8tFb6veOlG+PYX0A9034wZUz/yEFQVLHG8LhKb8k
/WESBHkX1JdGqXhpc9w+c+A7ZP379lCBLdD66P00bzWsPHLykNPOwvfk3ZX7aZbz
45D6COvUGF6k7ZIUYncGO8ObfCoQyrTSr2tPtc6HD3hFAwNwWY1k4SAO/vkIINzr
lomU5Y74jItnFyNe1UiqJRRbE4NTdXTZnamvV0jJxO8e6i9Wqc/JgjbpvX2c8pb5
WhbPZeyxsAIkLTjBbcaCPR5zabQ6C6IHH04gfWsFlp7ned61YsbZCO1DjgE/D8WZ
9ELmmzA3Jmh0HOejJ5Pf+dYxX1RfvH5sXuMPSlCawUdE1Srfc3p5i8yrGT8yrM0W
yloppuCK4ARGACMmdJdEth6V6a42Sb+m3aC0ElHXuhv8/GV95oCRMm9RJnzy0nRa
5CPc33kbjo6dcKgTk7Vo4N7BhsQKx5w/9PIDiQXqgw0JiX4I2l3wh5g4MjZSZCzO
oKYjNap15S4dEnQ7vV/ZXJFAhdqPS1dHAKjosRkUGI6lgCOnnlNY/53nbZKS2teQ
iKTRX5jEWbHMNCxScPqBGQckdRqw54dtN7f18XmYqOAInX1VpR43zA8rGR2Hb6bD
xfG6ys0Zv2s2AVkXxiMyTSnDlc4DnwhqhK4lynKifAlAwo0IU+9Qu+7oRWgFmXJx
W0kTNCR0xm45azwgesfrE0NR1VhQ2F7/ggx8CtRGHyUWVLeO7P6J9ozyqyPoZWfo
kU3A+6zrkGMB/qEve/LAN4WvASphRVQ1bb6droevy5ocesZl5UQgmqcFAQShqm6/
WjBXYW4EIhSoWOho4nlZ2VMlNaILcCBYTpC6ukeID2xITC6ixXGUb2wuNS/ycIkW
4VHTNkxDkWCohBvIwPaXmmr3U/V8j3MoXdOlsHXZ/q42dRNk9JdC2OzEHQoEfT2P
yx+Bxh4GjCMwo+N4b8doy5mEfAzUVxR1iaqtwYrQ8igA2/3FGN4C1yaWGY6QnjoM
1Grc9lLJT34UR2mk4IHdbZo9shrLfyoUODq05osgjw8cF6X/FEW4EYkByHy80caL
0YY6mXCmbgafibMkhD93t04Eb49nPtWpr9FGxKkpYH9Ui9J2qFBcTs5A90I8nhJU
IQ5zqO4Fg5QzhnMr0p9JCljSVw3z1mvXvkMRZRuhut1isVj1w/cT+zDCrbHwhkv1
KTmkG1rb7ZlSQqesoh7XN8F58GQANM+C6nLS87S8OwHdu6RN920lpJO8fiMaNjqt
TvPmGVEeHib/WfmUcXZ/x+McOnXY69XOqPSjpAV2azm7MsjYKbSXOx9DQ4LDLjrL
FAHtBc+WvIqz+1k95QXbJrUttaH3bw6iwSnaXcFiMg3f3UqZG94Vw3lGOvEnZQw8
TW30nM/nszYVkwAV3ktoWQ38tvxSbiyBssUIDfxvzo/n8taPGe3Rcv2tP/Z77RTb
YrDXMOG8AhZVAr0cyG5MZnyGYWmxbWh7NHU3jPhqqrMz88H3H/Hz6RL466a356Gq
lJ8tEdeIlw1J1ayzLdK/4k6POaAfQNrjgyvGU5CvHSEicV7jN3sMC0yyc+ufEynd
8/bmdNixUXZSKSEvU/9kkBC2JkrsO8O2IHixn2ro4uj/vYSlLAaO+evHH7fZ0eF8
nUy3XzCXrFphv55Cj+tZUt10w7mcOqV0+9qRxemAuenCZZNCuOYkmxdWf6T48ENI
xu6c/iTRpeFPD+C03PpTAEfCBcmSF4atqSZrVTXq6InuvUW9X9zM7SzMyv4rsTdO
uMSFsot2qAVFhhC38of0Om3ruSv3oeVqBwZuGZvCWCPIRQHgG5WL8/SqN9ofMQMJ
dxO9NLik5Lz4dR5j5G4bRJBWPtX0bWJ7d9XFtQ7EF/qVICa6Y7kG91wvaIHjJuLg
+DTEAxbuw7UKisInYS7qDl39OcGVwpWCfAefkrbcfSmnkcP7/y8oqxZ61jcAADSo
eL3XN2Qcmp+UzPKN+yfvBUzR8KTnTucRyidUhWZtw2sGx2AQJhTIudtPlW001yD8
b8ofnwF6tgHIQJhH3GVo//XCJudgxtPi4VxFGHn2yF2uSuvIe7oECUYEKr452hCb
FsMJvoS7rhNDGXPEKZBDreCNHSs6FZEJilpYdNsptKNKZm/aT5Bx6Vt4Q4FKF2IJ
a4mEng/xbGSvVnDkUe3x9dKu8hn0HJ32On5MaNU8Nq6G4TaNs1QkA3WHn+rGoKjM
zB543qvAubvX/1ldCsND8U2VSl7I7Snz3Qz3hnYZl3WBJqYebJF73WohP8HtzJrE
n8LWWlNpMwppn1LUwXsN4MFaRn4L6a3rmJffbjJ7yvSYxEFaFc1EuBkCwprha6QQ
4Qk8HI9y3z8b0ESfvNoMrfJ1Isa8Sz0tMobHkiQxooVX5rDPvmvqB1f6CV9z0Q0T
PXlf5s1icE8sA9wjeW3Dzn+P1PzfEbqPW116DIJOd6egAiugZId8Kme0QxaLxs6c
OTj6GnlZZ/YXv3T2n6XbJMLUpVe7gYRJ3BxDNM9KBQU3DPRv2rQ4OUGrrUxtWuoq
+3U8f69/OC/z8tvXRO85NPcmBd3W1jzdMePt2G0VwOpxxh2ZMpMK4neHp7HdSLgr
IlCQOMlsNS5hIdqZC44fR304rxtXB8xpHOzYxaXF0/scBgcQsfvhsh9oaH0td0X+
ci6cgXT7YB+dO/QWiOLEvVwL6m/GCj9VwdFP7boTj5xIdHXUaP8E8IqnX33wFRU8
y+r5TiDdvEgmeYRTEWjeT6yT5dQD2aWMEUjIrBpx673NGxhXti1qbDJD8TJfrfQc
QATWKhUO7MfPw2gU5t7QoLbd0+WndpIsN//NXIzcRdtqA+Q9En3WPIwR5GW0SRPg
v8VIC4mI7EHQ8LgjGH1LTugz1PikMH6kq8GPUXGY6uxq7bNuaJXz3rgq81jcSgFX
opXVCd05mUGIlHpqfY/taqxXZ0LhDYIw41QFAFW5fvkoH0rWlWPMdNSx1puruRCb
R7QMXTmAcI4AF8ptkbo3NuTTXrG3TuSNFn06LTqUZ6HzbCe99+C1wXZIaMQ3q2SZ
GFtD7SSQwLJ9Q41NZmXIFnNZvQG4ZnEol5UoyKsOCR5uunN3DlPuI7FgDqs+WaP4
Go2y4PVgV+GDp6O9sZJDrYC6v1UPlpJE+28ur3aWhFeDWSJkCSoUnJnQeDgC57cZ
d6OCyRxDJ8vwlwakwNBGlfhH9uF8viYDQDRehcgV7qmzmh0/hNHXz5PMe5h2x9KZ
6gpuqBl2i9PNOXENEfxtk1znJ2NsiJiVGR1M/afAvuW01mUiW0LfUGPyfxlngytU
2Hso7/8E7CkwrJ08mLYwTDbURQvZ4YoZx/hj7a8f/aSiakBb2Ng3H8SY4JX8GT2j
zWbnQZwuMiftLlGKVjvu/YDlSTEXlNwLMcvKNXNReUWEvUqZfFXFoF/Cs76iqmeV
MLMlphIFWjYUYYrN0xtAQLsM9DJV3W5sNcmJouCVb0lRzeng2f3T9MOBLQ+B5yJC
igED4/Hlzr0B2nsfBXXpMr2Yq/yksevIB/aVufQQK3bd7hwlmtfH7NNNqjM+UBaj
5WpKfDZRtdU77l/7JCkR5uxfFaEo4MQ6VYAakXQefqQpWOTgfyVIXSSZPKyrnxcc
jcjTW0FvIEMGCzHemvVGEOxG6zvR6zJD7ZcOT8zbELd7aIcWBwB6vn1Ak+L/vDQ8
6kAOzv9q8Dx5dHyklQAfk9vFyqhSoicwpyeKsuGqvM51sVK1Qs1mPYunSjXJ4g3g
LSruEp8MDXfWblBC9lwItcIL6wCwAgrAC1cmwIpYFydw7KGfjx6bYbTpInmDHAuy
29LGfFG1LAE//YPLjuvNaipiOPi+UJpbPkuwGY/KOXKRTa+v6KdBe1XsyZBp4lWD
x+UrQsfcFY6hCr7KX22sQlH40UpawxBRl9agyV2OS4+naBDj0+0n7Q+RRct7yqK+
YDUlkvQRzdQkPKRisbBN56bmMncoNh2mPd8JxYRHuzOVvt5uw4S+BF1E1MuoM+xL
BP2tOmRhwEH2/gwY7vBssPbD2OhHld4qSt5AqqffCICrpgJakAreTiPUXolsSvaV
hSO3ZYEsXBBXVcDGmcsNsBsSu/01tbUz5qfp5doo0tUJHI+OIyUKNekbDvkEGtii
OKdUHYMQ7CJ/uYFzLRY0hyTDYmFHzHLgXGUMxyVAM63N8QJDvbOWxEIpUN0akBCD
VQZ5lpjKNgLXQdrKa84kuUz/RkU9XGKf5a6H9uwUKNIatuQmp4PhNq4uPQLSriJd
+yMDgDzKN9zZhTgl7uqOHhN1jZKiFVG1donBPOGVlSK8fUYAeo1PJF7CBQvUrnZf
HjFiM/+DoDApfs2aoswewOyhfhY3fi1bJrLfD5A5NGfv16ZcLtDM0Dasg3Dqlvab
AW8k2vNNKESC/ei/j1sl0uw8tcOq9Xd6w9kNNjnFh9N0GMTn80FbaiisgDC7iges
7XGMSYLCWBTeIjJqkopjsuh4DZOxv6sYPTE4trkDpIymb/eO4E/b4qde+wHFX8W+
B7jD24jr9pHtr5H/b1xxV/WGTI3wmTcm4PAJCtikWzXwK6GuKLpGjT8DgamF3N0Z
2yI3w5v25Bp6xbuHPOyJ23VVqc5TsAMRDCM9qLLYA+cIF5CKmaYQiVC7Z6as7WEb
NXL9OGc1qe4/jxeaMxtFBnlBuloYkyabwxvT6YLiR7Og2/AslheWogc7CVsKXx6A
5QlVtSWM5wGUAg32a3+YCWAJ87tLUmJd+1eDujtpnFit6+BfvDbEbyPzTdLDZYVm
RH5W+xYoAlIvZ+7NXV4++V+RmDsvphBNunvpjkAIxRsBK23Skt4wtxWcKKnZVayF
oEjLepV1obww5i0WI9UlD3TK4+C+EooVqCrXRUxvM2MMgY5q2JX0ZOuPJ6R7nauV
gcy0/Y1zlpNagLft++Fhf6bBwLxZR6dmQdKvHpfEEuTkquh4QeAvM8spxj2zPgEn
0cjFKg/F5VP0PneEidplzFPvpun0yDNhACz3Glcx1KzTZu04aPny9TznpwcYvOqY
PS7bN9upwlKQp5U+DuwoTe4zLTbocsvkoU1Ire9AKQL+XBnVEMD0sV+zFcZMrlDE
U1M36kKUkNKyqXzff1620deU7ynrAQpog9b6yi28wDhJ7lcOJPvp+hE+FDQDTFDz
+LsizncLbVoeFnd0L1gX5Ftrp0gRWmmb7N7kfbLQFVYzmUzHP+2JMIx7ZzLWQDLO
i9hAPEQN7Xv6fBK+Vp0vQqxIGojWtLyP+xHtcqGg25sEgI60eEMHQZueBOB01u0r
5+vEa7xko+qfyLgO/M+PMQ4qIeJkhnSW9z8fP4KmrKnHCwgzrESas/3LhJGV8Wrb
fhjoHqUeDEvKoIRDUXiJ73kluZ+Cm3DbCQgh7WAeWQEcQaqpfZjPS7pdx0OzUq/G
47cIjHAzWh9ABIhaHyOgZeSWIJj7k6TVbDnIOgSn+W5Hpt3NYPBnHkpbMbzTfbGI
T8luwun/fQkYUgvN0WFYaIhVJfchz1Q51XVwXxeOZt1Q7/j8T3B/oiqrhTFnjrUr
qnQLnHEBrbRMZS9EGWnluOdSOz8mLnU5paU+7KDG5GqvHHMi2P0qTl5HsbpwGsDe
Hwg4Rx8XFRAPCjHwpQbXR48amDbbprVkBARVLjwsl0Nlx+hazISYwSHKWELYf33B
Qn1P7zNU33SZ/UtJLLOpOvuv0Ob1Qxj8rTThfla+2gaAvnXcOZaXqdFDx3LQMRLU
S49aBB/RYgv4aRPuUvHYJreB4defC0y/ay6ODyBcC1d8TkfbNh/erftzAeE2zgUa
XlpYB0/WXVdH3Ye8X29FamODZYXxpSL1j9X/q5H8TtYB91uIdeVSXMWpXucp7UUh
eJYdHYqb2Ahaf6v60BDY/aNwg6QmIq8aCkL14GAvnxQx9V+f92zZhj8dKpVcAG3t
D9R9vhIgA9GebdNhwgN5XaP++HwnZklViOJpxymihbkFr9YPPR5f00NGBI+6C4AX
cJEFHmiq/6ZWwmcsub2SZl5WtSAvrk3rOcGOd1TF1pgYoRelU2p9yPWv/+tkZHG2
JetxU7mHW6fXPy+zc0eOVGbLFknEx4tMbshdZS6SQngqLiTwrjM8UH1HK1haNpBA
SAp/8Egnh/O9Pbt44DV4CA+esNGArjioYu09b5upyvctG9sdfwfhdic+LFDreZyR
sQiizA1Y2WWyfbGEUjXuCyy1E9vp23ILFzTWjpPiUnsxKD0NJfrlrsmLHeurOyxg
7tMfUNnm/xR2naMKlKbcqTdVmDKzKFXSwB9Dn+As5kF8JsLeCYouYh6MyBnllncc
QlcIu8xbUHdcTXQqDrGUXu3D8MJqyveSHsoqP/8+AMQrYBBRMOQtJDS11yF5GvN8
LP4JkQ7QIAPafzO9QYcqshvQJp+sBPKz1Q5kjp9DHZxnUurQh9mCMmKZdi1YUIQT
XyfL+JInvShNxBzxOvZgOygyYWy0lLyzwfWRLR0kwfHUPNj/UiDTWbP75sEg9/v9
MR6Zb9MW4lkk1pl7lUVkcRU/tFAlmsfrlaytWGfIBF6HEd1G9Iw5b71LGVa9plws
S60kBKr5XVM1XMOs32s9SgXIP+Yw8zA51YnA0O+dBxmWK43PXS/c0I/ec+rYf2Gd
yoOiwd3zgMVaQ2Iu9pegNgUEekdzqz0431cleVIHYvE6UpPD7DdeUgf2NTSBZPVr
mmYvCwoTdzlI3GPpsmfKoj7Z73HsG9agy9hpCU8RlnLV6MUrApBkk5ERQVlGOjmc
u8TYJu3nhOYs4SgsEKTsJ/O8qqM0XLurhdpoeOo0StHUYCwYFjMqayMQe9spSxrl
0BZ8beMokSncWaw+in+bEETD5I+WO4LFc6wMDa7u2DhTOjYyjzSNRSyiOy3HEjJa
OVmJTtzhTJ91Z84F2c+146nB7xvjQD1f9U/EcrI2Prg0ETp37y2IDvnRAKy+LbgR
8k70oRQi40sGnRXmNuPWDu1LBAEH8wIGeh3e9g/Bx1SNVeKJx3ApRpgUz5z7rqD3
WRr+dJCpxvYEhqkD3DXL72zb5fyzZR28/oskD4OCHBtQZJ3S0YOWZuW2TFf/Rwao
P7WuH6GJGNVxjlxpijB8fukx0JPPWkhXZUbCV9zD8C6wbMSf0T2tIdri1iWx2wp6
B20vIqYAzJ68xyOaCnY62WlKBysBV+xW1kNTGnxsSjP2qXlSh/DC2p6Oonw7/lHy
/xcbsi1TWuc30sSCPpWJb7/NHKj4ww2TtduAEQ7CJKLrYUkPueA/qdPYKvj6rA4T
PONc9bFWoftRmJ0f8Bi4y+kEDMShhc/tJzMqepPqbePRn8KXzMa4ftQjirmykUAc
9aDdviz1yP8n+1dDWDWoUb3WTvEoOXLXbGtaHCAGqRu4E6jXPVqvVGcvvQMCZOQp
tjuxk4dvntCiKtUQIoDdvyoLrWEWNyW7IZDncEtG//pN1OIdgOt7BHTxETIyJzHh
cv+nwK5nEtRGtusBGbR6t1Sh1pjKTyshqmZiVSOmcuGiVcwsEP7Prx/5ABeXU6FB
B6hQah/CWlzExvWdJUWu1V1tZoXDGtydwbsv2W1Nu4cuvIH/xDWBb/q85JdeoFkE
FUVIX3BVUftAw0abU2cY2npqYgPwerQF2xDtU+c4n3d2G/WcvDHDV2wqizVAUMSZ
tNEnsaSD0q/qTQ7a07GZYZ8Gdxjorn10+d9CIxu5nzd1X+sOVUpq6JcjRIiTtaKn
H5UCget1+7CwGKoKsUjYJVxVQBo+xx4kybVVQSV+0cwkfCFqqLKFnDunyqngqBZo
Ay2IXnbbh8rh3NaiRFsQqcPXmAEARQOOzU0OYEKaGkJK/W/UtEa2RGrQSwyCHh7d
Zu3qGM/KVOC9qGm+yq8lPGWzH6/vhKU/Yt5kYEpzi7enn4fJzwBX79SMtTPFOP9D
WDl92RqXOH/510qByuDULi26wZAkLCDqX7CwvDyg7ewiO1IRUchlCGgVmUArpuRH
R+5EzQyAT1s3Jf/4wSFZyKq7DXh5tbTEZh1fPIunidalEEc6Vs6TeTOTmk5131X3
UykBI61PqC5raDN02Jq0tqO9hbGRYbtHHwUWSOuPIxBXQdVj/aHwIflTnYlqD1Jt
LaB3gJcWWxmgpyCQ5JkC8H44GDJ135/Yq25QYXcCtGeLj8ibV+Edrcr92+OO4PoG
pe61JfvreCHcVG9pf7nRq6ipm0EcT+oSeyFR7Wiydk5Vn7eoqOsqya9DaMill3bk
LU8ythqbHCAb1q+5N+aT+jkiwfv7wTBGJq2XBFBcB8POFFvHbMSpFTcNWvqwVBiH
rfEYZyliCXOqPRO2rDGgYaQPUAJ77qXnrm2aQG6shmrqS3b21c5bEDjgN8wyab1Z
NHulSsl9yE4aPgfhSFEADkg3Yb5fpbIqp0yJFV78G8IQB8xFeRD5+96DizaItSVn
syRNP/DM3TqIoMrEDfvCE1oRpAljdjJswst+Aljbxjn0Tho2hn0S3SQlcybnov0u
1ltPrLOhN2iYo9N4+4RzJvPHJEyhXD+hK6MlR/Ua1HNSO68/Y8vZX5IC2FGn1qHT
6nQE08uiFWx+CbtSoa0gn35ZXGOWseJrE1cV9kRucN/tegko3sJuHdOEYFCb9N5x
BgPaWckt8Ks1VOslRweTEyZd6VAz9zu94VHA4X2OvRWpHZydOsZpDNREbL/2Ru6t
T9IrevUVCK/lpcok6Cz6OIN3PsDJRT6dkjcR9ePQf8KngP8h+2n9Xkxzx3Zfw1yc
p95wZV5fTlV8kumMkqaXqkANNupEuEfyT6IgDGNicNPojVNpiHbCKHpoKCW0uDqp
cJXGdA39CeJJDGIm3YzW2WKFPXFxx4NnxTXIg2MMOfaG+0q4O4TYeTngKCEicqXJ
ToGU/egh+4KBPKQ83yl7qJ7TtWCkn0oXZvtLxH7pY+HJdDjiH6I9UEppEwsBDGj/
ec0DFchlMgMaoMd+Wl43m2Fu2ZJpgGQx7exOjktAjXL7Pbu5f9EvfBZ9aTVQHE6t
jVi+G1csV1slN666bNRf4Xn5Eus8TVobrGnE9TmU/9s4SDV4npSaKWWgTV4tTiTO
OYq/zKlLnhQIKJbKfGuU4bjf5g4IzmvPvDq3tDS6G1+nOBP49G8Prd2GBBhlVMVE
KrUeD9h6G7QA/n6kU72UbnbHdo8alrQz+hsbgrROX0uOZ9XMgc19yN7ZBHdP2dXK
ZfBDVHT8JY3edSCmgTDp6wlymNusexAFkuIn9lU8E/wmEWLrRRBOnJzoN3e+6EZK
3WwUujo/K32DVbXViEjvRHmgJIpT8VukI/fXKs6TJLn7Lj0Ca6j1c2gEC3KX2IoS
6YkBxawkKxmRZjMf9vwP5RBtqht+alPS19E7iajTrjP4VlzUPyEQNg+tGQOG6WwP
6MXzbX0yrISXgkpZ9NX60g2UW3SW/Cj4REvJVpL+xPnFru3dMh4MEWY1UKGmMPQF
sklokclIVRHKZabNYZIVPF/ngSC8+Oin6IMmpuMPvBMv/B0BQzPp0TY4/Qlzazqy
FUDbKmp9J+xBLXEHibPO7OpeoR1GXrUboaeRY734yiI6FOSBOyzClCfOhWrQdaUK
n4lipdz3yLOvtCOQzZi0m4JDVnImZXsbpny5sYrNFlAU6rip3Ex4EkiKribyGbdN
vlb0eLsgizuFug7fXec86MHI9pKxnHTcwSDZLIxJBx0/e4dVRz1If4zKi2hR5rN6
1bGGFui0aPOaj2dRZSOguwfbp5CDGQazoj49pJ6ddQtClOuNaGQBPGZm87e52iTr
J05MIJjngwaNFoAODtwmekkpdsdMtF2oFlXqXlXaKx9RMZEcCBTfd1EJzgJy4m4I
pr3cVpUvUXQeMwJEZHVQJZtGjLA58nSyvAL0n/ruI6e2E7AeccLVL211Gu5shEks
FMK9Ac7xFxp6vM0rq9aq8R8NuN1w6WZ0laLpUzBIQgYfpczqj+8oeur4ffG8IR89
fW1umxgyfvQp5Q+f0Wc/gfM/JFI+uggrqxm4xSzxAeGuH6820iZDYRTw47bHC8LR
5l8OkTP2ouSBELQChoDzhIX8Hv8hTa4eRgeJJPm3mdbdgT2+MG0QJTclnQibu2k/
77GMXmzXMhUaE/DIAenJxUw070XYJCR7RYmPVqF4jxclZKJYdIWauY+MrtiAZck/
7JmK9D8yDOqe2y2k8iCkqDh3kkiC/eOVc29uu3wjfu0xu/FLwbjecJ2h7Bw/WgyA
ZG6OZJFiTU2h5wr7GIL82HE0Vi5aXD8SZyUqX8Xehu+aVvE3N/2D/9ycWVCeesHW
DdqLLhQNlQBP7oFOJnEeoRd20n+4x+HWGIsp+rV97m1GnMh8mSSUvwbrv4e8+A7f
9zDgoT28m5d3IncPjhNp9bFAKhnsjyAKkJpYr/czdpl9KwcvqZbJDrJs/FhlJjts
SyHcWJ+N67J9ON1oTVjKXBZGtEuAav3+WH4XsCe2OMrYGAl8U5yYnsamdW2uIiyj
jgRmXPGfRXTUYN9ngCBjdvQKZDlW7zTZrGU7B+LzeLY7p7djMkpOIK5PViYT44I8
k4CJTuk6bY5TUQzDuItTHpMR60M89+MCvSTCEvmilepLlg585jWFIyieaw7B9X9y
kpA3xHUYtzuIU0ht3Y25AwBqJ7jguoVma0IqBk+zoJbakniMLtk4OLH8NNomMwAZ
VDiQQ7ZubkjRQ3Hlcfw6KyxHVL4nQHguysBU2KghtlXZ6y3pev4hGWrZB18i4aov
jvh1BLAsVzC0TcqtP+EwWGk3nGHyBB78bhh/djRoqz6TA8jDWTHDEv6hIxwFFuGD
QP8F29orZQQsRFm486G2wJAwRwT9ps+qwyF77+KpBR37N3kM/yhQCzNbX/WiyQFD
v8MwT6jHDkS04em1gza3Z+zE9saNrVtff2qE+FyIdUcsVyMWvN3WLUtC75Qis15D
3lAKhx0KNdK4gX1QN6R2Jwb/3F+LWlPJ1sHAWfOoWcFMZV6uyOgroL2MLTyAbHmq
rDNzKU9RFnQvw/PVFiKqbLRTwt0Tmiozz+8CB7CZlNWbtCF5rXYlzPGFkVYkjbfK
5l4J7k+q3v7rpt0ZImPJtRhWpkuCZMjaXgRy2tI0SWFaHUk03H6siyVTDXIXXbyX
l0q0f3U2Jbg3cVWUFeGcZf+wgyjR7meST+KOg5PdqLDUY20rr0eawXOoTpjwD71o
yo86Wi4WyoOFC38/4XjF0OuLgQK3QVBnxtqkMXN9336mKW4phlei3zQk/7u7DIHk
eilZQWS5G/X0xMzsBAru7i5Bj2Uhu1gj2l3r+ltbCk0sOBfTJFQKV54DvPZPhceE
VhEgvkiMN0fbkCYDIEOW8IMAXhpqOeD/lXHPhsPTCGc9sNZ2tNvrnSZmKnz0rriu
wyFtXlAzR+XSnkXPvDb9mPFkrJG3GGGrKSL39VbNyzNQFLMyRMjr/k1EjI4XHJRb
CQEbbaG6JWEih++dXl0WLce84xEkecoIKtP5waT/3s0MuHHUpVbE1aqIXQdFDLDy
V/+Rc49jNQZAHxXzDohO2dCElmYw4db9t3tQAVOI7aV/qSN8Ub+K0ZSVtyK39gql
j/Elp+ZdX+NAGz9Isk6J4TBgQxmpB4IYmcKiZbynPbxIHGYTli8e1pfR0oMEs5U0
ZVMs0muAq6z++n0CrDCFt8m+nfCQxrFlMRieQz+jH43urtksSnNy1kqx+m2vGmcC
ry0ImgeHhqHTiCf4wwfWDWv4lWYv0wthnu7QDiCyLffKr4QS54sjPaiI0DC91MHy
Ng5xI86jP55NzLBF6iNYbu5npkl2hlyMOQAsM1pKM2fiuIaEfpv3+1E6f5TqyK77
nOGTco668G0JTN2ejs4PGY4sFi0EPdl5uNciUQPKI126hQkNuuqv93v3Xvkxktnx
QzrnXDIMp8RoahKjB7NVeFVtsNFrsRVtC1ggn0Wxycco3HBAfg7FAitXOCuMuDOn
RDCitvJgXTB8vO4CeWk9aW622xmcwF8ClzBojELPI97Z5V+U4H/YuY/M6gQdYQcB
AKmwWpLmLljx4NjN2ES2El2CHQlT1qHKOOOv6p98YJnl35fabMP11gdqUXgbC2Ck
V9YJs/2fuThjk033nwVyxN060sS16Sx3OEsfHeIzM1bz7yvCsJzx7cy2NGC08Hnc
9+fooGX6jmlNUWGHiFBHh2zaHDDieg7YxR+Q5HvO07UKBf7invAksMewLNoWUI+R
BCrpNxqkR/9Ge/Gg8tlIkg35R68xYi5h6B2BLXTFq1EfrcFRhOkhR9jMOYKy8IVH
Ou4C6RUQVCzAM+QDIXzTwGhNt1tKws47EUhEz08X+l3gkJMLrQj4+gymC+9/5ktC
zXk4A24fwI2OCSX0Ssa2IquANvFVxmP9v5XcEuYTpUiclekSpPhBJoL8wOGyr+eg
fP5Hd5X22Hut370vc2GdEhqmUgI+yn9Z9uoFQWbnNxfwBD1gW72a2HZph4NV15l8
FipDqYO0UGMdsrkuoxMx3EAb1iKCl0wUyevV4waOAb6X42J58Pso8+43BowJSVCY
kbVa4ZYG12mWgs83zwCz74ylmiB/t7lJ95JI4pCHPzgE9k0De5UF2BJ7VkoDSz+m
Hl6NrLM6/yjDOA7u5Wo2IR5UckrXphNCudFIelRUOWRSirmjdCd8OnD6CLOZHNBf
9d8R3azBZTvrSEdGockpRkSMYLr2LPR6Jk+5wV72OG1JeSVF/rYfirGDGTWvPZlI
3LVvcyTlY3roDft48v5GtR8H5eETvFYndAjE5pE0W8Hf8F4cQo5ysc3iEPGUqy60
h+EtB7tTb2J7qZI6HS0hK7o/lcrkCy+eKHm9C/dE4+LyfF1FsCSe5DnJYqcULlhE
zdB39KvR0JZ9Qoxmie9Jhc49kHzV0QbcTxUOkbqobC+g9a+k2aWX8Tq9U7gQ0leI
IDZaC+6JKxmkMRoAJqM+3vbWnOuODEl5Llww96HHVA5FDqgaNJx2A/iLQDChK+QZ
FS9Brxu8TsYe8JTE0xA8DwR/4aKLeomU05ZahQdwTHH1T3VEvoRMX9+eDlBrVllQ
KzL9r2WVIINi5sR/7yenFoamZa7sYaQt4vc8aBuVaDWG7Q+GPp9nNdEn2WVngGy5
I2u0UQCg4wj9IDQIKXWwJeZnv+F5+qma3DFqGkWlWFWXAne7+vbuxeBtvFzdktYH
okkqC6v8O7uEnKiIxZAPVmjtU11J7tELNC/XZB6+ntgDSDFfxLvXy75k/t9EfGJn
1e7MeWR1WhJ/mjs2plHz8NfwWsMG9d0SsQYsIm8VvuXyodga7wfo4psDL4wOLgk0
1WB2c/0t6fL+VPzAmYze5wY4b3RTG7/FT3+UkfjQ70bLyC68N2aS9CJt/xbyu6td
pM20C8DDFiK8UtDb3W1YBiovI55XRTEpR26A/I6suSsuon+XueKjoF8LvK60bV+Z
LCe+gtSatpLPenUGqO77ejDEM+hZ7R0Em3apSeHLwNvJiuYWkMELDIU267HNzV/R
UthFfCrppMgG++JI1LjmBRto5cTrVKl8RLH2Ij0G44wmSg2/OzE8UvQ5uVEalxPT
J3uRfex9qYfDJiH4odRhsEOz1+5iyZayd72T20V0w2MGjJI8lHGxghZ02LKoopOa
MQDX8HKe5USS6jdJubfj0IivuxIfWmRHW4Tfx+rsXSSupPT3nq51wUcfKJhqX9CY
9m1OVuIOAXOhw1Ftt74TuGtvQP9YhiWhfdPMCjs3yHFAwFL6jbTk7aiI8xOiUeyL
QBkBtUN3rru2eStgycBInW2AsAUzkHc+g3WhAMor7hIqM2Vs2kKKoke6xH5BUVV0
vJC5lGFwQ4Kbq8ofPGWrwuELmtaMZol0yHDjh4zjpGRwXW+zxGDR+QoWmAfYjgwF
FpX5UIiUPbgWc3F1QHWmMWx34EcncINfPCnTcITxxq/lpvVlreDb0Zd1VUBAc4am
ywE8ME2D8PRIxNahg5LVjpqM5x3bJ7Jnq9CUHSMLctMiUU8+cW9Mzfe4K/ggrS1s
KuYKdR6h1VXY7NTHDK/ki702rNO48K1Vla+JHo/CviFHex1gbtlUK4Si85/6g4oV
+cxrGf3XnoqwDlDNIsWyacaubdAjS4+wcufcvv9KJSd5F8iFNEyLSGCKHrdtSKGe
S+gA/VIoFm3A0BC0Awv7O9z/84vOacSR2BOS6uXrMdHrWbfc7eYGq0XxnXgFmZke
ZY7gJ+xoMeXn7hmLANf5aTcoJtUOVTbruxoL3ern2SchHE8TZvua9M12ZN8+0k9x
1k8xEXhwawH20sXDtqrLh6bcLCJ20j3RpvxaDDhpmgUR1zjfsA+Gwt2gNl6zkrzD
mpQe4Jeto/jhyDwIDsfTY5+xp/I7p65lyOP4DlrY7Ncy46iTcYGrFaEmb3gRDEsa
Pw0nao69MwPjW9tRRMOlyPjh/89mxtHL/UsVD7VAGeWPt4BZGxgvohdLA5ukx64k
UGsNx5azSXKhyL+o6lbhEbNtp/7GPrBBjG6jD3m6lWbz8h2Pg6njdv7qmXITF3UP
OsTiyt2QDI8+EqiY9pLaws/EupP6gWl9fUU2DWmTpAfO5dmb5jm0DNRNebUOpP4Y
KO/+P6Dy8v/BH/FJcDvqtGjUY7s1heuKYslEZJBIvHILd6YJvG72SmEvA7PJks1M
WUHI8I+WqJb33rATp0sFgIVY2dRV8IgLrdvDmriN72q7vQjvNPpCMoZiBUb/FR7d
UjyjsO3wLzV0AAZXNkuNs8BQBRsZ7C4djvWxYyu+fSNdtOwsi0PEHmIQ9oT3Svp8
GvO1NQ4VkwJktHysu+GGYH3dB2sqZmhhiHEF7AoIsf9SIBUwx9CG/R3jOdiBHxGH
J6KFBFuP4A3AF/Uz2kzjre9oA+WVhSW8eOE2V7uiU28ocX37KQx9Kh3/xm0bb+S6
X/ZLvRUUpaJk/Pk5ddMwIHsR9CZSsALxCTg75pUcubkrH1mbq4EbpWo9U3TB3h6I
7m+pWZsr/byG9Vwhvc56P3trVz6wTr1gF4TkIgQFgIl6Ij27MxRR/LgcC1dwugTH
rOjsSP1GGl53ilOHFJEbUsjN5urDkebJyi+VJGnoiunD9kTMlqnVed1C6UguXZbh
MHqJjPHBUNSah7Ebr810+xxMqDKdUNePpDK2DekfJE2y345U72Bh/F79qBIzM4pB
2rncjujCfB8vur5qBu/zoZsLwWmycHrQRMn1FQt1qoADG/RQDVM/rF6uGsbcor2d
+fx6pu3/kBzcOeg2ySSGHIaNXsBceLF1FPKl0rG/BDY0afBZb0qn/82z6ml5PWk/
+yox086xSxDkg48OTpeUhmc//G6b86rTRz6U64tHGoHVvZxIUWBBLISZOBux/j3a
tFyTGOcsFaVJhHTLLfucTSI2PIZ9Im5C9SWzkwNyyMeaWqnB1bxxmKLnDKFKcYRa
eIRxgv6gX8m8l0DNuVWNYkQ+qZLH/VTdXEbrnRCbUs9L0Y+5Oe7ZiJKbXIRyQ5bW
8hJfvMgeNuGP1gTbeZQ/dQDJ9QNBgWJjXjQh15DBGzG4GbEp6iHmD/oKbCFvtn0o
fxzE4MhUwX/IG2P6IhRzFSQTCfZ0oAnTzXMOnZUR5ZKvKGV58XYerUENOQbCf5H6
nwXPyG4n5jMRKaatQ8GtcYK+mgUYrryfCl5Jgya4sncdrZ8ZcNyeiISwuKI5MxgH
nD1xB1QV2UrPDvwxh2eYWw+fKWwPL3SwMNHOdsTUm085xnKDmpisZgzOaRoGM28p
D/NCOMpcNKnSakvEd4QIhBHBN8znDx9G9nbFD6zL/Oo3UZ8PpD9fibLTaftG8QjH
G7BYyND7eWmLPMSxWnUc+QwCEUCctHtIAEAEBMiMzqvu4NDDwtEVdIG7ZqjUlh+t
l6LIWT6PHNCHhbhZmqicbLgfHmCc9o7RbErOMx6Omp1Lg2yxnMSCBE1kjEkPg51i
RHRI3GhFq1fGA2ecM0QGBgmDlZewRGnoyCoOvuqhK9fD4xb1vQ3TMJxdYEJQ7uoh
7fnmA2/04238FAhBsXM/GMvvlVUumpaeKLEwjh7U01ySkjqJ6gjH67a79dHHy79v
3AKto0vTyD4HP5Nn+WW8AYN5uWzCEIwD6DEHj36Nyv64kubjLILpfYWKBJS9ikqN
crSBCD5Pg/uTlT9QUWZ4s7l232sd5I0Zoc2RjNzy8aCvPfvbeHIbI4glIBg4sjqN
KDOTIytR+uIqvrNTQk4OCZhgsGIq+hAS6VF+PJA6FZh5rDrWeYqaEwjyyChFbVg4
ccXOyLTPVwDlOq84UjDtHp4Rv2WRtasuoG18MSMX2BXW3LsC2BW2PLEQrihu0a4D
hDuIGf4VLv8LBFQuyY3agdw1JtCe1xmMtKLgwIj8yTfgmoZ5LuMVGZRRK4+wmULR
JLf9i5hAgmvzu7mpB6uh6dGeGHAVdXDYdNqjDW3uxw3Y48CVqzwEYTSqTjLly9RF
3IdmwEiqZh/9uTeYWYgJxV3fG3ghUYbLQoDdTbDtuOtPgzMkZW/ae207rdCKb7sR
qeO092fmYAxQ+wBkQ2UfhaJSO4EwJaebcRg71+MH/IU9wX0ZllayrIurer8Wpk3D
erESrDyWk0PPIFFYFmd1cn7cv6TvY3lhK6pbQyf9u5TYrfQRgSAJiADotWioJHdf
Q2W5TUcXcFcIy/Bd37WRRsDjmFSW7rEka+bmntJrluDXgk9jL+vNnKGrovTPKK3k
9V64TnZ2MTb0HZsfqXGShlWX+bXW+DDyZuzBczpMBGXmO/gus5+Z6qOhO4EXdFTy
W//I5xQHvq9wbtKVBXK1c885JVYFtoF4XnoZfGsoYgcSNfjPWb5xFhdxNMXThTbg
Dv+B+dirr6HFeTFAy0lvEt/qtDi5jjguEQNRAm33U9LEvrHLeoR32sujikGhXoQe
0pFT+Vm+YorxowSEWwKsqTE6kRRpDjAIkW/D32+ay6dE2Yx3lF0sisfE+lwSSVUC
/4zd8H11FJ4xSwAkL05Ck2KGlN9gM8DkezxNdnhqv3pYN27XRZsQxOtIS8w4Vrt6
C9DKJfFJC00bNKpEzgeIPncdQC4clmIrBSsbYgiH8+aIocze5o4vTpD0Koh73Baz
j5MOsRB/P3XT4p2wAp2KpT99g8BgX2SYiTG/J7fTvapBVhx4ncHE281HthJBqR4p
3UNm/s5iHLz8i3jAAuKIisA0WavOaZ6piBGvVAvT4QZP8+AMRt8YxzroYlbZgdGU
cJkKIQr/bVKrXOYuGWNliCPeAvDosubLFi74xCDkHD1LMwIa9dUbSTijzZhl7gYr
u1diEpKVQiilTALM88qkryzm5sf5RLHJrcxewVAQGp4JGddkB22iY9sLLN8QKcQu
rUSLAAm/YGqZNFwnplGokXsdB/SzvMWsdXYvJRMad+7tgeUsXl75D3XYw9MJdV58
OJtTBHDpgdQIkn5kf1xyaB94a7iNTIZcW4mG1UaMwNKLwstyVUM08IIrA7NYyHeZ
KZ0ypZM5Y+UxWegFqllyhuR6Yf4pzP+atrWJhwY40pf865yGqlurDDnlpufwhVk3
qjRFK5/UcuiBzLueu9jrYyllBwbfGy6bwmnNUwHNuElUeGWvjiyeExnVCXbkusGL
q538GWTLSp22y8zD2F2gGQFy8vQD77IKzynB7ts1exYRpkgi9rUl6UdjBGkacona
HPNYu1Q6cZtXLwFxQtE/wGUfJKjOuCv5I1gRx7jqE3+9h8X+REZsKKimUIp+7nZZ
NWch45YB26IOZ8jlUuxK8tM47YkPLs3hFKOlLHc7dnDDFEBuQm08cDCngC5uHI8h
eyHqnofaEvS6baGkE/l4PshSWAo20kX0p0IcDekJsx8jXz915lpSdQpt9rf2uQWZ
vvb9aof4+n17akHiPB3af/v1dgHdR3JI2LxjYK9Ed7ehi6XLzyXixfHNj/E4Xxjd
GqUkAjyVYxwEzwtNaTCCLmaYvP6DFS+WnegN2O01WIWUkpZ3JdzTMEewhmKNbVtX
4/KYoWUvAtovhlSHuvSaJeqGCVRfNuKY1tmVjA1XFqhaN0YAnonVM7cnqoBI5+Gx
MXlq2WTKRqsdi0Ly8Qio3v3wf7vC+uViD7rcEphX3Ru2ujfTxpsNOmjPwIa4YvVY
FaMAmt9et4v/aAJzvshnBGPzrmVKaEKZj4zTyU//amxgcPkOZ4l1+UBwbowIQcao
9TNE5fJvREQClWXKgX1NqbPdPDoGp3L90SeJExKXm+nCyHVEqd71wqGWnR1/m9Hn
JOu0fVaB71/P0Ps2lAZNSsApdY2CM+DP+S2jjloaqGnobogNNzBV7bl8aXAn7YX2
VwKfhk8kmd84yX4OEsSrQZYjPACkrMsRc4lox3y1HIXz8OcFKfZSKHS7gMFyjWXb
zxbyjP7Rainp3w2n6hkQptCfoBnZ1YUzAgdMAxpYfRzv+1M1bhY/C3RXr35hW0Ps
kJUN3pZl8esztnZwP59bInwJ3zmThZAC6qhWa1iKoLP3z8cNJMZ8pLukEfcsJp3k
SZtRPC79ITTj7uwi67MDMVJUcHHn2t1rjwEl8mZ3L5KoHsGwra7yzezVU7QyQpUc
1jmrU+R6I+FYBD5VXHrnwUqE0nEt/XNt4rcPdj6agCzSAbnee96rEwAsXukVZd8o
YHdECVE92U6c3vAA0BLuTlSX/uGtKVwkgw7v+wgQtFllh6ov+TKs91RU3YRIorxa
INE5NvwWoA0llmuTMkHcaFL4GqKcGRrMpt4tN2W5+F8dgAe1v/yLnvSur/RD/K21
OOXuG/Ev5z/5bV0RYRZ3oCCAx4xYzNojzMECssr0bIdEyeHHUFxd5R4RrCnz28N0
dIxg6R0+tRR0fdlzHqR5HQ6+EyPzMUbnpNxF4b1iUJvcFWJgWSTQmFDRkWeC3U42
pakt8QebIqXyeAdrvgkttGj7FY3Wd2LO5t0knL+oehqHj7jQrKSH19ZbPUfEd4Nm
QMAtObBeMUe6kRCGpqT4XzErY1i0r7hJM3Aw5DK8DXX5mmXRJMAhEyX8RxRrfrDz
TzXfVpv7vXCoywkUnecG48FTwh64+MTbAhEb5CZQ07RK4yaRLTT40w8DGmMNodYI
fa3DyDJSWDkoeJubtxxDL4mjane8VL3SY0q+jLPb3NKkCNoV00cKmhimz+Q3hC/3
bxVf+fBX335PC9nTW+pF/JEnHxfP3dgc9AvNyt4VjaXC6uJSoy4tzVuwNPyvWXWD
fveUYQff1iXTPgaFmvnErKiQ3OvcZQxnxpzG+LAyInYoViOeCr6p0IIKR5KE0mZB
eF+lAjP3uoRL/t2toZ6vjj3RKHPOY8mnTDrm1fk6XXOWAVG/wDs0V28cbVnyUobA
GRz9oy/aoWQgsg1Vf5FCSrQbDOX2AYhBEL7aaTXWEv66CGXzlQ/F00L2TX5Qimi4
C5LDAo4DzGNGa/5olCva+JnGTVzBbGftnJqZw8qgfPZmoYRkX2kKtO1nQBRaCbfh
GCiRbAszetD4OU1vSXe2mhbfUtcCJH4MI1JuDoSWVNfbu5Sp85Ym+65Rp9sVHvZB
I4zkLCF/1k9Vrehb1CZwC8PD6qTk6eYEAMrEjWKdCTSekHoHNdVxwRFuxYFmPBjf
XtVfVnkhLih7VCKEECcqw8uAPuxtJWFRqvw3hCEUrlGBufbPwrY9aRPBL86yVkdE
ST+eWKsxpb/4GkJ+0d0XxXh/XwPNGoso8ZOD/ZDzXzwsgufpwbf94iawPwZAYa6o
5eM1C8bm3d9rzFSjFBTKM021lZwHPhsj5k/Q5SPkEQXlhZEXx+mhXzfE5eI83AXD
adqO6RmT5bJ1PdrxIztCRyvjiZijb8tYj5oF+Ys4KobuN9wfhpvV5Go+GXvnrEHE
XoqdCraN4rlnCODqywF1xDAUVDwpzL8WAKBtdjii5nzCUOafo5W5EmYOp91qCikB
eJaG1Uk8UcZEVFkOoohcXE3VLGHeBViK3bhbWcLLx10Z7KTsZ7hLw+bfB1xKGmZ5
Csvs+vqB+nAKaz/2NZ6vyCwrMpoUbOmEGXX4l0SOjOytmwkejdt8LPZUhlMJcSgt
OMy4J+NebdHKh2HW1gq8wjMODM+TtMK6SIu2/547OFRbmJFqHaHkZJZ+nwXXPb36
/6eRqnn0IppL0RQ63XvSVPc8hCtJHFlcVB0GRQ2QgqOmGdo8hTLnMvDCGr4DzQI/
+eJxpFnGZ9ttyhx7I2v7I5oIjKwQPN38JL9+wdvIYhPJXYkP6AxdmUpQIIUjcUUN
b4d8LnOgVLxGs3WXsjvL0/kekKu4uQc/V2gg36YMm3t5Ewp0EA6jJcyVRq3soEUM
UL1LS8YemeQGJevcTVrWyPRhqozBgznu8D+sWzufh0a9noXcON9NmixqI2y6Hely
StwhvuyZgiNseZJD3d5JFtvSPwFF9l6QLOdr6xdANUPsJgWF2atMHAvdETD8BLU4
CjHQqjiV4u4HqGn3V8krRSD0rxbM2KjFhp35BVv0Cg3vpAI8rHbV9pJc2mx7n7/N
EtnOsmoC3uZ47RQHbepDMDx25VFlUYp5lqy7x9Jc1e6St2pK5CIG81I+I0/deH2B
trSzBjBYG5Vj/lc6L1lMUNQknFk8DjBIJh4sDhiDJmEaxqG2QjtbccDQmCUsftXT
cpXporxM9bw+TRPMLuIGjcZ/pFinRmK34UIFtxik+HmzfwXKsps80lxUNfKJ0C6G
8WskGdNigLE46tbwrs1D50jHu0FUQzpLN+NRjFxX/xXr3mKpo6ShKR1S61gwlWRC
5/KdidwLLI0sDDV0RqD208HChdcLZRLXv2TjFAC5nJIxyw4VX02E6SnFDW1H09zy
Y8R/ZjQ2sOZVaQ2R2jdIVS/76y+J7zxhljH+O5RRN3dKiFg1yzYj7aS42HJcBYfX
i5KPe7uEiuepNIwLDate9HgCMT3u07cGaALK74OCz89Es/LcLAqyKM/+e+IDlblR
myOnWZcHR5n06Fx6AydeNnvFSw/wfJEDuuNn9257glLK+oeGe1JViNiSkcG1o+1N
KtzuLya2/U5c8XNp22UmYcbhAF3kB4aX44ycWFO+yW+nLWGDkCuZyMkel2zdAQWT
qfSmEnIVsrgspIDNaXegXKPMDUupJ/yd5urSVADrazhnv6edlauRAJcmEYRt3tNr
YW2HQk73n/0Vqek6SHlJUQjBHgiT8/VHlRHVDh6lGl+UPfAaIQjJEB3aNUo3oWk4
wAj8qBLRVe8h4aEpJH/NtYmGZ8s17p8xEzSgf3QQAMnqq7ZprwF3zer41gldYzMO
VN9f3uou+y4sedHaWGdWgIZR+x/+gGHUyN2UOSsjGK8ABxzzfZLJBdQoJDG62NCx
aYtbk0L+Tenm/MXL0S0zMDGegxC4dPEcMpMGpNVlBvP6MwinTY8SxWHeD17oV1H2
j7PQ3xPzXTUV1CbWYtan7cGBMqy7OwisntikXw8XoWTIz8bHOQpdzjP/6lN1dUs9
NqjGTQMhiG/fhu80GsoQ25Us1vrMlHMg/bDz6lkvRnNxrIxx17w3IzbDmRScvenZ
OrrMuDerQVXGv2ZaaA3ZKaVlt6dYSshb1LoBwSYYhTJ0QHbxSdva35jW4GBpUtxZ
iJpfOflr8yMNGNZ8Eqao/iLgxoVUoE+Fz7XrXRJdlDbOfh8n2KwtQ3QQYE2ylJvs
papQNJ4Qp0iv6IMO/Jzm6VTg3skp2Fz6fd4JC47y4G14LZd3fgMp26ksw7TSjj+D
AXDdbcDyBuI3mn6PbNt7KRkeI8+jK6omxfqjdGAPXrDP78X702tuI0nDbHho+qUf
o4u3HgsBdU4GGPqO7Trgm62UnGDiipMXp4K8oHrXBbWOmQV6DgN+9qgvNFJsIKDM
BuGrHXVS9viAjqlLMIZ4E+tzvntcUzpg5Tc5uFby2g61ole6mngRcZMwlqmIqUms
v7x8neTWWEcioXq9wFrO9smWqX7GxYf9eskMP4UWwX3aBTDfHmco0RoZ19qma/9U
Mu7gIUZmP4QGt93x95+km6XZrd/+RJPQvx0qI5YN4cJLUvYOaBEV6zIYxlhj45M7
I+h9mKpFesOczJlZ0G9Jk+pGw11XOUfhHDM10CIQx90GWQmS24uTO6/HniSDZajt
QMjrTh88kuepb+qh9FO0ml2pfDbbHLmT/ZaaEyauUBDifV8G01ztxjjAUufSwA2b
erbCD8iLTzmNqkf1RhiTR9057h4f+3vVb+0S+ztSKVR1uumqThNkKY0uoRgGXHnU
42DAHKgZM9ZC5rTj5Vz8Tn6I/lf3iyaAXeTBn73BGmnT5hlE4Rpbt/M4V85nnq/H
IyFIQYin+3b+engSQ1PQPP3S68df/sLfrN/LDDgFCUyI6st67HlHilht23NFkKmb
T+REgHYEXPjLuUwomHUfWfJereL69b5R570FUA3gq5FKuOT8qD/w8ujBLHSPY4gz
uH/jlVIZZW1efeMOd5AiQmy7SozT2Pvxi77eh384KjS9LTXR/uBSwx6Aq4rbc4/7
50pIdrcEx92ToQ2LE1DZxYBF69IzoCoTjgjjXK6Da0VV48Bn2sovt0zpuP0Z/fKN
LYHpro7m6NVRIErUaMitzIQ3S/0SrctD6maRdTteiWwmtwNd0jJ0aaHJs/dcENRn
gpP6yvoOMJXcGQNSMm2suOsOA9yl9nMT4iv1eBAgZQ3SsLohnEjFtDKzMkau8DJK
rV7SEzr9EsUAJV07cNWYlcigHC3iU6ZOFjC4H/JB8zukqC6QTh0lpEkIobUJUzam
aABJjYN5Qz7vV7dPrCHFYq+/IXDiKq8UjXRLZhBNumqoOB/l26PxeL2TlkL4MNre
aCx6xR2kMv5waY6Y5lWF2hirxHuBY8WbplOYFKKhy1YjmhENEg9g4fzljwXJ8wQQ
SkHKTtx+kNCahS88r4ISocIXhq/U+U4UN/P5kkWEZQpz/XCInriybl5cYUsVRTAR
OZw3WfA35AzoFJ0Gs/ksv9mSKnr/GNQt/Sl+ur2I1KEUmovlVUiQWLLMdgPNT5vt
NG3OZ0DKkjcRRw5c5rWP2FqCt5OV+xwAk6n+XvPzdaZKlxbL6vnkBqSG3Zt2uwEO
Q2SUdo+HZ8zHcQjVfwabTRuvHgOpTeTvJx9URzcBG0qthd0QNkUd1XTsiVhKo7vJ
Mq6gTrq9OUT46fplDvQqzN7ZFpAxoleH55gmJXt9w+cb9EmZ1rdUyiNZjY7uTHfi
SdHddhx0YJ0Pdw0mlcfb63YFPJdFWXFFk/ZrLjC1ITQcunghPvMtJLPG3Jm+WCYr
o/T4sdIsM8JPSWMg7AjmgsIk1I9h6Tux97bSVlhTkQsKxHIm2aETqTF2b000EUOi
5ILSxa43ORKMTxaPJH6jgwv3ja3BTTUMhMWCcWTGK0TVhPUn8LrEK1O8APFgVUKX
V3MKQa9Dzv6cC38kJtnp+mcsBNa+Ki8oOB7XuDkn0Rjwe5BjEs6CIKZrlX7Tqt9r
req89uLykG+597k/QPnbk0nA4bF8yckfeGPYEcCk7fPRvafHgY/tLM3mr67os2zu
krRjm7D9gZQ0mz+CdctZFJ8rgKxV5f/A+eF0mvszOqk6JlctAHiMCT1RbyoM5Fi9
nrK2zf/zbltX7HD6luUp5itv0P3+dz+u76BPdQslRRFA8SxHvnqxpeCAFMre6N1f
D/7atYtgIHeNnO2zQqJz+OHgOqAAsXU6IgJs6dN5R6V6jnlZeAt+WW3Uhr2s9D5/
6bxO+TiwYJQukDZvtir48LLvff68TWlD9zfhc9na/ErUtYalj6J1oayoQCTKlN1C
vddXsq7YJ7KqvlA5iyqq+xh5RLmzzvqGIMld9c3eTONwuR02JSIwBxkBB92U8twn
DT2OVf8HoeIBUR+YIQojy1TGYeYM4vIKr+1/udKJ+XuSA9vVurxjYXuzK3aYT37k
6eUih39WVaF9iLkZH6+ItybPBc1lw24fM/VJQsTyxWAxWc58TStL4MR8TaEteioc
dLOTjS/J8wjS7T96+Ryh/K3NEL8UhYTPKPIPexV39u/inkHs25HmBEY6tjDYIi8v
Ydz9LKsItXw2t8KyJc+2Va4ky4NatP3TiC36E686Plr7GetthgIp+pHUTfzJMf9P
cyMY61Ika9zEAFITRs9Lk+o+ZCJbnRMN3t5X4kg3UXFXa1J368W8JD0DNN4+G7Bo
SLRMgcBER+mP6D1TOmc4NKh6uREh7cqWA6Zo21t9MiJDBGo1Ue55LMOCtLyblVX2
llQksGK4fV49tg9nEip78eqcRUXM0BFVQDFfjnGoninNU52Q7hv5giJd/9IpNKPJ
NuPANEEBLCsksG7tiHGpudPL/tyn1p5UIe8Li+3CLhKfNej1p8ghNbXj4jJ6wOhQ
EE2DUQ9SON6DJDxzhuqRi1twaTW0sD764fAtr2H/Vslyma8j1lQKMbiGdI0hIvAy
KhhwFUGJgV6YCavC2FuLpQnwxE7AJRj6uXH7wgb4BTyjJ+fMO2Ip/VJcCyEjvYsx
jl2ueahIvvdxWVUQnFmYcn98z6somW64t5YS1zM6OOjhZqMPRd17G8r8nyvuT3Ld
jU6P4POXUvCvKwEvKjUtXw8Qm1CdJwg3ojNpSsQKZ5Ftm6igHPOn1ahDs8rZ8N7j
5TJG1QleXKafDd21/J4rGvmvhLE3+qV1HG9FPXcllz12rc8fxcB8XPdVsaSya1rF
svEzofGS75qrVWpvZ+OTlHnGxpHGPIGobG/j+ihSnHcWV8owo8OW+zyoyVV0G6gv
GlAVkqiLe2erZAMx3b/+Avr50HwXowYhCs26yxf/8Nb/XXhxVJiu4R2BQa0w5TlQ
prfbRqaCmoUl6ixfuizRhSY6CIs3zWu1RxWpEE7SdZcTbmssFN7FPDZ1dq7f5UDc
S1nh+TowXSVQ0AkZNjMlzfMe5+A5R6w0K2tselwduPw4CRF8E9LqzitKtz0kH8Xo
iZ3MnwAc4Zd6YOgfiA7QiIo9dmHwCvTbySISgiaulDxDUl1480Fv0Av1HMUFJtho
ZS0RIXhL/0pq+IGhfTcFi8me0ZDjkbCvwijNqTY/RkLyS0bB/JgK5C46OqRvFW6Q
7fpYDGrXzAR+bTD2wXGLsGf7Ze3o95skKWHr55pKNq0vi+sWSbZYqklhxXRudjU6
Q8prA804VMylv9X/ql8kyjjXilvpFPUSpYKeAXGJpblhBYT4L6ICkJbvPWRJ4NtM
BnH/dGJYFftSrF/ttgAmXVj8xNVz4LyMkGoR5EeIFaLj1QwsPYUXW1f5QJEaU2Wi
boIDGmuXYvHsokE/fpH+0V1bS9ZLUDbNAgwyxczsBLsnAiTgcn32PntETmJpzeqY
GMBwxiDmsXUJ9Q+8t0ZMxwzRZS8I3QrFZDX8D4Uf4wamtS/WtI+GhOByui9/1MZz
L+KwMp3HQRXr689CD39vdCOBGGacJkGAgIZtWmosRkF6254EdA5RkX30KrI5Awh4
gfzes6MuZEMNd/JKlsoBGmHrWk3XRxpmJXGudfk4DN5IsnuXbIy1UqiTpuDXphtJ
FKx7JM5nqQulW8se5diaQyPzr3XdqyKkWAyo1WEm6XCGUuON4KeafTZeU1ppaqxr
bkw4OJTYOQPIhfO+ntZpZuAanJqUC8biFgBEWBoSL/tGCIj1n+tdQKVfmVoDMJtQ
CROexsUSXQAHSKz2PJ3VVMAEZtVvYsGCKZ3mXACdcOFOXjuZ+Gg9zVl9owUNLuFA
VRPISZY8Hzx20OvyXDCv7HNxj26Ewy7XSP0lI6p5k50hi9SDT+OWYXsldxMHq34i
OYu1CZCUy7QkfVmB/LcsNfvS9cA6R57sqGwcW2+zqG7FUHKuFXz5HwMXoTsb9zcf
mQvVVZmWXz7WPZnuf/flNvvxzfZPbEIvTY5g+AXIxa4QdLw7R/0Kysi7bnzTSSlv
0XqO1VSiOENBsOBVRQXS0Ka6d8qceMCbRwohD0YG98om/0993RUTLMNYSqeayzD0
6BJDzElkw8P8D2o/U531h62jwrUvgLWvbzeRAkgLavsrEuLBP6AmVhlyE9FAYeBB
NlMwxRWsCobbacMbHCORqG/mELa5Sj3Zkz0Xy0BpxAWZ5pumDaSpNepnw+cuJrP9
7ENYd/dO/eS1mUTEj+2hD+cYrLPK/Z/dwYYnFDUddAEsYBTsX68qGFMaDsRAWztO
StjgQ0NGveSIb6GGx248NgAOs23rl7ZKn3SvpsaCYNE+ll9qtLkcu192nUL6ZPdu
Rc2cnVxRItWTm5mK/b2VWS3z43qGlNpkiePptyfsA5goS+DVXMWStnYkK414C4Pq
zS/oZmNHvdMVKLeKFjhPzm1RVfdI3XUEI7AmNSXVE9+ihgwB7B8WiTmw/llWKg3b
tXmPqR3mIeykhtZsm0vTNhNRF5PFEi3tnpNspSiiHcoX4jLH8gG68Y+YdYw+SExD
YQ1PtaHkAkzo+vGx93A2k/o9t3yPHREQkqn/zONI4F17RamTnA9/h+PrESzJhDUw
iwm4JpBl0n1LY8BAPoH9nnjCF+OLsUS+FwzkWNwjndOmQ9btwR6hei6Jqt7So0H/
9FPXKwy6C/5utoFSq488mTmQpXFsRtBuMsmsnoauW8ZoUZTOUn1QCLzQBht50Ydf
6sIDIiqUxTQKdu4q1frX2Yqw5Xxv+cXNacOMCx+KxAfAawpUJhTrdWySCxuWQBQD
vHH2G+FGQArTXnf6urPqbirVI9NpzHA59qh4TTSi6joplEDuvSNJadvRmpZaygNq
VIaWUmjb89kzeCjHg6m11+MXzvViBhvoq21IFOpyKMyUvq9/mnOTY/+NjecJxfAT
h/ZIb3/7Jem7ZLft8Ov14IJe74x6iD3P2chSQyfBk3v4sobPi7ptDae7Jsfioz4s
ggmmLGqbqYS4yAqsBTq2h2bPSdzV/gQc/gDdDz99Wj3W0J3ft+rKjHDV4gYuOQZB
SJ3D4AQUsoll2e3ymiFpt6NZMyGrR8J8RFLmXGyKmiaUtoiUF/TW+Qz3Eyuyj4FZ
H3KaNbAraeLCAoNk4MJG9H3zpdlRh5wzv6j1+2kK5h6sYdPmlpzZsEBRP3mgy7np
HmeW9CH6stGGKg9dKvXxZl/l8arE7pnmCpdf15ohaKCruyFm826lwWEUVDTEflub
nh4hqKUMm86HAaZp2fdB3Di0WlHJizCW6WDsc0ut3/z5LlE69/E28t+Ht6Rojb09
euGJzfTiGC0biw8g+9eAL4vmSXykfTllbmpP8EhTgRzXajbsaof5v+4JFygv83fk
A3IEflgJsXVN2y2dzjo6HiUAFyQAlSexJHBkBUUnpnBwWQhhQs/Pd6c+zAQv4eHg
GHAUnE9ts5ZyUh5c9xTlUBJBjadYj0A4CcXP627RXnTrIrTnO0InUefQ3bAgEY+7
WSEefkbW0W2hSgwdqCtwoPmv70GsWw1Ov8EBMLmsa5cZigCPEEBJ7g8sxaBRBxEn
ZfLj3GvPP6lF5DdI1w3Df8DoEhXS4dwysv5OBE05yUktip+FZtHuZQiedmZBvM6l
TQETb5SRAaGeMgiSYeTrmNd2R7VYejbPTxtFVB1T0AkAnHlwzbCtoFUoRmfClh6k
fcpz4kWqKEU3XUOWFGPBAyC7WhEMuLibU/W3BuWfMJB/X+VGmqW7G8zcaM0KlSRS
bggknkgfQr0jFq4D253H+mffHU8X4wCIz7bZsH5N6NfUyRgoIjnt+GDZnRLGjPW6
Cgcml5qReJ13/n5eGtxMLIWhHFBG0RO5vuPFY3IvwLYsqmcADj+TXGMe5G7G8GLS
ABAYlOflOFBrT331UKn03TQskqEbfUVnSVuQKRclNH3Ibxu9pQqvYvS/hcdviL80
GxXgiD3wlPNByWsOojXgUzOtAlv0mrBYOPX6kWhsV1SLbGH/EWRGftuh+VkR4VKC
LKSVG2m6iUo4V5Ms12Cvh8VXsZyIqAfDrdQrROWUxGnlO1q3GR6gnDUQttIV/LVn
EDcrk008wjNHhzq+aoujWQAb68qqMEZhdMOXGg80iT4m4djytKWD2DoK33uFBZa1
GX4e1fzeZXysF4Ci2J9znbZ1lTaZLh6Vf8yiB9V5OInx0zh2Qpqb9Qt6lOnXWTXG
fQicIuoRshymv5CDK2XyNA7wc+rlPeWnJ9Jpi4LB+Ykj6pNE7eAV9I4u5XNCbJJh
JyOB4H0SOVkqgqmR3r1q0yOdvJNnGK2PDwtGck3h46YYzzuh/rZwiSx9ic1Eashq
HceuDihNVY7hUpgvwIbMDusetSKghMn9ovbvwChSHDyd5eIIdw62xvBfdjuK0cUQ
hLBRgaf8TwB0+DUi7JeyRHAlYX06j8siBQUef3P0p+yZQp53cfCui4gB7dOLr4/+
lM00Sd1RsEFuhp3WXuEgY/5lZuaFrHF3P6I4zQp7gNKZgtIqGgFE44xUtidWeujj
idHYANoc/n+YXgOGrk+CJ2fcKZ7JBuhdrExADXKC4YIHjb1cD6xqCHbhQ40ZvSPz
yQ+7LaZAkqANfM0DI5S8kNzvZKDoOX4poe2jmXkBKgXZq8K5zvwZmIWYXQ6gtdfH
Iyq6HiWGV4bzU8IUYrhMC8eBA6QV7EVxT2083VydpKDkrAmKpcCYoUxHpEROUDbk
ia5DlFnhntFafPzsKATEr1cFx/UHAmSJQT3nsm5CLNZHvvbvn8savl3cGDTP7Q0k
X3rHPvMhybqOdwIgi+K0fHN5XoxnsxaRzoIPJ2PtcQc138PtMQAdGiYBaVJ54r0W
SkiVPlw4wHq+keQHFkXlhZk9T4SYTr+ymqe/tISzeC0j/X7KP+5wpim/hSDSp/Ag
/FRiYDKO5hBlYGcLTCZVZGcbIy8zsNtVESZd/lLpFGAJDpovl15Z2pPl0LvEsDVY
WtosGjng3tFiq4YUI9Fyptm0NAY1NoHPgzBN2bJ+cZmLSIYXjgky/yW4PmbvLqmu
fomoT5m2IYkxiw2Ybn0+9hfpFF3jvKiJlbDS1yxO6LgLcvHrC0/UQfhMh3+5DuJw
ICUebLuUjz+i2wQx0gRco8E4bGxpairewY6GTqIxRI7DH51deLR8mbLGwswsP1q9
4+f78numP2iV09+bVPrjFvkEdI4SUMjjI/tKPRdZ2E0zPyPWs88PHmy5TrFapkgx
8fLYmsAIX+5SiO52AgKtu/FFMo6A8DOc4kyshfBh6whj+nraGjuqBKHUUdXsoodr
sdyO5zjcfHE2pwZNpJIjOrEC1cOwLUsq6IZs+qTv11U15Ll7Mt0atGN11C+hOaRO
3cB7UzME+34l/q5hHb7wI6L8qMFOIpx7A2qkfqx4yRj0OoQ1wP5sCM/KmwsPqAYR
wpdRH0zOHjPIdqvP0LlhMwDIOPCIrZe/94ZG+vaC5OeKEtDLDRXsjZa7SWFS4VB4
KgtVPvp9Cl6GuShj2oR+kSk3L3IpFSwooF6gP+3h3R0GZifd+VhvlQJ7YY/3OFF8
QtCMdSSaKLhdonm162qltzFKXFhrW5ImwbOuVDDbCPOfnfFGMNfMtVt8RV/Z83uq
S9d9ZFTLxGZRmMqsY5bTZZnAxoo3frWU6xR6xsDfKjx+MFYB+2dnjeFNY/mQJp2C
9akP9aMZApnMFFRTMXJ6EsSOQMgkXD49qlupctY1buczcQwT1QgBbD4rciDp3Tkp
3vy7AvfpKO29bGDCs1kXL/5KHQ6gi8zjauhwHmZ9RMnYYYsy7c+PwZVK+bqPuzGy
XfwjjiQFHJpxjjiukxnRKbICvX7IFmAeeBfk4zHGiMBoR0Y2ypQ/ya7NX6FS4MAa
PJN/eF6vghw3yzaXyyTP2WQGymJNE7WNDFKBdJrHYTAtvzIiSRtmqe9wB6cyfCPV
uvYNa6eLW7JKAzUnpaCXUlk4Ef1sfW2mQJ7a9t9x7KNTviXvcnVF4WC8kC6lR7Ur
hQp5BgXODCBOX63olbxenzxQWE2xqhty7Q7agU9OO/JC5DvmiepXnz+823tKZobU
tKjwHvpk1rF7FswFrOILPTLHSJLy3bowGPKPyyvFGaCLRo6qVv9UrJHq+W20KBL3
/UFhT7CF/wekq3TQWYNNd98diCbTLfanWFFEIV5QpJGs5HvcjOfMarykUvg5ig7/
ryDAf0NEF417bJA5HC/HjFPrQnkyj4dstK+wORI0aDL0M3iyr2sSWoFt5HyDQThq
+RrylMdgCt7Hb+5kfLiwpuxEFm/huC0VMxRtceWd7OnFyipE9bbzNoTSJR6SD/Xa
unLmCilPXgGFSdyXzIKEfOreH2nrV/yu0tQX4P4nOCyJE/YNimpjqW90KfTKAXe2
mnJ5WfM6m3yZp068/ccHNaxGiXY9MBkVVVUeyV29TrT4T9mRtG37jxylyMpwYJp5
BLWqwGJ5DJ70YftH+b4Q869HgXLbIGL9mizERCxD5npErgkgbi3fGeNkbxUWEefS
tBLiGhWPKQpc+oT64zMcYSEVKx7ADU5tCvtYGX0sXgTyzab+VdqDvBDNmSSr+Xo6
+XNuGurSbXXnNsOCkXqod1MAQWdsLbE6+RLxiKWy/nRSTOEO2AjiDr5VQ+5KOhPu
dH/I3swEOPjjEUrdWodLqSwSvLPPMEw6b6zAXhRxEE9gy0zCc71hQC4ayVZa9xWr
N30H+CuMhEhF4+hQcItbnqmWH23y5ZXbH+YKgofMZCryI2au3a9ssKiap8qjypNy
6A23vQiCUePX4I2Kpx4QUUncKb6CoCagk9uw48N6SBSrBTR/+e00Y0CSYIcesyRX
0ysKlrf9dEOIwTXXal0JB2Jgjx5NFoMJEOWGgFhAWzPyISkSCPsZ8VdGm8J2k+Oe
9ZCBZiTpunTJ+g7ofDbZdAp6Y+6XVxD5IPQbP9gp5sJNa/5yzExwYB4WqB7AMHxz
HDHacN6KYwXrP9jymClhKhgsnTNLl5BtFSJpWxXYP3LtdEK0HUKO+++Qc4g3oRAf
HGef8BYnHhw0cAewWZD0qSgN37EKNW/xShZSB7nR6mw=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fUaXMWYecqpb/VscNVkk1+Lmm/Rtdi3EJuYl+JGdIwg4oBZl+zZXndVFy8O5uYTL
PFfS8Cp+/ZWNp02ak/62FkOkzAqqq8ZaKpEGPr+bB6r4vGRFqwOSUuXYCi6X0sl2
69Q4J50c1T5b/eXXopgQeE0rN/PJSP7Z8k1/7x18WKqTOQZIxXrN5HRrq6H34W95
VNcxFCBQqpkalIkvPL9CC90QK8H4MA+8168ka6VrAToNLGMWbWbr3vvjh7s67LEO
d2DVNSb5HTzuSMypwzzbuSbq4qlPt917+ez5PvA++gN55JUhuniRI2w/5pJ93RlV
T8EYmcKLtagW2YWbAqymdVEaz0CeoaA2vkqzZFuKEIOjmyYOLm7LQIxnb5kd0L0I
40BQdH4wQ8YeiPzxKwpP/3xl0d6V+uYSWW2m+u+SkAjNQ5tRnu6+5gIDo0S4z5Zx
1iwlUrLNiiMaCBXiaze7XZTiFUUutEIuPtC20kgrbblSbh9Hwy3cQw1X0dvyHA6s
nZDBHkU1yPMUa+49IVZ6HpfYH9JLO/ngGmUTh6uqgFpKqpmd1ormEGdZzSSAmzRr
qqBY1FLowzvwptYmnWyGpKrIv/qZrZjPbQyHQZ2RyMrIUS7nu3VaZ74NuoCJJnl6
EC7dZ8UCWAU95+BEBKi9LTM06H0VM+sY9Ij/8Inc2eG47ZDmCt3oYkK5mvl3FjCm
v1I941bhb63Xc5tGks23g7OhMrzNuLP0xw3abeKDGkHCFq08BLc5qtxiMy8lGRV6
Ea2tgmVSEyOnYqW0thwJYAhXe9xjxw9455othAN8Z8rWnL94B3pUzaqqrLjI/wKW
L7pwPIVS7BsDfiCCXcRpgf9WvimFfpGxd0RP+fV0UFTdnyZztQFD3VPPSv8fUuUD
yxVOFw4Y3rs3hPCE1Jw0h2Zp1/SXhfHs3ZYMeFee1fpGRS9XrpUN1nDWycH0Bd9d
Jg8OW0u0hRtivV+R7YMxus7NBXd3UuxlMrsUh+50c+zx4pZebVJ4nDtNHunFFEVw
nLcnOJ0zRsSXnVMz1pTk3Nes4pRSNrvp5+Xp+I+1XMM7RtFj9zfpZ5ajQQuDV3d6
bjPmYFmIqfz/SvbCaM4a1DhOdxXly6EezNNBi5SyloRzfR+D6ayiK4zPtEUzCzoI
SsxLGtYQHQnuyGPmqjkph9cjCQXBwCM9deiDKqOTjni8tDhve3/B/Tfy9hDVJpIu
2X/nXv7nQ4eFEjLYawgXqMfGqWirgkREqVNPFCvDiA6r9bDIwtkW7GVpEc5gHAVl
HgdWWkd7A+R5dDUTGmMJKXEe2UgxSOT6oOuLHCETLghrOma5wP+EfdfLXOPzlN/F
HjEQUM4fU+gjeKh9qtPnf/sU2Y+Fd3AkXxX13VnZRTGWq6IQ8HK+PJY/zCPxQvgi
+N5Y3PiBtlp7D8fSzEUIjFiO/2Ks3D2yXgxCYvJCCvX+ry/InMTDiyeWciUwl+is
cn857bGqdfvTNVtIJhAtXke96VJIr5LV7mpXhJExPFmA0ZfxuXdjY4VQhJrefgSa
vlMEqxXDPqReQ6z5G6mbaN98EXUGHuevjFRajpI+PImsjBCzhYDYyDcXTqY6o8Cg
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Go0LTJFfkqEo3vJP79GjOsp4jjlpneuwoxAujBODQEPBUX/+DryhKxrNaiR/b6bV
8+/Hc5bEk6kMCUHe3mL6ItuQGpabm7XyRrZqrAnY3lXOTDmggOQqNiSXDmWthVFw
ORPMCM3uInxFafRWzXTHhFdKKyY8MSJAAHTeERhIJo19IfPIvNYQ6WuUW/Ur1STI
kUyRFtNQ8FD/LI7hOM9dj4yFxHVbEtDx+wuQavlJYiup75DNilEZvhCoeCY1k1Qv
4J6R58sYrE0t2L0sE3fb8FNUMFHqxspCD30rvwbEDfLusyEFi1KwdQeApbtiPkuN
lXCix3LCZZPHkBdCgD9IOHTw3Mi1ZYwVkZO96OyYoDEYQclUOTr9xVipZL+zB9I0
sssONBjXmFfZ3KAs6mF/0hCvqp/+vubreY3UtCnVnY4ZDOIldwov4wTBDhr2HqHz
yJqOTGIlNihMereR3ZFOp0wvsO/EMGcH5EO1zjiUCTQendyUkHIhxCGThEgYCNwk
zZVTFl34LI3zwW5lVdREZ2CDaVHeYNd1vQ+l9HwL4lHVAKYa9zF67MKxzZYNwiel
8fQV6+5/oyrW8RK25nk6pfoun/gUy7LVgNp9GM8zd0eyKfoBkJSVXMoafT0qd352
Y5LCQaQG6yYYpAdhGye9F8rk8CM95Usz1mQBq0rLUgf5Meg2sBHeLNlsVV7ni5yn
A4tTMDRAo+Iwbz3sV6ybpr8W3Z+2EwJzT1V4Uyv20xgRpZAZss0117WBgRKxDIHN
buuazeIiVkB2JirM14VEgOowtWUBcSNDoELF3cstEiM8izqIuxfRSQhvVJGltHkF
6U1vunu+kLliWnPxW6FHfUrZ3urrjUXEa2gkkhRhxynWGIythiK1WfKgoz5gqi1d
DEaIkDYJzfy9iKrNmKaG8paDnUmcuVcLe5CNDcoqmcj43aeiPjwlRz2WG0lS/20p
ouE1ws3aBMNJ+25YEF42Mtc37eu8k+UMufOE+hXebmsVJzNv57xUy+MR+PSIhuvh
0Maob8Fn5BZ+kVm/EAH6etwFjJnpPR3WGKFH/XkroDu12m6QGJAAUJlL9/kho1hH
lQ5Vr6F/N503lEDrlCw01NdLz5oRQwXYLv3+9lbyyBwa7QH9D/GlSCM9WEpBFj+M
X/zI+mQFX4Mvg6y789AZhuFfdc/nDbO116FDkQ/coueUImfHutkQvYHSxo1L6B83
zkpD3ljjXF3mjtTLPtBl5rsVXfCGaNMoseClOkZbsDEUvfLrlEzHSf8smQPmGKJe
lqefOZz2KC0dV7o74eygXkcnMe7Qix8Pts9Pry9EORsuKAIY+XAB0V+TFNtZF+WS
CZLNO0Xs1yif2P7Ye7WcHwx2rAN216mXK+XbUVEcdVQTrPi/+5MRh3OGcLH9szyj
6i0CkRPTyhh4I1URh4gVc3OS6vxjLpi7CextY26VMvqE/Aau8RUPX4IhzCzFhCmv
7C01gWu0+jqNHaN20RGZ9k3JaH6CMnWpMwFiLCNGhLvWk87gMCXaEOQDTdVdoHLQ
JEnl3LJfk9RcPH7vcM2KiADsyjgOaD+mt0ATvmJeAyHjtTGkAr7Td+eRpXxu5jOf
3M5wHImFdOp5lthiBgTqLh2/DSotWZjumnIlU7Lp8b96OAbY9/l7oO69kVUEzIKu
78EaXD7VaokXK7G0UVzf4KWrSsbvNkySlLP8aQ6SNPle5EMDCTeIpJIA2olb/63C
VxVnQ8jhGlQYc0/s50PpSpbJKczDdARYA3h9TEuM6XBiRLfFFhuTZH85G21qn8tV
uIbc7SB05puuS6J7NVkogZDXkejZwXGCzt2VZu783s49gxGohMg50qUescjWO1qy
ogQbMHvQLX6I/nfbSOP3sCRlT6akAyoyRD9CqTbFcxc2voHhXJ6orfKlbdf5jYQ/
e8ue1KrcPRSnFfA2cdFpTB3+a5NlUDj6OPK4/Eobszr3GJSi7o7kV/Go2crhQzEp
QFXBPXAbUV67jMo+1tG50XBTLyz5wN0pShiFhRN0i49UJhFBDCDAbcfiapviwXc1
WIGRWjUVkGVTDlK0Ao6X0AhDBz2gft3VVKg+YsXTmBng6c3DyZ0mFhhNDhfc3RXc
DkrKQmATbGvZfuW7D8m1yC3p/CoPjjGIsSHqF5jaBjfxyU/V07ZPeXXrAdj83vOZ
xZFesq1rrmF7fCnJPn7/d0Bs89Sn8rHt9HbJO7iLUj/PErfL8c0b8wIBzPoOrmTT
ZcpkaOQUIjyfl0mXrKBnqBrp3+VWTQ5/+Tqbrvk8bFFucJJpxJMKiB+lm2Cu9PDK
rho+W3w+WmRhPxPN6Ds9njKLoBFRBi+O6599hraB+Ouacv3utgJI+hH3LD7dpDHn
146T1ETALZKaaovCy/iqikNFE+9SNwzOxCP73+vxj7xYAJnKYwNs4ix7DjKSxiuz
Swjbe5QLGrf5YYvdNreq3Les5aSRjg7/+21j09mUbr0477UvvxYDhrJDN64Cym4L
wkm1ZpiplF6ugXNi3dQhesvbWYKcdnDwWjRol5vw7vZl1I0whxdJokeZPEMGQSE4
qSt77vrBFN9H/hk8hEu98DEADLR+yQedFnx2mg7Ps6/RUH3hKbcL6SwJsAcjT0y8
K8e2d2AKlvlCvtmuJNhVohC+ovdqM4EXXl/ruZ1vdr2UgSgwZkRdzcoE0Omat3vp
xBf6KFyf5a1mIfEgRGil330jsJ4jDWOlax7db4tj9Wds1VFE3pKWRv9m/EP3YdTi
CeZGK/Ea0JdRYE8ryv+PFONCWvbg+dCaB4Pf+sciYRA9VKDkdq430CDtWuj9g2ez
NEuHbD9glv5VdBzE0Pk8c06FLq5unmGEk0XALMagOk6DkNnSyuNKoXGs+EEp+G8E
T9yIF/8NanJxfsJEo+K7Q3VMAHsRk04iSf9HFSiBWpUp/eoCZfzSHmDdo2A2JCII
G7oWs9KcoKXu9fGeeO6/GY34PnDQdzf93pyLIYQKKCnomZms1pct7U0E68muvFTo
OehsRbrU9zFsLCFcVJ50hb/KidJaUHBP++zsbwZ33m6W9BNotyz3kfcN7ZqjcRvE
wzkosvSjvsDVhI8lTOkyQXyNdG8h1nKhgbxpYKyVuyCnWC4jXEXDCE5/a/Er5ECh
VVgBUPLLQDDC3wAkrf2NNU3biscbwsOX53opr6nnml/BKrniYO6/FJaVHe1SUMF9
McS8Fsp4jPcd/TwWjIyf3OiEaQDIKDdOrjxkrKeiFmVnz3AHX2dNeoD/TeonRxcz
Ldl6Py+Tg6tGVfjbOM5DOO/HrMvcxLXtRMxTDKJWaCr+KxJzLj61/F0IqNbo+zbJ
IFWXkrraaWnx938oEtGkUov+GqvbjLyB56p/k2E0GK9Iz0LfD2EnjzXlBqZqNd9V
A8UAMnyAEP08L+/n6xfgSkDCLePfXFnuzDipvD4lOCbp/XRCsHeuj4YbsndltkfQ
SDGDpT3j4KkpDrp8vfYvl788NQ6Uz99yk97s8x31psp26chllAAyIkLn4cZMXSMm
OojCS6ZHuqmDK7HLftGcYfymEEqEA9ZAIiAW8p9kjNIH1IR69wTo2t5V0npI9G9v
JeQB7kRT8ZMfLOeaNC0QQ/TBFx2+qA5VR5thWF1gy17pxoi2T1kcqsoVS0pCCxbp
VHD4PWXubQWMZFXD+tuj0kqxU8VJvWatY2UzLz+IKsSp2BWQn6hgfQ5RD7/crAh0
jpA6Bj6dOcMwPR9m6suPy8kncTP2VTFbtFr3pfLrOZovTcj0tcSZ4Efj83bnKw0G
gTL10Q/8uF2KEiX55nL7kSuuw9w5pycJt48l15OpMFDzJqskKhVF4CZHdiWSYBEA
ESljMW4DDRXticjMngfzgcQqq4ZKGuWvSs0Ko+98xouyZQk6+ZB7OJ6yCo+sRhMz
Mn8u5E+sm0Qqe1ol6UUtOZpmEVsrYmk7NDTIIFsVSW0HAiKYGLDlW8+j2+RPzcUz
ZT92/Lwvowa5TDnp5MIXMg4PXJ/qqi8ogf38Pk0s5mfiyaNCQmqRAyNKnrrimEjh
HcwJY8bbM2vVVn82LNg4NKYzWBAt5/Fr9+kJk/5ltL2g+g/WfYxIIHhwsVGMPtph
uK8BTr4OmxAbLKNx07e9aQLCuNYaIBqDEKPPdjvi3LbmOCtdEIF49Z5CT032KXND
j81n1qsfVmkDuly6On2dt16dV2Tj62++5klxZmuH9NCuUpvGG1bDuMu+netjUpEn
Pjvf8+5WFlNuRH8Am47j7S3rn5Gq+O+hCNV2v8WptsHbRlszf6EcKfTAgrogdSiC
0ux4bMCwFQEJTneBZEMsfZojgxbJGviJZMt+flZsHENp6tyuM9ywTUMemorl8HGz
xP6kgXKQ2ByQ6YcBetpfxe/QLT+6fuqHrAUP/HSh+79a9pHUPvMpcYJZIH57NAFW
CFzUP4clTUC3W/eSih6UW0IU+20332m+29uW14aVFlzIwLIpleGuJOXqt1slydbd
yYgecOoUYUyyngM4j5BYRyPepiY/Xh6KAIyn7mjcR/ODS2z5VMeiq1g1mwDynbLn
eTcab60gByLPBnH2LRCSOPIO9GiiUgDCUyO9Qu+QjEz6ecSEmxwRlBZF/pzdTx/m
G4hFP4Pp9hKz00Ic+Wv0EX1KZzXPTHRmCxKZ6/m/OmP/T7HqnnuAokzseXqsqwyI
RZ3yN5YiKWVi9dKUXwsIJfyy2UOy0uVxqqxpRi2MC2efOGuO7ob7iBZR0V6fu1bU
1y21zvHxF9nS/DKot2NGWZ95/Cwcya0l79tIsMo5lUaVTU1J975BqI1u8oHyK2TC
tGMJ4K8bvqlcPA2nYguDoodP3LBNgzYFpAUPvfR0Y6Rhdl6paNOG2hA6fWlNq+Jf
3vCXGbn/yoNRiaFvCFOdGRqPm9I849Hxh4NBxrTO4C6UCfDw6km6lWg8tJBy4KTe
29etDp/VAau4K8ntdvvSgcchfsgyI+kRMR9yFkqI01ChImacVhMwSc+j244yKoQP
8YjwoZOC9Og9guhkOL/gzEYTJBBEXtLJKRpsp0mlKsUN0DFBgSIHajeoGl4WSUnY
9Ri/t+rj/uQ8iKwykbSoRRSOVY5/aptDCa8b8oCZbta6jeBEvOJf46mFcJP8UuC9
8JCzbqP8PoFf+0VV0fmA8b/PWjh1+PvKjbT2CaDE7kai+mBEsHX6uWK2etJu+sar
7JjHsqRdpvmKePd3uEXTyIvnfRmRCjM7dzD0naV+zMXgzbVlad9GNWvD0n34JELI
Z5HxX0lAWuJJ9tx6TT3QqlgcibRcp4fyaw6/76lQ6RezP9r4IC4zxjkCUSCWY2wA
cphPQVVcvD4nILnd6LoDxz1InroFjNjZ41Dgi+kjino198or2YsOI+gGLF0ls4Zh
YJgjG4qwRzep66z0R3Sh5iK7WUcurGX/5tmrIsw5KoEq5xsf40IAZ+YYeE9jwaiB
UT7UggLeWUMVYyt4JgesWU6YY0y6p6DaqFvRNtzRFBf79ygDxCiC+AaUKq7SxhUs
sHfOSRV0MIYcVfFP+dwmAC5yfTOPi10dXZ6C24bJoiFpL4bWDxepNXgxpiQC4FH3
HF9rHJSX3JLvBrGmea9sD3z3m1/LCkWYHL1Je1Ir52mQsq7yw9RwtnfWK6+3UIPc
kTdQlB0Vlq5/8Tei3dx2wmbRgZWpWA+6igriSSaKA8DMgxL59h0nkPtZsWf3ouKA
hvO1Br8C+6/uy3aWTNhYYqcMT8XUavkAFf4E5or1dDUzBBVwmGcQaA67irjA/Cqi
LNit64IyZ0fSh2vd5209fGGN/AV5hICClV6jfndtFbXmAEkw/JALrmh9cV34VZzN
mfpUigUERX8cgigtNVKRB5WfNysnJ9tZnJg+BZqYNHGKmM+u2ZR6IctlQD5jdXgB
dHCwoB1OuMc/p/dLHzS08aSw1hAdDS6rMAp/s76H9MSshFfGaqWaoWL9MllF8upV
siGyWMyl8Px1d2OfDNGAI4ppKFLcAYqTvcFbtf7SEfhJbeE0kyd2VRfo1DzS75FE
cH0J8LnMCV6dP0hTWeoLldrosrqAjypo1TSHf5tnNWO6A326vx7LWxo81eck9Hdi
EitJcstLVFNaxNae9mBzbEZL5+gfBC97Bykv6i6u1RnQpqKxENj3P7AuoMI2P8bl
GniaL5zUAGWe76SXg/+e5gXQXemaC4pPOdXaQ83mxbej2IwlujCA+/7/S+4JyJXQ
txMj4eJDyvJuozyMwzZj0yBW9/gZjFoBNP+bbpScvjK1mVtMrfNp6/1TKNf08RT8
9wMNRWPfct9Ogd8hscHoA+j0nWpIhA5Jm8+h7anJ/Hy1g9PuG0EBI7P+TcNnvaa2
E1RojxSpnYCRZAWoWSJ/lfg1wb+IYUcat4MIuZWQGHZykWjrLUZ+8k4h2/sXind1
Jki5j1yEPwoGy84cg5Fwxin4mkUxdgT77XvDiYekJhogvipe8GsxYvlkd0U8rJH8
k+CgG+RDD7SZE2OppOzBupoZc55aBKj0QJWMyXM2HWmTN9fB85D8WMm42S4XNz5o
WU7gpwjUH+z4BMFfSaYzRKOzfjoQ1MUEvkhaRPbPTI0BUd6f5hhoDEFvlj6sxQrZ
E62RO4rsXIcnIVilla7qgepUzLSS2fst4buwOzE8d0Zw7LWF9S+JcMmT6+hBmFK+
fSsbNCEaz04/F9VPIvSzSgmZf0RPTN6Ipopm/wOiA5OmzjISnFlYJ5oNwhKLUswY
cjwp5zn7g/sDFq+snSG0JGyT/7qn67OVh8rzlp7GAyLtr6Rr6x5n1h79fP6iXrl6
FvBqiMD3TG8KF/oxHUOg0nPxUAjGgz+fWEJwv50hnmv6ls3BGf8jbi9Rl1tghUAH
F0TlqvaADHck2+EpQkdV6CEjOqvI8Mahtqd4N+NU02cVgNSTehTFivp5eVRxQ34v
PP5b6elNCiPnVe8Mn/XTyWs5FWP/0oyZf392um6si375KmIz/Bs1A8PEaXs/R1M4
er1ENlimkyX8af2iDNdOfw5FY/XXZJiSTWKVfENm5o6q/9mZQ83zgiEhU8C1o/FO
mBODcrKaKJ4C3LJ1xw4DDi9BSemaJYiu+HORTZ6an7ibjmiVOEOH9eTVpRtSXysY
kLBEa7jKStd0W8zZdJ5POqbjOzy1KtLuDL/h3uMyNGwMt+Jx22Lmxkc2hziGk2wG
TLqDNXagcW5yjzoKoe6En1Hx3Oi7xMEvbRTLOZhn10S2mGObKZT4DvzSyLx7AhHh
2i4eKQu237UmihHFR4chqCuwh0ECHi4uvYLayfNbGQh/d1tfnnxQDaDz8L0RV9V2
bKBOcQyCJp9tXeZ31dj+MmsMQlXyc7wyH/5L13c0DdlHvSKcXnHSfxnydUe9iyh6
zV86vZtMKZ4v/o7JBJjxbgo/vKTsA0cQDuTaYawi92z137VFDiF/+SyhHcIw5rwb
5E3xq8cSpTv3zGc1FlJ0aDJZXxWB6ae8yFb/Xv6rGex8GHMUBazt4MAojXKaFSng
ciyQvbBWG9f3rpOuXCxwvLTSQC4BMe17yCdEDbEhGG1nzAs4txxuNRhMjQRo2+4+
o0okVoST7McBjp5TR6R7HWM805jiFqxsTvm/FkRpiV0BzmY09Rn0zd+NBGjXOCuc
w0NUMTJacplqBOLIwtGOhC0WKekRiNAQ8E9olTowEgfYy2LkGGtGWOslL4LnOcwy
HcRCV77mpvgmJn/rel0XQBVTRug2Y/idcp7ktNkZFNpNj6Ch49jIleMt7df+idsB
efd5KrVo0guk97RRQriUbELtQBHfLMh2lWhrCceiz3E=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdEPfIwANudUflXTimIZ+UH0oVs5uGjD0lKQCGuDQqFt/LticEfQzYMvy18uMRVj
QM5AOebqujfPJrO/gmkSkvWdonRcoR3CT6ZdYEhEFdup2JBFohDkuc1onb7M9VeN
4OdqjB3QCojOn8QIDTTLs1wbNnbTTUXj4R343l533Uh0ebp/gQeoMm5DK0LetNC7
lGkDO5Jek9Q4JkUgbj4oa3RqOHsQJI1JqfwCVOt/9rW1vUnEKRncchIGlYCz2y8r
xlDKWlwgI4ONK+cv3OpFy3KlbgZmgyWyeRPHMevdOYFpk4+QC1n61ubwrBlPVjMc
u70KgMtW7P5XeaB75JlGgm8UN93aMtcMsE9lNNxWXXTxS13ZgAKwyiWZE8HBiFBH
3++8YFlwKdvj6GenVMFKdwN00OhAuwBwD9L5SIlWCE1RSAJfWhK5FmuvGnLKR9i9
IsFBjQbgWu0EqDTVbgqO9hganWVxkkiiyMnobk5gDLgOEQAbtYE16PWSSmY1WtUf
gelkzWIK7MjyRFjwshuwSSoEAC09i5pCqynffNZ4h3SW8ncpCJ4cunTnRwCqli7y
yyh1Is+Uodn+K9BoW9GKH/RN2raGGgvHIKq92zvCt9224I4h39Ic64T8OsMu5j04
lVYs8zLS3Y2mh7zRD1cScH4DpHcqDiQsCXqB+Do1dBjRYpAfJre+pGkGGjdDqC7M
C7/BJbnpMl6ffJCGvGVlH1dpWwWNPRNgGdc0RickvPuubjcxMz1O9xn6TScd8xHV
qC8RamSiC//c5zQ10FBdsjS1/ODTYpMEQTV9eFo2xcnz2xioehNBw6/MOt7WSSAg
jpRPU8bvAGKrLV0R6zYECygUpKO7zl7C3G2NU4cXY6GpcwIOKh4tZ5ssYPdTWGRs
73GnGvXTzZRKDNVLk6ZkzZf+YQqn102Dj0cw/KW+FnMstt7Uopt8waNKn6x6pFA4
FKopFvdLcwgr6vo4YPnPxBzNw/yQfMAvezeqyj51Zl+ID2HVuvzu1bx9gaCaMmZg
C5td828YwX4bD6NsHHchHkBHTlV85qoRgZbrztACGM1rWu4eGsjAAM0/59IVx97Y
hdt2XXiZXx1uJtzw/u6mm3Q2sdyYuoqTOOuILCAwe2rXARujtuwA20dVWibx0JeJ
6dQ57wG/pMQaCCwkaYr2FeQnfb0fY5y5puIxCoktTZErBTURk/K3Z+3pCi18/CAr
pMByiUiLxok9kYAlz/nERAhZ3caRXVsNVGBe1xQdMvXcmqq9MDCj6VzbpBGa89NS
urfPszcxJFDPBX/ePaMACh11L+fbwV15BthC84rKPwgD0fInjp8mOy0f89o4hU7Z
+LQdpScciUXw5gqefLQcgNT58/ee54gQ0N4NRDdFNUM8TlJcqlQ4Bf3cdQbG/ndr
xGWJNwMorAJryPahot6rrFl7lHaQrIeCHXi7pbaslfPlWXYOdBDZ10ST2MMbqANz
lwaB2aUC89AccFDroK9upQMqyTYXu5t0HLrJqJvFaNZz9B+Fplip0E3Rsun4rOwf
QTS9P3fRFaEaQ4BOnzzlaHWc6uqV/aH4HcqnhXabp3eLFrOT2DRu2FbcvXhCVTFm
dM8eSBVmxC0XoKWY1rmzZvVPM8k8hnh+L8XmEHp0mhCzRc7i6rot2/OGrgvx+QNE
VNUGkgpUaYtoFerxxaVZVQ==
`protect END_PROTECTED

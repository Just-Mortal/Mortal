`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5RT34k5r8a5HujMY7GPocHj3lzd8LZ5Ae8JLdJ1ICsTdHn0KBZr4wGOyAWJ7S8/Y
bU5vpM9cwjoO8Oa+J2VKORajIrIN+gbJw2rMiFyerDv3OMx9+JDNz6i6EPVntSZJ
gVR67gjGVM2Q0gR/P/8kbg3//1SBzC9qByvkJTYQ91H2/FvbqZmWiwgWLQwNTr0F
Fq4oOOZIAf2VvUe7V1cbqf9gPjsO9Tls+TsLyu0Gq0qvV7bVwcxRXkxJU1HSNhLW
M5XpUwGXHctECWklWNzIyajMvbppJH6NOy+MpskRaMHzZejlJoiOcqXnSC+PzcnL
fkDmsz/e8E1LMT4TPyP10e4RI0JhnYLA8JdnVgxaWd+cKcNAne/o3FI7truIpY2O
RxAB3ysauSZMZAKTZf2lAmHaJoJaFWESt2xH19XKRNVML7qv+usUChIkvC0ZQ8ES
Me3YB0eoAmjwT1nEdtwKyr8BNwFo/DO9xsK3SFM4Jxo=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GIMl9UvkkkzCNHzaT4fr9ybif2B2XNEXGf5lhSEOvcS/FyDeUJUzZ/8f6Kjj/iO
unqinhmdt5H27DdmJalV5WSK6mWAxNPGfb0Jx1haZwfTzdh8pS5z6L/e2XLunQwu
wujYA5+hrcNb/Dn3pnDt0aojSCi+h/t0CnG9F9axQwI42ToaOz46m7EhWfFLC/OR
Jezpe2OCf0RogTB99ODTe3vS8iWcMMBQbXfdpPrGfXkac5qqL4njgegV9joN4Bas
SZ5faTkOgOnIYIlIZSlIy2K9Rlxf5916FH0Oh/KLfoV8bZHVgVKWoRUJoAX00zRA
piSV3F7h6XBnK7JDYEDND+LIRLaZi3r+rxnCox0F/dl9hHKZiyKoABOnOyCHlCf3
TeowmY7TQaL5doRXYs5XjYCse22f70Z5b5eq8tY319lZzkUJINTQPXqKChVQOzfr
MBEQFeULkF9E7HhvKjYG3yYWLl130bgLXFCxEkozZZRTyXjlApMepjpKmBhzJUw2
5Mswus8G4P7wgHuRiJcGzqYT7n8li+KCsCv3lm8jAD8zzkZUmFggh+VqwW/1reCp
X+2SiNjaoNHrQMzHtKmw9Dl5zURoCBCXyZJquHEeYQ7RaMW7tsBu9FB1zfD2TirP
+8qcxZzanMtvjFPx+SKrT+LAHaEUkab2o3OhJvwRlg/KcCHpkyeMJQv8mDPbQ/k3
ST6/uYjjTqsprTX0ch+bfHifFbfkwhatoFOfjbmpdFX8tmhavfzZm7IG8ZEaHYMd
taK2N0q5J4f6wz/lYar7LarOpXgKMLtrHiRKN+FDcQHLFvkrdvRp/fdWyiq232Tm
raxsaoKf8cT3Gn7Yi2W2dhEm5R0lQ1M+vg34VW2kU6fS+fcA3uJXQR3UbIfOBQIC
7H1ze228zm+iRzGhA/bWqY7XSCtqvcGA66MEejHfgxm4MlgnR3x5LvtlMYCg77nU
vj/B+VCW2VSlaHihq6xlXDuy7vqeUiPq85bFwA/miltCrBrPmC82ejL0yUoCH1Hk
/U0MoY5egl/u2CqFRrfKN1f5/G8FEWOwRYfuDG4ubOXTirURxvbaDEjdG9RDY1WZ
vZzOo9Vu/hDLWzCMCVEGvw==
`protect END_PROTECTED

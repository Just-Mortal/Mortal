`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
os0UClfObf5NDWG3E5es0SM65tTgUp/ptTlsSOFo3sRL5lY/Ak9VsCXzOctmtsY6
9Ys7hK+BNHDBOu9WrAz0xucGgX/WpaZfjCurX3wBqV5KnrQyfgsiuBJNU3PEiyKM
Nj7Pbb4WsRTKheKOvqB5p/wDBxnb7XywwhRK2gYlicL3pZH2rroKMOmRz+iG4xmw
4PYsecNbnfPv9BEXxLP0NNb9r6E908sT9nyExqkz27Pdutri0bSj5cNAX3uN+Pp+
ANcKgjZ8sY+CKhJcXkN77CcbUNUXC98j33k9jYKmOQWISkG7fDWFUCvUr4EwlgnV
XZrZyVamOyluAMvn4+mImgOgpwpiSEcIfheFMDXhArdW5lJivmvRWDuXreQQhY1Q
mIdS3uYQscRITHZ3okJSgUMz1vkJqgH9K1+SS39aNdj6MUj6u0d3lCfeTVF+GRA6
xvmQU10XGrERdAzMKcEJrzsSjpl74giZ0sdScxC5PKeTaKnPTUHUNIQBXznoX9lP
eea9F3fkS9GA4slDj+SlG4Tx9oo9p0h8WhA+NSWUnVRML+ZiV4qRdzBgzpjQB/NR
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
40eO8k1u+Z82K3pUUt4SF5GwjRLmLmnWbpLkQjeMQXmKFMrObgav20AtDz3fqoug
qdNVyT4UPx3FmrjsZ33NK1UcII9/PPUaV2n8myL/1YeguM8qhafiOyNijEfOKE84
hp14oHcxoD2AMHiRSfMN+tAbCnk6hPsTDG/IXTHuUAsQA1Fcn/KAxloU0Dpgajcm
N9Hqp/KfuLemUbodSy6yQEn/prZKp8fA/LoEkvEWzQMyzpF8lQ+8K9VKZM3uqXlm
npmZb167m0MzzyOF7+krPI4uxy/uQcgRDieJb6Cc+b2cFpqARmiCaHZ4t0++BTCl
W9kpUtQCF4skZhY1tVn8RrxCNCAHvnYHBpX8g+NBC2JWbOdW+eomM6WT578AJYdA
th6HLX2eQxMUU5SMQaQYpwELwPMxMkPAIxKtPewTEsCxyaw/g/GJrxlcnRBAm13W
wQrwOClnpbnfI7RMUqV759minFJNl6AoomzwWg2KGRnyG4klXf+tJe03dMBxEdpP
7kRFelGn250/StNF9yiklE9BKaEob25fVClfeT0auISo3RfvwUUWi7SC2ycUGu8Z
GrfOu1WCAlpFliPiAerS3Wpj4DU08rj7E+c/t+gNoHnlwpkgvpa0pzddRIYgkDD1
X4nIyaRO/J/j7rOlUMSxlUHlP/7eBf8XJedg/piPLnFZwhOFByxui/J7Zb1+dDbp
DFvHqcOsmIRvMAVYQTW56O/VuooKV+a8BijLs1MuRpUoPlhxEPhw5sWFFhX0tw1F
dtbpfoUR8XzeUwHQGwSgW0dj4yGXJcc61k8DqASFV87ptn3WuK/zz4gQiZWtQWO2
5zDt/7TFviKjcHH5Bj8JhaHaF+x8ayb4ZCc4I0T2SenrHqEMAb5+w8Yvo4TYVAuc
+uWGzCMy5nSaWd/0CzxryZS158bUWr31tjh1Wag5XXUQscUbA+qTrg8sHqmHL2ZN
/kDSYfhErLlcjUY8m7evjV+o+7b/TdLxByxdJ/iZx9uxUYQu5gq0NyPRPjAcRoRy
HoVA9oZeDF/x1amFVrGUUZK3lBZ5gykicJU26geJICiC+ZGzflJDMK5VG+wDMB6X
aXqG0eGyc1a040sMIz26i5vwxfjBZPLf2Meu0rcOHuN0zXdm7a/qb0CxCdAJ5Fn3
bSAYjynjuWxF9CuUnAniJw==
`protect END_PROTECTED

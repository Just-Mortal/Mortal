`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZQaAGHh7KXo3S0MHwFQoIQ1QsemFN13ZoiFl2N2/kEB/We/vtP3MLp2eHy8Id6/
GJlW8b2wmtgqklI6UqNCVjVDOhx5u1CGVF9rt+OQjOksILsaxICVHfKZpK65ZVnu
ih1wu9EXHS9O8HyTJ+IPWNsAdpxVW0PYHOmgBFm1DD3Vrzw0tEuUNwtWU9XyK9vo
piOoUbH7RTYxcdFNd9X6KzVWBl9VbI0SZbAlY5UI49NZrtA8h3LSx/Da0QSSPIwy
rL2knhfA7eBWnKXEaduFucJRT5LD2BWZW+YgZEbH0rYoNbdXnfMufsufSK8/4VYs
J1Hzl/3B0TTx/ZAaK0TQp07H4HLsiRGcxfIPm5TQ1Bt7eLdK7AexeTsmfIuy4EhF
4khIg/30npRNvSWfjW5H5VCAgy0cYH3NCBG2h0UC9jq3TiWniF6XzhTCyoUDhXVe
SpkW3vonLtnxKdyBZNDrFJV1y+qpft67x95JqXIFdDvYgLaeak1MKahQ8RcTBlXi
O1qvYG8c/PO4dYd3F4BG+Aa2UmC7a61Zm+4A/mPn4CGFHFLpohZj3ZtAnDEgyZ2A
kOErpvGUUOLCV7qid4tb0LwEMqC/Z2me5z6/0gxKvjurzrW8o4HAcMvZ5EXrYSDm
05jZrsm0EUqv+VFgawhHDUDr6eL7OuxsRRADSWQky34ztkRDUQDJYWLsUGXlEpxL
0g8WKR13SIfxN5oRG9MS8hpPrfVWA4N3GaKyb6oeJ74bByXK2PVkwHkRQoN1hXSv
XOH9pnIk617504mrbhUJjAXG7nR2DgnFUizgsLhaHW//nVCfAdWJAsY5xKSCPMT6
3Fr3lq18n8inyI6qXJmX70dwQPYkmLMQmjD1/B/k+3ID4huJKXTmxWDQ3NHYc2Mt
g7Mhy8KVNiw8Vc/H5qqm/HhRfQgZwE9u+vyPX/KAzvm0VuAatwj9Kq9j606uIhHj
xTdOlPExsiMJw4UP/fQrQFqftsJ9HLV+7Gz3pKvbHjqbtAz6luT4FLEquZy4eo2E
Yx0YBfzmXlif0S+1+I936mJqUCovA2c6/oxSKam/PlS9TXiPWoW+N7okdAJgoIIV
LzB6++qBsWtE5TOfGquQVMUiZk7tmm+fX/C0yyMl7A3QkPO4ps1JPxRtwEnubVvr
vqBYNzg2ZR4AFmyunqJPXgd+ejBWcoeFWDVGqlt1vcmhp27FPpKUcUbdr1fx8Bil
PCVhmr2rkOmfP0inVExCEnDAUouryU4nci4y6nNUGlghIkP1OI3JqtHhpa19rVy8
vwB3uYU/S8kxYPe6hmeUIIlnfsexn0DMMVOXXcbQrOxg2TusypsVdhurDEXBPSK4
ZWqJq0GltbTiyI4UvReVi0tEj+o475t+r8qpFAAKc9FIGfYb0k+MvxpdWh8Z2CT+
fL2ZKCYH3OFgnl2lQMZBo5UP5Odv0dUq7xDxyqRCT42vav8CJHwQZN8oQ7SMtUI/
vYWK9VqU/rqwCHp65EezckpYMEpZ9tYNftM5wYKuhOWGBXy0TPmigUMKV5l/OKi7
+HVDL4I5Iz+ncj6QY1McSA==
`protect END_PROTECTED

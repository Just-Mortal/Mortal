`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
32YQAbqXoIoxp1Po+no+QaKuwUx9gRR8a7ApriqEGP+InGuWavSCQNUkVFQE4i/q
tGuDQOwCb6nqg7bQkXaSmDpe/fficcgrpQ6l43x+6NeHL6glf2ipzWei+GQ4odxc
jOyWf1uHUM6qJhckDLqa+VW6tj+oyjqCjN6YXRh6x+NX3lFaUfiAZZNvpJZsP/EM
7smHMtFiQOWvLsF8PHv/TQiGGLZbGMZWTkcWwTNgz1c9V4CRS59lWA9cKmfMMKVB
6e6zmzTeGjlIdkEO8fD1x+XGrtkV0lnBQiUPFa/xwDGcRvBP1Jt7KijcUpKa947N
Id0zZOYRruy22Gk0pQ+I4QNFEy1mETKHjA96mwUEHbtKkQ4PXkOlG/OXtS6BWtii
ZaCMfL2kWMw1f2tm5HKDkR00UvMxh6I11RtFcL5wvJwk2I9+UtNo6d4A1EEGKPC+
gs1o8eVKx7xO+ohdMENmkTeBp53RbAPz9PRaTAA3DB654ddTUIqHf0tqrFZIKQ0B
Hi88HcOtuVa002ZXiyrXKAevrK6gSzRiKAoWbRhdKRghoOINTJCvRip+SJshQ2og
f6M07nJg06dxJp7q/GlluJE++mNFoWFeRSG3+kzh7Q2Niq1rYsIlLoBIBZ9pOMyq
ZuYj8Rj3HpbQWa8miuFtqQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAXH3FZk/NAPZT0+5g/Ws+bBp8qJ53pYtCXDmqIBE4CWPJvKHdRes4A49XhHtFGE
zU957AP3aVrZFjIhk0KhkJmk1JzA9CMrmPg0JicHrdPVEDQSgqfSUPt+kreyhcYn
mjU+P9b3m6Dm5Oybl0JvDiQPYg6XAE3qh9gvObUUd7Q5VJYxoWePksftQE5MEICE
9Jr61sKmNpZQOABGXiVg8ABvyygIMrZie30FYk3t8EFVO9v5GX+2xZACX/JIDQE6
b2DR01UlQVGf531cbLyk4ig0fK434qNoSJZAcw6DFr3BgqCps1GEhKMtJojcoaZl
LwBuT543F+bZxeXO88B6RuUtEs6q1ZUwJoqdMBJ4AOKSvQuCXfx/oqpJwHixtkwg
03eQ/RnTxxT6JF76b4g0p12nLFL7we/+6KJz8ET+uWhzu9BLY6Y6BaJKQi1AQOoB
wzsYeAMooMd/qrLCQhAbXzL5SlX6F7ORVnMM3hP3WPIVydXyP/vsz4WzZSc/KYsy
852AiluqamYB36tbF1pxm8u0gfgKGmAnFkhDlauszkD7Xt8P0OyWiXbueno39R3W
ZvvBr1S4X0JdfslkL+41cg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GMCnH2h3l+k3hpFcbAJyJcs+RRoHybhtKQWD45W0FgZjDVmvxryY8RNIBmnPfWwQ
Gojbw9k1GB/xxcVU31Y85KCOGEc7FB/YacWpn8KlguvWkc0Bk33FDEZwQyk47o3j
1c3+9bwOwILHicAd9OMgL3mzb0nLEXcChg68GVcQIZ1w6qn3dZ0KUVOwDXI455i4
nh8uqx7UohmCKl0GY2onSn9oEEMRhBDv424klJFFBY2a0EidR+1fJDABcC9B/Ult
jNhIsYOBlXyRM1aUeoN1DpOdPgQyeKOFsWljiULTfMjHeo2WEuEUt3GlpggDSv9I
WVjga8+TcNApNHQ83GrLRvjsnFEVOxfuDjsnc5Ilp+GIi0qBdv76vhy4DgMs49Hm
xTRCIIf5rYZRehzohVnpyn7glsCBv5kJ8S9VyhPHMyu5Fbbq4UDQyQLihPKquEBU
CCDoJ9N/RbDt4qP/x8ftYvqs3bTyJM6pX52GBZUHa+4uQbW9dB8eiIwLEn+v66wU
cD7haBR+wLYm7uUsNX5gcpCh+Es9XXtiyt9UUAqwKA8iWNKzK04R3ZWvVlBjLrZB
EWaraBd0n09wDilePv40rzJC2rAI30x8uRjx0AvO3Z1InYhCZtlFalGQ7ldSc2Wb
oWYBPLL7OGfCiVgTdyyTB0PhGXx8yUWOzO+i+8/YHcRaHj+2pNUtkfjGmEFKfmgZ
lA4UzGq9ltMNvBgAU2s8mEza3eF6kOGk03S5rLr22lHgKGIBryhHPDYTStCAv1s9
YjiqapK0FeuXMUh6xiALnhGPJhI8NT25oknSc+amP5l87/7fXoKeSgml2ScSpyfC
uVTp6gEADRP/y62AHJoXpojee7LVIxktqcvXO0k+dj3D81KBM6UPOxpVjY+YEzen
AUotPCKnZAk/CDPOL36iNMLCNdYJckbJWK3SsD2GJxC3eBZUGBK0A5O2kcRX7qU7
GLtWg6NCNsFjlQYwQ7n4eo/Zvm/Pjk81ODKP90LPXZx6YrdBees4FYH3USvs6uVJ
CYawHXPHDhpibI91sW+N9K0rxRtBll2ejmrUaK2PTBbSJYyRX1xngDZTybqTZ6MC
7EBOP/hKNfvxcnQ2kO6t3ZzUpsoEZnhxwnoZSRYg9tWS+0v3fX5MY7kS5ID1LGfd
jqnxU/GQfpjmMTjhQaZ9XmVUNO0DOf5jg8fYbTq3ISWgkgN0XVSYGmQ50k6KPvK0
bT+EWekAtjgr+yd03yKCAGLeJx7vTRBqywBFKJVFu3b4FKQ44yq78y9fPo2W+DJl
oG6KCB0yLc38QFjdjGN2ExIZ9+HC/pwXzmfnQrKhGmr209tnxvOqTxtf+R3Nm3Ca
iPfQBgRXzmdqNtZEYzqxHbNhicdCjbbcT+sXVCzEiX+5rpxekwFe4qfODU/rM5E4
XBmtAQCtECfT5S9SM2v/eYdG7zzpe6yPYM8oaCpoY/IlgRNXGoVixTSLKY8BC7v0
nlTyShqRJJqxszg35ZEgI8GlbTtd8uFLr1qum3Mdj7dpy2+9Vq7xdFgQ04WtQwHE
tXFDj9e9KJeaJy55nQdsxrUtlNzsHY29sSy+aGb9uHTZCcqzRPXZGnAT+6Yk85LV
VVWApWjI+QruL8SX4r6X4p0l71G/xwyx3LCwYtD4STx2tIoz4kQdXtl9KIvD422b
WqPv/4ocLY7L+99n3J4QprSbkQHAhD9NynVpOrNA1dv6dMRpHWsYdmG/DYP0sQ7N
Hg0YN/fNqm0dNRcfnGfER7Llk/DElvlmw9lyr9ln5DRtwZkfqU2GdnNRITMAW7m+
I813vMhtkvudecPabioNLIwrgOJY4BCv+m7Xu3r/gg2Nz/r3oZ0KOA57HeU6ATh2
uai7vptJgA7phWsKn+dWimnFiQEXr4uKBv5MR1fJ3F4gMWUwNJ9QdGBBmmtiPoVa
mvvDcuQf/Rf9TihzMMb9XzBgPaX4raMeq+4ddGpiM7j5Jyinf7w4LFMZT3gSxNQx
p+r6l5S6MzwfjGRUalo8fOOXF6OlLd0O37BZdXyC/Bn0VvjFzU3P6goP/Peg5vu6
00SpI3uQT5EZF45dzDsiUUEZqvbz4/8yavgjNWkdl2oQOs5cEED7cx6qpgJgBqx9
UUnFksjKOSv/kTmq8hi731eO6x+DCXIpds0uUGZakCIdfVb7rPYEBH1Q8LPmDgQX
6hYgm17ZxEjP3MTBHW1JHOOuiPOuNJ5fUvfR/zGPYT06FUPc4p7oc06Ux4D4qq9n
ujz+W8C3tGZNERg6yYMR/LGzDk9DpfpjiCxLqpw7/kv6Yp27YIHDr1NOQpDtl67H
wYLFKHbizlrKBRWtylJkEwkFMCETB98zYQmUDynoBDD6Qt8OlbSPEQGPA2+aTN87
66frSKZJirG2OA7cRbiHH4m7ClOXhozR9qUc7fGvbKBMUpUO5+cfnNX/JyHbJeqM
6nLvO1HNi2WD6swBEEA73ahKapzpgO5qySr2fu7ETphur+Yewd1mC5w3klpv4lda
RuLDsHEAdKi0PECKj8AQJl0y/Z3fmJo2xnvlngc0S/qvak/7PrVdLNyET+tr9jJk
/WqJXo2CFT8LVduMaj4CeXSKthtuelp2WgeGIM8YRc76BL9lXvkME0Y3I46LRqZq
CNFzuo15gL2xgFfl+4hFyN4ZgbYTpKlwzz5wvkvnC1lHm4YQ4R9w4p6blBp0tuKX
bNhhDBhjU6Wnde09OG33c2jk5BJ8WySBi6fq3gXRIclz16sLjuXNnAxMWfnUDmv2
EtKHaDbRe/1OB+FqRB7S2QkeIxgQ4x3gYLicDjp7ULRN/TGWQBp325Yz+AENbs5O
kzLeeLzpl/1PeZUZm75Y7BJH/nwRJw74vEPTAhesLR4F0ScRP+d3qPa+R3I4Alf5
hDfrgTlKf1vBzn1QEkdSRcaeXANnk0F3Yiy0E0KXeRQf7RRi1f7HiEfuvHVL2rCB
1lpGBGy+XWgtoZM9apjrmw==
`protect END_PROTECTED

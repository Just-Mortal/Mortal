`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
igD4z35fk+sn3xaWmPqygB1ui16Dq/sswXWI1ChD9v9IOLbmUDgdjf02ZqYYmz7s
UtOVLE1LQuJplH6ED5n2/DCP3ThtVTl399IkqEif2HYhM8YTMystuwIEFCibQ+bR
hxRUY+Kh0XRrjv0YTZzH+QUJTfjVzpnp5zmmBOr0qaiXZxCzUMzV06jpe2oI3M3a
OosV4XmxgAoh24moI9c25+ZJ0BWIeJbA+/QeN6J616emAZihQIZnQ9IrZDcpeFh+
3em66/DbVdWJ+hELiKHGNcOD2HJhsDaHLQGmkEtuGY1UpI2WRClcmMrpcEkUvXxo
072JP1S3AGEpEguro4fac7PHu/Oa0wrVkzxDH5PIOvRY0wAy6XpkSI0wfNMmEKZc
NX+5TE/or8c5icWgOFdAUDjahT7GI4YjWF6Pn5rAwTOCLucctyse/7wHT1kDm22I
+8kjA4XSQCZfXAdEqXZ2RZnibel+bbrLCkB/4ii55abXs70OFXalIsk+6Fn8fw+p
x1n5b9LqUsT3+Eg3tGD9P0Uo57IfYY2Mum6v5c6XV6yrrzfnpjBqvxHlGUlrx+Ka
m2necX/NZ0hBXGypmob46DNqsrpWrvP8PsaXgDor53YssLPvIkBi6garcMndFFGO
0p49AIpX5dct00Grbm6ZVgGMspvBOkfiCKy9Uud5fOjMlBSJccWq2Fl13SJe2zja
DnQ0lp0XXztT1w8TgXyilh1glfzKmc7rKdxXvFoIFjyAx5kiqRX4e7KJicHrlPYX
MqwH2tdWJvbWwG1nLk9WabjM6qpaZyrMHe53rboxJyPqqvyUGEJgRGcQ7OcpnLbk
MsjsQgxjSlYuOdyd9Xl/aeT+xKO3mesKHCT/gRn4wOPGWAEklYhh5oXzZRirp/cg
62dADcwLfLeXii8FHurNlT2AOhhGX1O1F+BQgT0DpTRSintrI0Pbitt5+zOmEjjy
jLtFD6q9U9NkVEXGiHyr/wm6eqKSeFmltWhP30sKsoQUEYLO6wO2m0RN56+oInBP
TaCcfT2IAHjRRnDufS8CfB2T1Kzw3a8jhXO5xEfT9mXWdO0Ua880bnHgUuTOgjn6
3DMpD3DzG0XswzswU7DZysKXp7WGhekFjNaVY0qDXhUkupILZ33DWKvtYXKbZymh
9wjD96/O/kWFH1IeS1MBuWqCETIL0REDgqFicfIr5hgRnwHN+ZEtYzxmlAR/hqCY
lZKDe3L2q7AkwDwlPoIP/HEWbbpNo6dOm2AxcOQv5awxHET0aPhtIwMdPRwMZA2i
TySvDlHRqV0IKm6C7XRsbsUQyeONofjoxjazrqbAeNp+MBd50sfH9TC8cCry2I8C
O8jyGGwOTNUmnE4OxtHh8u0e3T2iZN3l6OdIVZys3G3sE3XcezSLrjkd6z+CpGWd
cN/9JF/mMr+2Ere7AmwPgrlobtRLGTZR0CpTyuJ0rhNZ1bvnaYfDzbq2TLaLOQAy
3UZ5iqx10GyVcBsIoMfy5vJeUzXvIJB5jNi8CUuUfywqkBykr9P559UpwiMArMwY
QU8AIMS4addOU0/SuhefOY+uixqWeCN95eS3HtirhRovWe6JX6yTdQkKxWcAkiZ/
PXckpS/Yd9h+FzKOUjLlit6NShcxtRbcYDNplO9zaZWdn5emjzfqjSAI4movy+WG
2V6vx1mY35k48TZbqgSq6WRfH17xBrCKapttbAjLwGVCZkOM4d6pOfxncTJn0p/6
q5s4k7+SZqdm5SDSf33xGJ1O1uAasJXiOXSBGcgj3JBwT91f0Sm4JQZxpDRluuuw
eFfbJjwg9wycJB4p+SVJ268FzI2gdlCurjG7y+RkisUK5x6O/sKliZOOeH4F/bNc
1OKeTBqWvWIOXsjKKnXc5osy8Di3L2QCjCVokpSPp5jATonXcUFfSINAROZYkDVd
WLKLABXhUXuHhdGGELIL22qakkE7bQL3ZLPkbuTh9xKqZcHPfs1EStGZVA+diPNL
MjiOx9bhhZj80Jy7x2v3PyF7lPamM9lJWjjzyOBzyA5eBVRj1HCt/S5Nukmi+ll5
ddTj4CbxgdcEMRe7kFONyC/gQkoiE0lvC25VrvCAtABWPAxEq0MMJX///YVdt/Zh
JU7W3WhUdR6vS6Hlq4T62ThvwprldtubPNHjSM3/uUG5tRIKcUvIv8zgvlBgvChY
2QdU9RvYD0C3zinwuDP2sfksnZHYJnyLUZ6akJ4XKySdHn+7PFelKh9DKqgHedZJ
JGxiUujAfvBZRIG8sGF6aV6xW1MfQsheRBtw8CWiHkSWAJHfV7qgRVuABbrRVBjs
NE3cS9Jn0ZL3jT8JLePfH0CeCNfiHiV090YBBxY2A1mTxPk7WyuwGECDUOAMf+hI
RW2mRSX7noXpU7Umj52r02LEoREY4i70sFoUX5qN0uSH1L75TtqFi60a0316Se1J
FLv/QhApNtCtsJXg01LPVKB9BWeB+Z0SX+6RWjS9elXd5Aw7Qulx0Og5TzAKqidG
vdasSQewiCemiB05EnaojQ==
`protect END_PROTECTED

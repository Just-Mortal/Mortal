`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5zWlBXCCY4SIq4OgRbhiCF9MUNBQ5rZIawjEl05P6N9yVyCTB1ZZq/jEkr4mt3L
HHK524FLCbhCzgReAO1UgjNHEwek+33CwuwoFLNFMH182knX6sMq7C7jJsnkZIB7
CU2JFSKyriv9cHbga0Gw4YIKDpJMZDLQdW0ounzZBCT5FOPWw8PQvtw8pqDjUVky
+Cgt4mYIcN4Df9RDqOjUxFglSy0BCGPsiGWahgXeLNpOjxFypWXWGrLA/lOqMBo1
J4nu1R4yK85leDqOt7uoQdBYFKXaPEVa8x1u9lBHXujNPsNN8OOwwsF3JMrQ5gtL
G9XYOVqRVedtI0JgdVX7J+z7NdO2ItTfGp9VVikE6nv/zWU385lp1HyUA3rGA08q
cY3LYWFzgkO9Cm7s1lssfpET4rjE+l9qI7lIleJDRbIfAsCjuFCJTmVUvnjNXxep
YfbQyecNIVOeilq3d+IVqoPq7Vpg+LbI6AawHysGyWppxGiCzSzKYx066/Y/ecYh
YfK2i9Yl6eX8DW9E1jkKy7Eyu9cdLOS863T0+xqFhXE=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4toshP70MrnqMR0O767+PYkLkBaqwtp6xth+SNpmLKq++G0OsR05pnWjJXdaXH72
OtnOqkvGnFlaqtX4TbR9+W4o2FTejAPFFwN3yPf3oB+A26Sxt/slERyM+nGKmxym
7wnjdvnTRchMrY+SlIZUQUVCzdejkufEQ+d08cQIZVGg7/jUPwU7CRURwFcMzvdP
LV/jvXNqJq4aGEkNDagLWnLl1FgRMjuyxDUl9ZrT6ZQ868Wmmhsrr3OKdBanTK6b
F3iwuBcsZLdXVLlgUmo0wZ19dHUp109QS4lUAsOTT2H2iBaRU3Bvuo9oFSThmijT
M4GUlRV7gKCwgHjm5FIJzGJqwmdi/AYbIyVLo7QTUSUytkNWwTeR86RYoztLOASJ
myMkpuso9sJuE22Ady+NmFSZLoPOOrx/lwBBwufDbgSdWhZt1Tma2Memk/mBk7Xf
HZEnOmJ3gKhsZMwrjOnjad2UB5xCyV2b2fycJPR410UuE0GvbCvBWhjjeLqWW3pa
oPi8YI5NNrfMvm3owakE4wnMg8fAlrEBFAdeoZUwyUyILCRC0gOVVfbkrJRUvLcG
AL4I01gJCHXKf3w99gewj/o3P4qljdNW0ICP7qRNSSEV3I3Z8K7lDjy77gf03e7c
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CNeY//B5aRbw1vV2mgJF86PCtWgS5481Boa5TZdrO8WXTMl6UX2lhqCjclQvGApu
VRl3K4/rZ4grJiW9odklPpC2rXaIjxPwEQfE6BczQAVmNVqryVVY4vz247xnaAUk
LroZySVhR/3mYIMiW835jXo4iRcmIXlii/7Aq3oowbHUaoNfVE+S/8Et6XYZzGcN
0EVPsd50u+0wrLvyTpHONZ98QtKwC69/nHWvBP0Rf38dsFxe1V0MqIge/r8p14jz
p8I0ZhWthMyUGkesmrs4kXGQaEPVqeX2TRM53F5PFB66PEGLdvT2LAQd/YdFDyq6
Zc4eFR8UntlM8vCIj9pRTsbL13f619CnmH/cqTyZL0iC7BQub0uBJqDbuosMMMzf
whvn5T2DjgsZ2TWxQ0X0Vp4QVza8UP8ZsH6g8rEY7Hlc/vaeUuOIrG1uvwilegmy
HCzcgj6emnFxrvadCeURusvaYRj2ciLgPg9hrWKhlhOn7SDUZOCp2jiN61fnSeYM
RHbkH0/Ewl7epkFJW0h9A25cCmCiyHWcTAL5Vu1jHmHU0631AgXFQTkdWvEwvuNX
fhRFLRWufNP3rrekY4Yj11GRxnkS3UdW+ckYKsxgBmHP20vPutjrOUtgz48xjtYL
5h4G9aw7Meos8dCyfVvDaA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/WoY/BA9vPU4gSItJwKuNwXtO/WgISpuH6xBmW++wDNFtcT0iWRzh3xt1ev/RLvP
LU4UZDZXUUlOhaeGyrw6aDJq7r8i1wdao9jQDn1nAWY+0UNoM+LfjWmcsl6e4L2A
hvCWrWU0jYFOLvKMSSvdUJfmFEdarKzHE6WlTIJ0/X4qmeBVvd72DONdT+Jqgk2r
lQPvImSjIpS/BBgow+FfFXJsEVqqJZ0g5kNjaABtrd+ETgLmRBrHMS+ZMmljrA1E
HEHKlooUBqwXTjuEbQQ1z0sZoj8P6tQWLo9ViCyPOkVQiDVC/apgv5hbgIV5fy5G
Hf95GJbdQvvIMbOQOsrN6X3VsQKFxupCuT4Z6ZO5MSxSbshxDk4L38T0BoY9gplo
XtZO1QkvNTFFfaG8QvYDdjfn7yIM8xLK1plGW14WfxIiqKPS521DD1t33eVT6cPT
oXDH7dZt8CtoRiyjvWNCux2BuGctdiLmWNUs6yb0kzUrssBjy0D0PaqdKrMPbziT
Kpg0FOqBtFRhPymlNQK827yPy3umWtnEic+OsN04ekby1UDr9KyDN/tvjod0JTWT
Q5/YVBfRnPYr44Qv38UAE+jhSr4D8icT+MB7YMvjyJI8FXTFZJhcyKRY5wHWDNOM
G7npmCHDNIgXw/uVapFfpd96nsij7ZjpmZnAkusArU0GdlDWVz7E8Q2jjtXUXCAC
aKsml3PjaDJppGcU0Ym4CUxn8N3orYsKUaD2CGS8SJ+l12Kj22K/5lG3ffu9HFbT
XSeqOf5cb0oIc7FsElMr/Tfkn35q1GYTzyHiWclc7oXY6cKyBcelOCCr8N8C/aBQ
apIy/c+ZfZz4GMn01X9n7FxU+0nZBirgP4i4pSepmxzly0scyQxaDrSnaJVw8h0w
4dSBbhUQ2CNHCIA1W6Bs6xHxwcGWMuxa6c1CMlcEP1imxzztdvc8eJZeGnZFfVfr
q3B8slrJvdKvAHh/YEqYrhxPmsFim+BS2/9rhSWreMGsV1BpGTC0XRfbCJa/3dW2
+zVHu3Gp4+Fa6eYxXnYM/Qa03FrH1wF8zQlcVnwkeflJZiHqYA8XzH68T1v/asdL
0V4gJQMv/E5dt8bOjRy0bM4j2j7H95MIlZqikKxIZXMcYHqS8Z6Ca0aBjkT1apgw
5Z9zpIQrgbIMNvdLeQzPGK4SxNBovlJvW5bHPJgpJwj0zVTHK501ZxIV6LOvwdiy
kVN9iUffcBvQjhWt/l5BJ0bsmzukc3wrPuUpBsfVcrIkTFfvTI5OSaMV95U6s5ZD
9RhIbBuqOf4VuSGLvePg2kQdcrATGh66hfWwdBT6zeQmPWBB7ifJq9BICyiHf4Qw
5D74uhTn+7dNAynfpQtUSDPY0AVnrabmEDw5Qp6dpcKYfzRSWrRltgZYmZ+UvziF
6TLq6+n4WAZu31eA9znkSWf+8+zme/JKZc+0EMMMMtyQ8wRlqBaUAIufX5I7HWu3
6oTpUsYD9t89WXK1WU36tcDcvA3b6vttPmgb2dcE1DRtf1IBpn8dgnocAvw4G3gY
904DjAlEbLwCGlA33zF3SsEhU7qgiU9SRWNaQjmoWArHGPeX0I2Sa6RKGQ+3VSag
4x2N4XUe6GUzSI3sPW6xEVpkizUTkRMkAxRTrsoaXFaMNq8h9tnrOOpYwdUBYMst
NhH8QnQiEylhJgH9dw/UJxs79HHWXVVb37THHiID8FaSAjCSxvEqjDRMWZOLtStr
7gBM9W5fYY2fLOQDrcYrl21z4EnX7bN01WHT8dTnT3qWJeuv8pKaLQVCzpsvreNR
0DXPadCgd+C6s8UXVgK2dcuv5li7/m9DhvqY7zD+aBXTBy6TskRDoaLsmYJgRxVf
BgbsRTilr6io5ud1gV9gGSrNw1PpONZGvePnbBkuKDTa4klnf2MLf/mBBNO1uYwN
OFEkijHTPR4mhct8Id/vVh51UfyYyn+iQqyeATfrzyZ5JKursIhfBQvH2IetkUag
IipfBADOYu+q4iDoTgE4m17SOIBgKV0lMgtx4U9H6EvN1rzJFmt2IcYQkcnGOj9P
SjcrqXExnFS1nVrahLPEtt6U1zALGT/rHaHl1iFolE7nMhQo8hxzihafupZaUXIO
bk/0xslvXKAOj/rfPQX9L7KP0afO89/6l7WvnbthbT59/EYR3gVBYVYuw2FOh8ay
VGjio5bAT7bACoave9MfGWxKC9phRplH5p80CjHW5sNy27TlJWeQS/BkZgJmJ+Np
bR9E+/OAghK2tdeXAnpMSINoqBrK7vAb/TWSQcjWOWfFo7bR0OzGsVo3ySN+go1h
RPsy/6Ks+iYD8D4BBTM7ni5CQMX+DuXTfC1+j4FVP8hTZnD9sxBcOJnrVOcAQXNX
DpSk7nkq5gZwTSWog0ZJaeKqq7wRr3lCl5fuoo0itPJhPMOpZNhPplOowzHqJwov
9DR6MzS2hFesOTbyOkA+DoFQBw3ekZ10VVNRMcORoHXZQL/qkgHTXNI1aIRe60J4
xwLW76ZlehGmbI81IW+9BA==
`protect END_PROTECTED

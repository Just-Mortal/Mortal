`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYJDhY/fKl/0X1DtIbVHcOnUUSRaVMJ3jw43jWaiO1y/MAPcvLCCiFxxk9vVACcF
+MuMsUEuW/V3wBJQqdZuinzcjqUZeSRMjKQR22CIJ8Cf5IiZxbRdquoZYRWHs0xX
oHmG0W4g1OkT/wad2EDkIm9NlnhFac8aCLH5rrg+OD+xVku6ilYSSDqnn7/Fh2VS
ZxBLzXoxYnIXrMC80lAddfcayeZnh2bLrRj5ajSolEn0BjGklznJsaEN8DqEtu2+
WDjVeN0R6AM4aSEG/AWiUuD7OoBbQFqalqghh9CbtEO4ZEPGmvdMt8dLHGBxkcoR
WRcAZHKt+FTFukuxQxWnWF+TRNtAn9L5RClti6xGQca0Av5dze69tYdD1/Rl4TTl
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mz31rIuqHoWo0Mai/w/Sk9VTTOaZrrN4eGH+EbBCdkpRhEok0GcGXYJY1uW7Yt72
+5lceTPZFlJ/XYygTQZUS+NyqeK/l+0tzL9cbchWEzp6rYOvXVpwYwWUKFAfr2Nk
3HOwv9oj0Y8RJlaBxwW7kWDXfQrHD859KHpFomfCIn3SoMFeNT94AoTYw/HKFEWJ
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KLU+eSPx2qB7kG9aXjd3wYFQAUr7iEpSprT+h2BekSTvB6w6Ct4YhoaYl2JnSFl
rH2Tuv1A0rXiB5jQ5o+JSGEYmeGIh3Gm59nNw9YWKIojfV8hDsK3M/OCpKHb3pNU
vIvTvJfnFk/POq/uWly/OwF+Emm6S2kjKYVZF/jIfIRrmgGn6srXoHxTvO563Id4
GGSEqOjrs98hhtcxnJ+ZrQhKOOy+OYgYrMGUDLxJxxGuru23PyEALm31mcJfnoWP
3mW/kflYeqRP8s0vmrVT/AlFNurAMWVxYkhwBkFZvUW+vG34S3K0qe/iusUPSBfv
t8VfrEp9fqMPLsUpXSQMb7kqLNaEbbXYGt+x2xZe0XldUd3PzJOGhgi60JlProtA
1XHMZBfkzYmBTTkS9UxDASUQPPrlZyAYtrYo5W37FfmpU3B8P+xTcMJt6i2l35Zr
uyC1jSpdHIPyaf0vaSVl//35/zx8/eVfp5YTZPMTCKFyZ/FO+L8vFYFP5+q32F+l
trQo3TXV2H5kWbgyWRkgguHQa2uc5m+4FDya6LICo1OO/DkFGOyf7te6L+IcOdpX
JIzQbxRH2CjZLVqulE4TyRST/e+zKUEKG/Qv4FvrFBgO3CVYAv79Hhc7BwjpYqqt
jsdsKLTfkhui+qenFtEZ5MPPV/05rb4/jLOfzIPR+kZTTpxGXwSgsjNVCrlO9tlT
cUHofnkk/RARK0Vov/loYBTOIDkU+l4JW86SU0zLydBl5LMyFRq5GkbMqfjcrdwA
`protect END_PROTECTED

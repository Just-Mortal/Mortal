`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uHKqozwfwgk79fb8bFZsYaIpgHYXQMDu1/hRcJPaW20e3afvF36lPBVadSCY3eti
O9wQ1cKF1IKcRHN//M3i0SZWhykE41jBtDM8fo4oNqvQgDDDXXYv9iBe8gtHBO3Q
fN9QcD9JW/eyY9MedAKUnyD6N64jce++WkEMGssyPO86kPvPBvGIsJd34j+Ah6aM
0Xc66lD9oRnQLegPkmY0Y8HW+LP/MyRFqVU70FNnQnhZB+0pifnfyOza7D/RUgRy
oYxCyh/wnk9ROILCrn68x+JWclFHwHEaxoevXWdUdIf5xtalnlgAdd2zqX50fkM2
OtMvVHUguELyIeKLHJPzQ2yl3oGnGkf1pDBUCameoj3fxLXWk1w4GUiPR1DLXwC+
zd0xFe7060cBQloDSMYIAQ==
`protect END_PROTECTED

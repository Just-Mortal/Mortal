`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mOjxRc/Qf/pjCaS85BSXRPq8wQe7Ao4wik7GTnBvPUEm9DxvI6eEjBcZpT1iZ0Yc
TxJ2HQKg9ORqHdTSEJB2PFx8OSEJeRlOFTsj8hHdgTHRurI13iZVzuqxHZtXsRhf
gwkWE1/JqnQ541aWuM0lhzE5wO6amCxzlG/tTifjG2/adxQBq3mEOj2P0MeiCiEy
iVq5Z5S31rq2gtvZoLULzM6ooMVBiyTXs8BrZDMMdKuxctopRV5xQMsHPNpvbwae
ioHDmD8yH64yHda7FYSTC02r3LUpZLNLcdcYp7D/3Z0qOywgxSAviU5UMkLNmx9C
bABQd6JDOBiJHOm1uy9YmzX7LCmVoz34YJumq3VosLETaNnv8+/WUnfzFlxVolAi
gzBuW9ZpPKWs0nz+vUU8dlI3BXavP98qDYoXYFCwV2zmiWGbmy+bivMPOutpM3kG
hoG18afSSe7rKv6pV/O17t/y4new3iWUmAUCqjgucNvLaoEpLf/kKKg0+/CQCg2c
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZAeZWvZGFpXV2GjAC/XB69wYffnLuC1MHc5g5v7JtOriizELlagL8tAQUF3r7ks
+LZkA7QEJf8SYTIvgzomL1SojgG1NZDKSF1lCPgmpW6RX0ETlS0OGHIY+yY9gX1p
w+cuRsKDnoSFgVWq5/MU4Bf1Y8jpBfkLB4mNCl2HD3XxZUnxpTyI/SBErnSK/EL/
LkPVXBIBcSebuoyF01vjv6iHfRE7WFAmq+ntyeEE4MF/H5cE+tJS2kp/CEcY2o4H
yYVJyrBggyObXFvnJ3VLby989l22ZHvaLeUmxHuMb5feViRhvf6aEufHaGqhLaKk
zeiFm9xmVsRy06b/0VQzENM1rEZkIKlo0BeUEIhJ5YF8wBP7VIR4hlmadIyV2wBh
C7HAG15LbfALLOnkEykNjk0YktEgCUViaou+EtZGnYuEhHvoyJZI4fYL1aBB2BPm
XR4EV8O0Ne8iWeh1bAARxbYeAIujMDXMYvxTHzxaJWung8PPd5FQLK3yH9ROuALZ
DdkbM9YB0XrPpiVq/C3qf9Aw162YhvdKmx2wMbaCII4SVk7jxu0Yj257s1pBerQz
HKuRclzKak2+lWd9dILe2s95C+5criIlY7cCzoEsCf9z8Lnlbw9oQTAiYct5avRO
TbW9REffbAIL0T6eS97KxvyEHKFHIwDmMbDC918whKh3ndet+gB9aP3n5KUlw/1N
ZfCiMYZM74+JYXi760OekWQ+mIHaoAadbjhUy9bmoSlIKOQFR/94/AqpHmANaZ7L
9L/6YLcmFB2uclJiXRkIVfqn+AizN5K3FFskLrcy3yp0J7CvqA8yZj6E0APfn9/l
3VHexi3plxzJafRLWR4UXpblKilH5oFn7kGE/E2KAIkJ1ye3Y0GOEHducKHrzH3L
vwpWkAnReNm27zxpbGOyYX6eFg42EzcAwjVAPAqON6coZvE8PTyyTrrqJAgxFzYQ
IANYkEWe9aGYgCW6yIoP797xm8JgIMVjHhUy/99ivoO9CB6Ud9B4gosWC9KAM+d3
xyueob+pJt4Por3QdshBpvn0di/rz6xT+mumhYSsfYlrchdQkQ75HHMB8bl7dc01
pPvyZgVaFzd5tx9sOcCiYQbX9JtPYODy/hcPGkB+9/VM610NcKcLYPaeC5opelj2
fYFC/a7mS2U4GZ2LcEDLtpbRs8SHfb+k4R+c1ImFSZvKWxP98GjTdqp/Mh+OOjZM
`protect END_PROTECTED

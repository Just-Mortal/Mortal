`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBCgwMV2P48ujdTxeNwnsxHTl95+zDBPT1NSib6KJZZDQ1+uUffKZJxBoQAV4iN1
gnjIDWGfRM77NVbGz29UYDqwtEItgZL/BYi24D/xag+dbppZHzJ91V0aeInV59dV
ELSiufPsuhx6LRw90vSddiA4W/5L73bHFoOvq8EdVrjexIW+r7/28Rd8rtS+MEzP
qfiX4d+17/shY8mtqjZjiLytOVYFE2oantzNfyCfBzMfh+ON1Xr0p+HgjkpBFneu
KFUf7yXyxAHSKLOJXLgx2ieqqAbmlX09PSgjGj2lfw6haNEPKl8cKeQZZ+Nqs2zi
pd6DrcANERhupU+EH/952pXqzvOUPQQyQL+08DVihk1gUvNwYuRGgdG0FzRRMxO6
VAv7ErUG8Y83MZFzfPi9JKbHnu35NRLR+J0zHY1mYY1wmT7tAPi9Igrb1jki4/bM
0Ea2xccKHFm37M7IRC3XDu5QzgJX47hC+beRh8zsZ9msvaq3DAg1KvMYOTiLzGFg
yIQMzYQmKiPEl0wEOjqCeKopuPpWwWQy38DxHhMjd8dYaf1fp/2NaCXwUSv6Gua4
Eoe870aIdoxFbpIcR86EGpfQuWN35alUCjzNLwcAcDi7qyBHmQ2UP1fQ2C43fX+I
vxp+fxW/CCVtR9Fnbms+yCMsjsUu/y8Cz56sB96Q+I4qCIZqM4d7hR+2q6G2wuSG
lxPi5eSgZcBf+uKFFT40fBiyDoRIFs6LPvWo9r4eRQhHFssbugGEHtNneRQ+iKpa
A1Mvn06a1XymQFcHKrsxAOKjk4VTvTb+wInt2fyqLXj7HLJmmAO42ERKSyyK3/Ko
yUoql36lUibZjFBX1ckpQnsjx+iHfWFdXTdbz1V2HTmVLhkH1v2sp9OQNkSyaP9n
0nDwrkd6EFMOW8rAkXqVnYP3AwBuRIFI6+NJvjkaSji2uUK/JeNjwSwb2TPctby4
qghEoWfs6gek5rNRUPeOpWsVqi/JMy75Z4po8jCVJRrTc8yPWQJn64+6h6cJGIwc
ZtxK1gNadJu3GhURVLGlVNQvob2056zICOCV3fkS1bPSwfsqVOaCfosTZt7h+xu6
N1uy8eJ7arRaKT25cXUaSq9OXqkqfXREmckqv5Eom3raVCQ8dDqBMa1XEaRPvJ6g
VP8oSXI8gxSiFgkA0Gl7z1wCFVUpB1Td0Sv5MGQXd6LlPUvUiSRyeWe6f8kzrKKV
/ISK/9cVnyv6wul7IABKs/5onyI5Fh+x18EGhSTYWz9E9qb9FJZgGaF6po2G5y+a
KuZc2u4c8y+1/lzxGJAX/YlI4j7P000pu5My4sDx/KWEeiGz6k9XsBw4GztEuUzh
posVTPusgTn0CZzKDRY9PNyENFAJbykonsSXUlFNESSXnb592NbJovqkD/zXOHmU
UB8MXfLkHSZu6CwGxM331AFZgyam0TB1TXV8qM0ya9Xu5VQz6sZ5DxJgG/FS+4gw
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tCSVRZouPgJ09PGe7GJWRKf3LdiJZWXLlNbLzq7dH5xKoQEVpU0G3iGZOFdkGqtI
KHvSL5aC6y5RKrfY5gHNqdfduS8/Sc9Nk4R9Amwa+gtIeLrtlETCugta3/Wolau2
yCZN3NT2txcakXeiJoBJ9XGRFyG7VmudGeF8uitKy0Eo0GtzfI5X+Si+0beSaq6F
WfdXcYTEyadkV2R/yOiLT972WzaF2uoec8LhDbjwWfcXykqnPcsKmQKibPZkh57+
gzzzEaCdLdVjCUXsS2oOL2t4HedXUe4NOktV8jVVSJg7FtOLmumcWABW9b3yO9D4
rwa+uFtosRl/povLTpULPAh7QBqB2yDXO12cnQK1hrfcUcNbuBty5MCwMjizAj/1
7kj325xuwEiC6Vmxf0p2Z/8CMmN7exArx81ydAMNDSQu2VgOgEylhMzJFHST2uWw
CH6jt+DdUbIUEYeP081Du9COMxxsIylB57Jjk2CVC7U=
`protect END_PROTECTED

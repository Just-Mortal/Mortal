`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7t3ahEnLu5dY+vhlRCc1T3gSr/uMe6UlarB4YBXdHY9u9jWyL+jwUUG+7rM/I39P
BgaRtx3eAb+aerSmubztUuJeIJVdB1Mf8D2NbJNYLcL9ENjN0+3+DBYhvZVfHhsJ
LjrQZQN7AnTqz//NiDhzbMq7wj77D5OGFoRAisTx8RV8xGAkb4d97or5i1tddDL8
xiMzfcf+527vqbaqBTtO2pT206AlwVkNiHmgVclPpjQtwMXUqdk4UsYmXRHvYNfG
CeG9H/PipWIS1SyETXUDq9Wt3yQWFMlotq4kV5mgNFN+RK8uQL+DtvxIpkEQGnRD
v8irwDeF72QBg3CQ06tXkAOIqCJzTDnSzeJP50ruyrD8Fp7+gOL/E6OMLrH9Naw3
0evHHJypGraM0P0msxobL8+yIz7tAlPdAMLzgfRgWwrRekpwF5W9vvMioLaL6Hed
JFAHXG1XdADOpa6hn36hnHnEXV91sdvOm+XQaUeG0ZSbwDsoC8GE5rYhRLw65Esy
3huommYyR55dwo65KeXDR/9DKYUy46IOluuL0wO9JLtje71BKfidntSRDNEUoFK0
sCpARzzC+Hb2YqUIzFYRrd6jH5kkOBy8jI1rKT42BvFkRGM8WlIfc4b0HNdvw4yH
gnzJT5sZItYXcOkw2V4DwJysgP8DMsPgW6AwLYOZ9niwLcOBxD0pX+ClGSF9iFyr
N213av7Ayfz2v+yooSuda920q9RGCwcBhmabYJG9IB2ivVaPGPhPYg5q99S2yM2V
1DGz1oXS1GFjXatuGnWvcffpo3apwTPtiqILoBtR3Asfpbff+nRqH9dVNzFZP4A3
LZiaje8JpyzChyCcY0rUdiawniR6yVHH903CcSEhnmktrkL6I/8r6l/8iO/dq3f8
CjUULoMpCtIQp3cxeeDU4lvWWzc4u7re0k88XcNySqiBiRCWlnMnd5Xbt78387Up
E5eo6aZBAWf5n4YAO0yimKlp9sJZxBwiiIPkuetu4nStDF6tOLIzA5W61qzSHzRW
JUeW+KQOSG3wdFNU/V4RmknwaY+GowxmNuy7PDQqKyt6ybTkpW5rHISaqb25IZAa
j8aQJUdoTx9oZrcPl/cO0FVihZhF0fl9Yeh/VuOnbZvcbqfWcXLClZ4Xx55ZBNOm
z/6nvGtaCn8frg8XtJ0RlwNIOQDLFm465cf1iEG1D/1ArtHxFIe4fMQhCgCEVRik
+cv1ekzMAiSmR5uYP+LuNQBVYhlO3V1n/DBoD09JegWk4BFIuM7bKSt8dFEA0D9V
m5nui0ttYRLuGe5h+6XYxwFIOFYJIEdzGQy4j9x7PDj0RuaIJC5dVS7hgUUOuh7V
VerlyUv6abIUSgxm3Qi2Nl6uPpR+dfkZro60FJqua3mZc3jymUIY7Fh+qaq/W+C0
csw3q1OCi8K0OWe1DxCIPdEZopcT+tc2Eqj19wQOVdng//JSht/19R9wkkH9Abo4
yg1cIM/22fk0UYe0EPBkC4zTulod70a5rq8LHijNw/s6KwM5V1i/Dj7fjCtudJ+U
Mjc7KHneAYpDsDZP74jPo0zXcDG9mu4GArO8SQeiQg2viCFlphFNsP8BE7Ko2A2G
p06Ko6A0D4PABlSoX4T47CwJA/aNnw+w+Jltm5u7XmILRHWYr1bckIACfU9mF8xX
8OxpuE+YkMfP6m66mi0xfXDMBRy8sY2F96h58fSxyOVRhueMnfGcpIwqMc88Ew08
dl7lhBkhcKaV8wRfSucX1Da496UlcOhkADA6HpJUW1pgNnkLc8yRQJZzJldhZ1vI
GojOnmcciOUtJIDznAibMEPAGPrnKK4g8fUfl1HAbugDO1HzN/QTFfJHK+P12crH
1f1E35Q/bM7oiMkXmfIKr1mfrnpfRUr02qBXkq1Hi/EIER3oaBKWLKTnGuy6cX4b
zSTZ/EJRiP/rYfXj/Wq8AI+U8wI00L/1VoRcEAyTtCKvZChkWO5kC2CeqDLHkBN/
xC0+Ep4HM+eq5CaECYZv1e5KYbLMyk2z/VfggZfL8/Gpj5GD9T796a9Ai/xWz5Vx
dwzS4MHYnKaLgIrq704RX2aMcWQE8t9fkZpaCW0cq1qhhl43wVppMhRmDopBqWEs
RoB8nglpdBIcdp9elPihW9KHYfusP94tcaWBfh8AWimlCO3E0BzwHLwW71LdErbb
npkTe3hJvM+iAa1ADW800QJwUWqLN40AvujNKQ2beJDQjXyd044GUykrWcNPSrxR
mf1H0P9woxZb2zS5zSEZXSfIXSIA6yqqgZpXQ7dYHKU8ValPMH6K3ti9aB3TuuoX
fpO+T93arvFLnsTIVZkRrrnxWmp0+Tw9eceLn38h2k7Nouwm7w0UiStl603DiW3G
3GHG6sDJDVciY6rHfhJvwPwpKG/7QvvvGmC04bTIsWsSgW39J/7WKW3kaF0RF1ed
8P06JQwm4dah0AFYtYKQD5KcnBNoZ5fuPhjX4wZwEv8Q2MVAtnPSfU3I1GyNMIc2
hWR7Rp43RaMwzfZShhmH8seA1+y8iKuf5AZ6bc5x+RdZhfJXw26RzoGyF4awJ5vg
OdytluwWjYqJwguP8nOk3RFpJaI+AkYKqL9qNovWt5ZPyceo6tXvOltrpoSwqBNO
/x6Ari/5n9tuCTnLiOuTLDnSZxcPfQnyCbMRzMsZFzpR3TpLzLziakoViOx/+51K
Xrz3VxHQzbifPbKjnuG8vs6s2OsMJjX/FFGdZKgifQG8ElO0Bs9db72bCP1Rx9Fu
iyuFEWk1v8BV0ZHv1qd2O/o5hNPAbwlY6al4EixrJO8TMsXdQ0DsbNlnP3pr3vWV
mYCSstdHAk9F14cNUTRcF1QVraePPCtwNJvSuyuKb27u1/m0c48Zy4dYOye47U26
QoBClWfgxx8M2UTkgJVNiw+91OxP0wAMUm6AzakEUjbOrCpbROxOcOOGflo6ohSw
S+pLTyN+tUeZBwYTHKBEXXyAycI+yHLMst5wGfHdoDejmVGfFuGEGfdvHxSq4UD4
Dt9qnF+o/+z2IbBDwp555jG9yNwfTTCui/TWi2UvcEsXBtQLL8kcqLUzZv7OJeP9
P9xgLPjJUENcmfguaFkVjJUJzjE38Lk9AMiUqFbC2v/D9zCcpiJV+CnKdQ/ZfPML
hv68VWr9NHZ/QILEVWRiaylCatbgFQ5LhpxgfZOlEMhGeaUY+UXdNaigWx54kHoE
aMo0t0UOC/iCPPgh/q7WG5aDPkA62mmzbXqFDo3renNm45rxwAuybVv9VuQtEFOm
KRsgmtVGTUytfwhABIoc39j4UsRaVtEg5xSurqVRdchdjTgjbcweeSK8Q/Ps+LPx
I+2EkGMzLFfuF1dYoTtcwhjCKIWsU/8kVUAP/3+CxDc0BEuA2vdAA/eWUEPnRDqM
qKOM+AkTy1MR5fa2+G1kMilplnQibWWpeXNltiUcyEZx6/sEu2zIBaxs6pcRfJZ+
rQRtR2c98JZtyuBEYLG70g0D8S3D9L91H2ay8AibDnCp+IDNo++RFFWfYnqapWJ2
`protect END_PROTECTED

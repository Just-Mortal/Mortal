`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQm7SjbC/iE/cmRQgENN3FCLNSADhBEsKlJ9WW1TdiQClYo9NSC9p7uxhtX7Ni+X
JsweGuQ2JqRTXpJHXm5QEAe3zKkhJJsGmlOb7E0MqmVWAqO1dnhvYroOzz3qKRzQ
PhEfrlbI5AUE969SfBl/R+gCM67dW+AwuVS7YEGn2ZDWe9dc6etfzr4EqEOn5f4K
zSEx8RhsUw1uNemzvnCyPatDukrWIshkP6o7t4VMzPfIUGlJDnt4FL1vXO5Z7nLg
wr3T+i21CdlaI7QmD6F3HjWh5U49QDaLW7LJqVnAWHfmeGZthCzf0LiiPKUyLPhf
T9zYJiuikMtCps8dLc/ipc54OY9tVm08E+hupPqjAKxStc0EqErdIKp/NfxrJGzX
UnUIZpcsuYH4s2Ai2dRaJ6m/XQp1/ZoAlqnJd21bQ/Bk+vzr/x9O6IlbWF6xiYXo
hA6wHeIWQyrs26P904P/T97m0ZRHx9MmusBHSYpjTGYe2uVMtJvHTlj+HA3nozvk
/yXnZp7Ou5sAdFJ8cqyrEZyvaweoc67V26ZVcdkzPQeawXCDWB6zrOrno7Xa+GHa
2gOMstAlMPEEpRIVkMvlCXv4A408FjYnYDk+U6/26q4QwVSyU4cTKWpEZCs/JFHX
lz2Q1sxnVqKHzlRSnVoorWxs7yPMDqRPXSb2pVy2ncE7Gl23gVcSV/v7unP+BnRm
qqH1a141OIWGmD7tzKH6bCCES2HDSr/dtyA0OlM27YagFuV99Neg/+cta8HO2pDS
VGXNb6SX8vPQPpVV9llU/p0Txbj9Vzfc3cC4+wxW/kTObm4SlcvMCyNrjnqeF0Ji
XAwFA6u9lwgG/qI8BQTJjU5iXMqD9LE5JkPwYoll6w/DKtQD0r5O0EtwySm3n+bk
t3EdOnoHt+plukLUVEHYbP9fje8bVkfIdnrWmTGcOjsGznH9Ii3s/GhyTSkUzebL
SuL+hP1g6b322iSzfO87snRWpptgpyM5XZqgellFGz1+xvQi4WPLkyAEq6OY3oCf
iKgH1+L+w5gJsJVfImgCUKuY5E2FFpXOsVnjaQFO0baubdIl0m3mwEJ9MM452WcV
Q5ZUEIN3xUTwnrGve5HmTRdiTbL1085sxXDo7Odzlwuh5E46A0i2Nt3NPVV9FkFd
wa694x2ce9qNduET/NjIRPXVDSwW1FGyiZNq+pKj4AIVyqIZDOfp6G6xiUj18DV7
I3QqUuqmskhBA7H42DE7S8yBDFaWzdTEaqf1SDm1l7Dm8/oR4D9TrQP+VwU9d8Jb
wBEQ6RXhg4ad581rp9N1pXEmIoX4V0AZtbsCbTS/a2O42OYsnlN/VrqabWvcZXSt
mCYAodUo6UlpqY48NqPai3fDCSTaKwT9nSFKIylAw+wallutCA922slQo0JnaBOk
JELJy/LFDvmN7Sb3VIJEedoWU2fgeGTM0W98As6akaKqQiae36YGONRdqWSELt+m
7xZElykrRswX1i53IxVqwdq5uZA8ogR1la3FfAUSbAtweL5r+oATDcTvShBMC5Vg
qp59qERGBfy1Q/Xbz9kFjxV8P9TvDkiTTnPDxQXpNZg03cxRSQjUkpz5wBJdN9QB
kS7uLZNrvLdStgHwToy0uS5dx4Hl30KgWi4wI7bVAzjNrsUa7FhUtX4qZKylSbxc
WsVBGYB3eeYIFJm/g9D6Bi3N0Sq9s/0urO+rpL+0q1LmR1rAAa6IBo/O54efhKyT
oIa9Iw7P6ltlwrb7mlL1gjOPoEoMiklZeU1/uxTFK5R2NU0pzjZuIoE2URhwcP6P
88MY2Udf6RNhKldi5RIaAj6sohMxvgAfySLcS08ZTgvMyjADLSnjAjJY9AK0hqqN
Ect1DimaMHQEgHLLeNPMQBTmRivF3OwuwCi5d4Ca0Lv6sWgTERcSfLhLZY7Myfy6
ATJm0wxyIYNHRDMEQ7RbZaBZlYmlOeDvVAz5Uy7ON1bFDR6L1z+Y/jI6O7Vvudyb
oDwl2sf0avClfqeno1sz4e2tay+zHvTSJdNhyxivT5HSuqPcrS7E3OxI74rE5QC5
5ihS1Ibdm8ZMLLFpTo8ZWTPBEvmrERh3sDczz1xj6yfAzi3NydEKkwpKPsTTPCxJ
MzJt1Qu9zJdSBfqq0DMY2LnkgfshRopfPVTmmrPMeyrlpZybEGbn/YHHvM/rKBfE
IYI127kIQwc9wo36rbfOAmRurPXKfPaEV8G7rQFSL2Kg5ZAxCcxYOp+57FWeEJnV
0Mygrfg6XXL3ixCbiKBarsTqTJTPrzuQR3WLvneXZiP8IkV3ouGLONlCqGHD+2SS
VxqHB+D9afc14c55o/fWZ0LsrzBnheMWZmi+2ZDq8wJCIq3J9Z6xk9kEXNKLa73v
7AduqfoYpVNuJ8fhsVW0dVuFq8OziFB63yI2Qrjo8Xwx5LW+V4374/2AoKuUpxxz
rs0kYiSZt/l86hDy0VZnXm2zo23eIKUxYd1r41ZxDtNuUddd38CEJRLoYKq1/QgI
FWmC8AbMQd89l7yNrKbfLzD8ReFVGPAtg87rMeUCUtpYrl/yHhhLhj3vHuOfM3QV
arEhvOjhDbS6SwohJxXb7W86tB44WHWZ6vl4rNydyYMTIloEkeKXFAeRlGvQh5Zx
aYguGUEsnntPHeneTEQYIofbWttTG4arUUq/4OyEyjIMkWkLH5HAR1Aj7YiX42nJ
`protect END_PROTECTED

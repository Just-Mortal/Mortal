`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRaxfYvYcyuUbHfpVOAGMxemboD5fiez0sn2pD58PH2n+JBsznGtuD9guQmB7Zgh
Fs+tXqAURoGgeGn/y0HSqKizDSaUqRCgyTZ6mqnN+Z9kR78vCaNFfpJg2s2xfaKJ
nb269sQBOG7kMhtE4oNHXVr7xbF5omAkH+cANRpp/fuF+FfTb61JGkDbkBHhj1oo
lrzr6My62bf5iW/aWcx5TJYS3jvRO6hzU4aXmwnHr8QYZiZwjMiAE6HuXq57yrHn
7GjZ0sfDwc6LxUk90uKhoYVaUQfhN6BRPO7FcAyUp8kxyhx39LgisUoMcqB9+MVR
YwUu3eCzepIlYjMjo0mwsKjLY5fUHG0ESjpjJfz9Eah0p4J/eJd+6l2i8FzQR2vE
TkU3pWW1jtRdLHvNWD7we/zZAXaK5pTV37Ae9zt9Hj2D78q7WfBnfMRo3Igxxj4B
l9LSVC7T4yIp/c1fjlO2r2ExCZCqfj8UM6ktKKg+5AFjnlZzzs3rUF6YfLVI4zYQ
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jt+RMnH8NLIcxh6kWKFhINEopiVbJOs45KJENEmnPHbDYkhUfdjE3rCB2kvEyv6L
DcgAvApfSK1Nhq8t3CPOubqlDJuu9J0436ndbIZTYXUouRyBHMM5u5Z1jMQgbML+
z4eOPQ+10wtrHfz/KJslVMcVkshQK9MNRJSAAKcaMI6YOYrq9gcC2UagPIQXEV3p
aCd7NKmDZxllSV972awJElpp92QD9z6KBTICKRgJeU32B7wTs54tR/hO94HhsKUH
htXPBNMlBLhuxFvlxwKdzphV4fWF3iB2mCSIWXg5H+ig9gakehVXGvqEn1tu4fH2
rJoVA8gJM/RoVvp8vXtl0JwaUbUWdsXWTlIXQpXemZKn7d0Km/lWMq0p4ZNGWkUx
eiDFStenGaflpne0n0etQJ5R55Yik1IKE+vDxnIVM1n9YVbQp9hSk0zfK2i7cZkt
FQNOqCJatCYhADEhgfQla4u8aW9Cz8DacxvfAQMh7uUcbSjhd0HiEhHOPhIxulGr
BE3yX+PCoEPRsksPBMRtSsQQ2+f54/drhRUvkWYogzavFU+PaT/A8LJKt+MQyi1A
7Pvs77XVwV3FhVNNX9ZePPlNoIg6VYc8Ee+lNfbgX0pcJbCTgkGK8duL+95onk/L
unAzT4DetMfZW5pEoc+nqj+LfJG5YZOn0zI1kcL5AuK605RZmxRr8v/sBfvytDRg
Wc6uifAHn0mfD1dUl93r5cY+IAsRpM+VxJpU7LauMSNtnG0cVYkMGluvBSnnBkB9
KEJtW9H099TjkbkUgxA+MWsmfT1j4tGORNrji1LjzrMLikYlg3Z0H+CisiGaLBX9
8MNiGxXXdcV2Xfkkt8l9dm83VHg0o7iWfM2sVWomHq+b8S9sZs2IBTpNHS11qmMw
tdB3geqhbPIHvEQpX1rlumr3dLvWKhBRA2b5gYfTir850jfwjXIDqm+zol1D/fJ7
HYkXqx5uskHjv+oQLCCmNY0VjjjTeLM9OKAX2qPyV1k=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lEV8bik7PfJHBWLH95NnVP0tcr4mR43ftiIIhwFJjL7Lp9QWvPaABorDbHj4vb1q
iIUesZUBRpn4v73VIdO9yz78i2JkoNQqSqokDc3ORnqkStUg2Z+Hr/J2y8Tv28Yq
pviEcxRaVbRzT3qknN+uzCdISYmP1awyl4mvQAhQ1zd4sK9sMgxYfUqnQmafDUB+
J3p20OADYDW/MacL0UGy4Y5JLNpcB0QQYouJo5QYV6xX9Rg696Z8fPiHqvll92TO
pDy0oStqJMCRdPt7wqzghrQtNW0JsGjV2WxPVijHjqrUs9E3PodGLdQ7Clawo/CP
r5EKrwhNAmEJ14/aTlsVr2+HGbjLYR32gKtCdxkM/TUeUnyLRizwjpoGEgSMM2LI
bHXejyj7qwDSXrp4Ltf1GMUuWkGRSYBbLPpAxT40MFRyqhfJkLSm46SYLjOH1QiQ
oNx/T8pcmYW6vutQwVZBxveMKbEgAlws8dJpzD3ZKx0kJu1UCjWGWKiz0eTYcktZ
zWJkDvqHnVR/0cKiu2zvFsv7xh/Yw3MX3c0HrHHquaLI4VFiTV4LfNN8Sv/iPki2
MmZ9cCWGO8r0WcbjC92m51/87exR+es8u5fHhmGhNXeIdlrqgUKR6Fvtz9ejH1OM
n+rjZ9aIGW13PAxzBSwYGXHtyLQ11fH4aqzx8H1PwuwZIKO5xTmLDsfk+LYn8m8h
tDhWbvobdBLl+ni0upobiwwDXg9Lm15J4fCwPJ+Cl7dxZYOXocmVcWPTDuWCzica
xQRGaUMcYzNE8I1qquyETmaosCqzkWWwjtkNEITBnK7+KiXc9W5KP5OgDqj9bAe5
KvKkmQYjG/+E265WGhODSClA4/vsqiRrtc8wUHpZraVeivTNyaA55UqZ6L2E5sIe
5c3BlhPWhyPC7ZHiIbnYkfkkV5Bvd5JhS8fkFdKpClzjnNROXHWROKVRFAFl18ob
oisLciVdtrNsRT+t25HROc317DCKPgqBLSpd5aLLBti0zAFK9SonQVrVqRDIIdO8
gQosqzwf5Ggd1UBQetuUwA==
`protect END_PROTECTED

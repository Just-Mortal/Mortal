`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8UoTSdQUHheH7VuBudD7kpE0h0H2rBn54p0rShSAstX25YzHPqapoxuMqunTwH6J
IG9wCCsbt+Q/iG0bzXMchj/pXiZlfUyt14gXxuVqFGKbqmUubek7LLG97+r2DFMj
I0Pcj71pd9tjcX0nbdnbCoeKQL1aMKwxgQXvgdTzf5WYHtXbQjePnv5cktx9tEU2
HajsMZ5B/VLt2ZAkQeZxoRDVo+MS13yrT9VtjLjtLcaS8yziGZ/WgT8bhtDQ6EtS
JzMYSkTfYCi3G1+VfQBuK5ta1V0wzCdDXBPqRm8/Jdx1f27nalkoQfRPUyEu4FcG
O0f+pmaHDavTwj2DcBVyhgQlghrctlF7ONfIXsWiO8r2O7S3t4FZTbHcB0cv4m7Z
6m+mEUe1XrhigFTcyND1FLVhZbC54bsuvmf0CcC4MSzZwmXJt9kcEWimFNamHaIT
7cacjXv7GCtcPxpq8QA6/ncUYyz2WBwc5UgTEe89Wy/lyPEFbRcLsB5LTQa/5Qtp
mkRBPhQKuWkes10cABmp1348EdG0sT35+MOSdyZCtfGfLhwmI4vp6oiPUhe+7fGF
NiBt/Bzifg8KY+GHRrVzK7BGFn+6pp1MV3xJEZsIv1u2F8yLpPs2ei52Tii8cUu0
bMIYgZeVUYO7IcDWPTJepgMQxc5GyVN+mCDxQ6LvOMap3nspMJogiVTpH6j427a2
iLNegDklNIRfpZnulJ8PvIl9ptWahTS8WCtZlbaAzqUEtHFcnqq1VlHnylqfXI1o
//pGItomrMN5T63ND/FzHhSNoEYnL8lg9MaCP4Df17g5Lt87G3DX3/4IN5gkRrG6
0UGv6bNQzccuV0s7uQAQNRZzwzSd6Cx4Np5QYh9BWuFevAOJwiV7uJokJZ5IFMLF
x8QEM95fanduFR9iDESLbNnDkXH3nF9rBhB/mTi03RHPzcGnTCwGMR2TYIEUAXnK
Lb61zTltJX/8dgkCl25YEA3lDJ4bCIPYr/FwyhS4Kr5bl01VEY26vnwOIbchsAw3
M7tYrAfkQlzJWzKwryOtPhYufCs1Odo3vwhY4P7K9TXkaSHRMhemY1G5gd6KhFEL
QvKxmZtuXtINwqmca1e1X82D/PfK+zgpvpsH9iKnmbmi/rQHxPzTHc63S+e+pSOO
lap3KByLqT8HVP3J8qEkcbaOjRxwZHsqW+jDb86mKdzUl5iRzuL3I8sszTh5/pKJ
CB6YS/g4bYEbCpOQMXIF6TuXtodLN4c2JMr47IcXBm8w14evzZiR0P7p0UnbbQCN
+h2pEy5hdYfGCfRE0s5WqnbCD20Y5CmqkZZQcLOIbrDeJnRjwuQGDmR80etsUS2H
hiQkdTvoOE8bG9NNBy9/cGdv0tnw52dE+5s4RbVEWqJBiXKjzcpr6hQb+Myb5c4M
k3qkLQxboQNFBVQQmyUe1ICONEeZkP73BIv8CXKe6aFOSeJ3i28GPFChNu2xylV4
mjS9dAJX+ZD9hgPjqTkUdnBqOctiTcg4jhHApNRp2vtlWyEhdgcwX9UfeIpzYWxs
DuXNJAyLAMXbqFEk5uljaOFWJQdMlqt15h7+L66NIvQzjAH6YmOVEcTaMRO0u4hq
QNVaQZ49OoyEcf7i8Zy0sYSbBA32uCMXe9h2Vd3RkNMUQHIbr4IfKI4rAW2OOvP8
C/YwxWyxgrlVne7RZCj3ZjODreFq1B0AZpvMilH+7DWf4467mK7Z0b77Vw9nHqBW
Hp47WJXtpSq72/pjY6VygE7RADL0PtGQwLGq/jQp80sn8aqiUSHryQCx6CvovW6V
rveFvLtrq8qhrfyUQS6IIFBgAZV5zm1f826FUG9n6u7a9RKJ0p8zAK4oM2362fjP
8Eymm0Z6NVvQj9IsZYMzEqaB19wrK9TuTIWBui3dffCecKLM0EzZiVA+McHbYGZN
0x9Zvd6at7A+O4EzXPjcyEB2QtjB4u5/Trg3tUYR4ikeOHU7KdBF07v44r9Elr4A
aYf1agETy5yI0giz+EUxiqBa0oFqD4CQ0z/sSfG1ZDWio6WTdh7GMZNIQ/l/N2LM
jkyGi3+KfPC2qjLKt3jeD4xA/9KoU2rxS/eWtpNHPmqHRXfVjM4jCENYBh9FtWrM
bJhuvKjobLzydTNG60pgEvWk+zycjKBaeuMgxW75PVN13ltzBplp+DAuIPi1BZQp
ZCqJr8r38oMc1qmfIdYHVojxpytIHHUxR2T79/5dexDbocHUtVW8y8slC/qjTvjh
1Ly0saVFi60eUOPgaANJ2wkr+xobnekjcX642+jDWeXPqIvn6bva3molXeDe3YPz
YwAlJbQrAQ3dWGPRYz4FJ06h8fu20nlH3bjRC+JsvHQwvUAdtbwyj4ce1cd1w6DJ
ONmkS49JWpEvTzrc05WM/ilv8jY50icKEsdeznWolOenNJnfvZmbp4SbRr90epn2
Avou3hgie1xPm2yIUx23wLOz5xpW4hefIkDDZrFJM06i0pontobvCr/7S8h6hMk+
PcTQc7PKTCUB/URNL/QfwEcQaX4PgfJm05OGfyEZz+VLMrzxPLNaWbFH5EVJi/4E
6IxL5Ul1wFOn4yVoTqLxgeCdm8oOjp9A3WizPQ89QqkwiRbi2sRwCZ2rhOuNB5mM
FRPOm0TklUoiq+iO7WJZzkPSrIAf1HJRGp+2vOIYAMIe22NN8dCbvaCbZuY8R/X1
IHgkWtBN1jAIaPpDYBqpPVA4oyDpTpMv9bkXbc52XA5I+v5h2U4sVWG71eeX3Sd2
cXSykX+Oz9sFPSDbErhgHU95YNEEloE3oRfCNiTx3ijWKWQJvgADqwjWeQmPTodr
aD+DsxGwuxwcoETFbOSNQc/GQBqNNVgNuqaQlNwCD9vvHQHbGxlls6WOfmC9yFVs
AiLHSePB3TSv4cvs0aYGnDCBAy3WuEUOtk9zLKT0QV5kMo7eeb60weRHoHB+hU4Z
klpEgLxJVePwK/UR9A3BLnWNcfGySzs7FE8pfdQWLHoXtHwzwrp5TMJxV6ykd6o7
6RUcZTPlpF2FJsvVko2lgljCPFr+HSVAKXp+eZmGWoak6ZZdXNBG0cmFp4Y4vG39
3CYzWdWQiz50hNAhFmWSuKEr9qzG33Fwr/mWQ/ZQbXNEVt8wjngsNP+1COaZ3W9a
dA/o8glkSkktQ3dnbf9i41PQINjr8kEwV8YKza6swO3ipXhvY02W3Xo/VIoGyJHf
ExjsYaOyj8yl4oWfC4RDcsK8wFQq/tF3mk/pExLD4WGZT5VUqy0K7jYsPY00UE+p
IkoH4kNMey3MCgCEy4E0OCDJVSDH4Oc1kyEnUlNqGrGVUMEMN6qc+soY95mS114M
nMB5g4IG5bcDexyxXjJhJtCyOk1HxwZ/NF48zEdpRWlnv/LFTBq/NZJZOP70BHtt
Hk6KvrjHOHbGHnmlrq7R3nquZ66c7pLZveGduEpiV7We1zK7XLueKpemKvDiw6gI
4qYvzyIiNR1+Uf8Zp9Nwzwbcy1IINn1/MVEnQSZukgQsojIqbShAVVD/bFOgWy+H
yiSuNSO908JfEJLmaEpIVtmfGBgKoJgxMUiWuQWGN+1wjjIJ9Qle14IoQBbGghMH
A/zAjE0g9Xu6u13j8UEG6Uc01qwyjM2geJArCCN7rTes0KQUo8U01NzQKsb9gLfm
wq38y2BOKQjSwqPdLnwmvnswQJ97utWUTEw9o0BLUotGQAWLv7jpBvCWQZOLv4EY
i4G9t4OLzVgQ/xozpiV7VOExe4aIO3b1xbIpzW10r92P+HvKJ1aa3h2WWJ0kQsIe
Dsgdfhi7oEMj059fTzCGm+0GMO0GZ+fV1YgFd2AgoO8BeMKYmEbE7zST7+DzEqpR
9D0cdKSZE5ENaGjqL2YLSKrJ5moOgzbSi+XPPYYf4/NE5c7YmVnI/t4l5FhpTYeM
45vOMUCPSTtinElPDzVVavxtN+he7zcc1vfAcoJbxNTpTA1j8/X5XR//9gt8gk9g
c4ybhvCJYsWP65bMKtT4IUNUy565USc6q/tA/PGi1/IRVqlA8oiddHNQ8QRdvkHh
1binME5npwkkGPBkEZnuTm+8DI2buzpL/4x/+G6lbdApsc9k28VmOtVYMTOSCuVa
F+2Bb3Lzb7X/2QstNtFYDsZHn8ySOo2ArJqih7o/yxpHZiE7fie8G+AUmwY6pmoB
ubJiPojpC78jZidDGjjF35k8sLcutsLIUdbG9KwXioiuy9Nmp+Hk+lxkHoAi68KO
tZ2yK4Hgp7YWPSuPBGRZXsxC2JJ2kADBXVAKsPV/qqxOMBOGrFexVSNJsIKhdCAA
+LOp0Uo5O89ikUaG+pb0MjP/MWyZtWFksCTcdy7jLR4Fx01HXYG6m8eWhxtsPBIK
LMhQ9+aXfrmFXT/QG8wFNlnViRwul+av0bRY4pqHKdRD1wFP3Gaqq82QSEyLcbhN
w2/40cfQP7ds+TPlE1yzL3LfkQiEZ/jQP6TdUW+bzKtrTwWg/rFiKXv+huxNIJXH
2Z3CeUNcl8/JGURsT8Ykp4LuiZmEYH7oCidodWT5jQjslRIMNNh3qaOmJcsHh30G
Yu2gWPoWC8TIaCOwd2R1f4CDpv4sXPNSfMGuQCpSpU4mS6UaQ0ZAor2W56uNQ0rK
CpQMtpLwra3rH+HwUKn/MXp/j+yvP2QpnZRWCVMknKY1bM1DgzvXRASV5FNrqbqp
m3hXS+OED4UtKLRZDiQSVJqO66OMIdsR7Ma3DlYKDoXrR7h0d/0eSjY3wZFVYftR
DFnSuBaBcYP9/CPcODUGFLV/fl3Ad+uCobyjB9nTrh7R2bJwFtKU0J8lb6eZUtf3
wVGLNNTkYvf6fQsAAT9pbv9imvO+izySW3Ce0X3bqtHjzDg8Gm+ShqB3zmEb1m54
0gMJjHQCciz8T6XQmKWWA2yAn3AmnuQ2pqnI45Y5xQSJlTM8UWw76ZBH/LyNRq8e
BCYR68GO+nqBbupyma9ClSIGyFxlUYzTHK0eTKN/6b5ZF3CFT+vokIVA+6y/Zpuh
BwAxYd2BbbCJYeau8JLb4h+lswUFmxEvnWdRysuxJGjF6ak+WFenwwcikCMomzIs
Jw0HaF4OATZPw6TUXIHkH4wCK73mizkJzfTemd7aXLdRGaZIt3iFFmVidN9kZxes
mNtetTFAacGiZYDJ1AGV4Kbb1SWrcGARMKx62nUnEG9r6IvELoolOXvo4R/VAIFk
gDX1gLKWvNmNDpQ5eWGsAw/o5QiZCKusHYaXIs/s8WAfXZr1uMAn2RGqA+80163Q
7I+1YFDJ2WyIc3x79vmm2t7sHXYC2ULV84vR8fMxahWBYJqHrtPokrpO+khd3fvm
G+S9siHxNyH+XIdwvcQMCjvsumbYYmFAS+2IrBS3fd9HJcPO8CHoKYqb1K+1II4L
4Psp5lXADtgjlOpnUllLZ04HJexM8HTVzDfx1Zoj8fMgd+hYDBcTSJMnWFKYVAt/
JVVEF5MM5ize2Uz3ZXGl29sQP0r9oQfLWEpHioYOn7jg4mFPankh5Hh5PLEBd7nX
9BQJsPmZ1etlsSwFWoBFas0UbURI5dkGUAKpA7VupK/Ux7L4biqvgjjyZasVuSmi
qi8x73U/vw9SlTlWZV+dmsZtWvVfXqh1hQ8UvXuONi2G4/tKYKj2L+NBMbOttKya
PfRC3Sg+tWgVWGKCdXSKaYqa7SYtnpo1p59KTf+jYWDTvjLMzGAgbIUjOsLk0rav
J5k5OPpouIpBO1vXXeyQOy/vKATGw/VDyBqaOqTkd46m7wbjG53IHno0E48jRmLh
xrtkmxc6iUp184BZt8S5QlGMM3X6fXa/dlU/QFZ6qC5ZUFCuqUpk3Br6UjradEbT
x3V04MuIOA+1dAwN4HQUnofgQlFEiM/KHZooLmREjvXejdwPVzSJxk56Vm0V4Rrj
9BQcxr6nxrQQsz4lMsyPlEZTrXOaddOApagn2DnFERFr0oiGng/bdmdh3gvE7zqv
Giic0SxLymP0hGuin7l/MTaPdWzWA4W+N11GBGUupOu5HtbkfS1GvwqgDRKqqAOH
yNYpjz/gssUv+uKEZfnhMtW8yOIh/YM8uXND1VSRAknyAdJpXJ7uJwG0vjbYHkWO
kjz85Z7/C3RCUPARz8hvhD09+D+mzGwSlrP4EF7eMc9x1wlYBs6riTEIjHAn1trT
Gysm5ORb9OUJGRLwGYCJBRhg34kkFgvZRLpLcEWb0fwfi0UV8Kl9zhOHNfm8c6rd
tSD473KEuFxqgvR/eE0UgoHWD8SVWO38/tloYCeTVHqn7QUDAmQezhsTuqsEybUm
CvARADs/ZNsQbEwyHX5k91F3vLspZv92k3/eVZtirdKGHXLVYSpbgEksCUfd9aoV
gAil3VHhd1bKwVHszvSA0KMQOiw5KMYPn0Xj7/kKZpUDLIGdxtvf/JKWkkhN/elR
RWtC5nC12ewxw+BCjMZFScG57L9xbaBzBQXm0nGNOGfkTcTmJ5un4PBVZyfI53cJ
UABzCLt/4sPzVV7R6lg4Gon9kfdYPOtZ/LvpUBUsBNCl/8hQqf3kq3vufCzgzaoD
islm6HCnmMDv6L6CSCdJZQsrg3st0Y8MdhYcuMO0kLjKvltz8ZH+QczSv2z6oOYV
ppzb1JP7T5WIbmDrwLGVI5aU6acJXsEVqqBiOkEwGliexGUdgu2auHelHaEMSObC
deuZ2U/caZQt/XqaNLjGRLN2pdEDG8Wrsj6rab+FCXLnFDDztb7ZvWDG6BEtcxzA
SYL/Yat0oLacycV9miGA7NtvSOqdn1fm+ox/0uAiKXiJTFQMCwt1Aha7LNwJEBCY
CJcuORP3LlZxFd67o7m2oIhwduDAX2dvnwXgemgD9I8WJoXeyHwM5jloqhDZhyC8
ioYaGbfhjbqqAZaGmEPgMqqenGnLxcAsqbFQ0zdtmPzQUz4cCC3B/9B9vY7lNiPT
2Nwsdl/a2UV8A2A4M5WGA4cyIhbNaMtF9OzXZTFHmjV169UdS36ZcLQmRx5gjUh3
C8DsmWkTZuAxIdwH4Yo1U7YRd3P1iYCBM+11SPe7z22Hw1S2ZFd7+VygDCLS5gkQ
aIVufwEQQOxu0fpGAigZGCLmetXSwNEBPghJ8fch1YBYHqBdTov/Qb9XaP1yzc9a
fG/vU3BlTflXm7LSp4+AiFLlokTdHJ3WYtdGlSz598MZBf+kXd3Mphc+txrEbeqN
wOYH93kI/M8d7I6FSBZWfJhh5fRLExN5QtYDQuHIDm7j4Kofh21TEhfKwO/aqh4v
TY3RRMCnRIHTfFIeQ6tvEHPhenS0njV1BC24uQFzLMX0NHc2b8pNSwB/8e0AUsdR
hfD3Kw+fJYBxqS2XqSV3wbSeU2uuZmKqvfmEYhbdFW9Xg+PcS2W9PUVvCTM0OSrj
m6WNQG6P0/1ASG8lBUUm8cx8yeiavFhS8uoWYfEqNYPBRHnocN+NIVR8XFnqTN2V
DCd8MuoADooaFD5xvfRCb4SKRmPORYUMYZWPHWmX6w31xxK554IwGqr+Aecze5TV
X3lwEds+aAT0QxXXighiG/aHdaLXPuOa/k1tcIMlB7IdjdbKsnbMqX20xXfUv0i7
yd9hCiOdAPGzKxbYVdiNFzGJwlJONWkszYP+CnQfAheSF7XDMOqeoIRguV/Wnmiu
SwvG+zbBE3NVPjicZ+EtgMO1hpx+R7R5vb/+b3cz6vd/nk80NXsvV1QWHZpMAg+S
8NzRnaKJ8BRCVFEXT81rII16YGy2DrLML5tPbkB/SITsGRusK0hoJmWxzrW7a+El
BI229e5WyZOi4WXp1fwzWVXt7okuPuxVZwwC2ulFWEJn5sSN6bFF/P+gHrucJg3j
dSHnevZV1QocBH6Ih7c+HahhJXG3ZLoja7nxzo4P52N8dQbrF4HN62ZBB773fwYS
gBJnc1hmjYYzrXwnRaHT10bk65gNPLO3gM+eJHlCxlOzIMIpK8mC5+sjXM3/PYyG
ltV1ChKrkwS3wqrAGDopnC7uuEzwByJGctK5hL9xgnORFjCnPqfg6GV5agHb2VmY
KqtucXjllVJUklMlZqw23Z+WXhPlHZpImqZvYzYJvtgkHdutCLXwvT+ZkxAhkNl8
Cva5cQuherNSowN9GKN1614JdGkENOsVZSfxYxv7FGlt2SMBB7u81fA16M9/A2Ss
iELK/2IC1GRhEFduoCEdHFl/GXvFMwk0fbF+jDuYjVwLlzaJ31YBEK4F4pxmpbC9
QJlu2ulR28K6okthx2F15ywUpO80lCe/ltJqUIUkmPrXtgsRiU+3doZ/Ie8B0Uip
bsp5LuW9wbn+jARjmxMSqRjQ3N/7M0wh7cMuANZ2rewuNBL0SC3rjGUftoLvORb4
ZIj94sP1N+kRtX9eD0xoZ/JE0LxR3sgSp4uGghXa4gnaUWC6FGi8W2hp/rQ+xmdu
toG1FTdfQURvPTR6IgsKQNb2oPOrLhiiwFbqGdLoF/xmOJMJZf4IOdzjQVvFN3Ma
9xwhUdLvFTF7QZPrF4LRSQTgGL+jZQFslPt0RJlFUApZHgET0oOA12kb2I3P++rr
uksPGdMaBDGUtsnNlWWtDDAgPtn/614dH3XUBN8mcLA4IJVp0Tu5VN5ChHBibJJV
5M6mgUrYDRKBGjLt9XCFQgWKCcosfBwSjwZCqsVF7TGqeohmn5KnyUpeDAPr1pmT
0RckQ7XM0FBFvX0F2JuTyyD1imsRdLIcjSbFFsMccJCKRG/9O7Y8KEo5caYGS838
xCwW0Exz0hiz1l9D2E33fmFZf4m6xw9pT9YcTm1yw9XKrf/z05RCCSiKL/SnMpHR
GTitiKZz75qMwaGx+eeixjEUmxEb4UmpV5YcWfXN/7QFNbJTX4FuasJRjNQWDZvq
QbTfa4x1cz4ITDpCpILaLci4fJB1eKYWc3b0yUgx9leXngccBInLZoVE06QglavP
R+Bi4c4Gm6yhaIjksvl/3pe7lULcWlZlIuUxy267JknecmePLRhiuevrhSy5mxPM
t/WU2WYUzLVaKmBTw8h7llq5n0w5/PQF8asR/16NTxslMxUvgqK2+qpw3laF9hck
NW3sEx+IZcZUKb1Y9VmVMJCf40uUbjf+9E6ObBnKuHg2SCbPc/ZuQNXZNC8sBSfo
a9UTyjQse/xRCQybIOuPan/RPgT1VbHGcEhJSyVnJLckCdSCFhcDCu/axLEeD4uI
54IFB4u2PJfGY8WSrPMaRNdcLYlFrz7yyUmdVsZ5PLhnwYZy1z+M2nR07tqzD4Yj
+cLx+WXX16xXvn6wayhhsw0kE+NksHmQ7RpZrTc+HXffBOWCLGl7c9HNa/8cpowP
hESSPYaahElV7qVXMTmPon1N6pf72ntW1hxAKJ6mdn7LlxlfmYAkLdrBSowNzOrF
6TgdBRExN2SS5iazRiLtThOdZ9ncvsJnrUX2g6aHYSeeOePRexCBdSvOEdlFL+JR
CdoC5eh5fBW81NL5PB4o2awDqDj1TpBy3nmjXMubY392gVufWILf8KJDo06KNiJV
rrDRNzZYINLjB4eRRAE9xs4TFUJLmIy2Ikc8I7316zxp/nAW3Xh/Y5HlL7VFIvYY
hfrGdkM0YQC5eePoF+03at7x9JdM4XyDdKN8O6Uv7JVVxO5C/wheapGq6TsnYau1
3X0FKfwW5V+w0GSAu1Q7LC+pAKQz4MzBPvrJF75PCF6t7cEsVQ+qNxz9wWf2Sk6K
RW+rvhdyBnhgHmgD8mMy5IyN3wdY+673xNGxQUKZkT7tzVKU0S9ELXLSGWB6ypla
YQGCUQ2hegENJZXnLl1ZCwqZLpjrH0M+am/oih46td5BTX9D01pjwL1glmQZ9ulB
nFSU6l86ppAcJTlJD1+Lg+AtAgY+vbG0sfx0jwzMnD/1OfER4gcpIdZfEpVxCc4a
NoBrD1tPnRF/C8Axt7kqKjyig50i/WwyZb4GxamkLUFvA2vPD+AP6a2hva4JG4Fx
0ia0MqK+OFtuJY3pZUIdSdQBNAk1nZW6sFGJyh3WBGCimz0pvRvXGPmiluk9oRe1
h0T2n1mBB7z7Qu5htk2vKpA4SmTDX+XQnURqoE+IHIuBC5UCA2r2AHyiSxYoXMeV
XpcNCUennEP1L9HY7uNSMx7ObvXtB6+zNELUDBAQ0A/lJJjg+E539FG3PfmlPTsN
MvrVKquyCmbu+JOJqHeDpgvzvyUxaLW2KAABivmVj2E++Fw9n+K5gRYKfNq7Trqk
1H9loFvneWQjoonhn8psL7HuYWAHZ+Sg90WQH28o+1ARCaFTJ2uKqnlnddfpXHI9
C3fCAcmIupzlvZplShkzzNG9bIETgTG9kCrte1ScuydOCTh5+rZ3L1UH0TV7Yo6B
OWbRH6XHNyT3u/BbPRtBuBPMqm7AFvl/9+5V2aBbyIJ26Us8/xc6kW3menRABdyW
bEN1BF2dL3+YlIx3rss0WJ2w7IhjbAy968AnTIFa4+P5u3P1c8wq0QhsZeWVHMxc
UCbgEfe0cCzpWT7BFP3Vylqf+Aze2/do9m64gj00jTLtVOk3w7fe13l++wIUPhVk
btsygPh+YpZ/4E185gTCc8EUX19rGCJcyfBFU8CnN7QaVzfbSyDbjU0RMXl6yjze
O6tYTUWcQl7g/WTfi13FcVAxIMrRc4E0pwkWs0jLNMqtPL3ysWxggqnp0yMDS8TX
BroP2VxRcNGu8WGQLnVBfwwp8IPBk5WPrne9EpGW4zGLuhzER6hVIDGDIVo6kkyy
gmmzkPSUOJRn+ryXq3uotxnY6VAsaDl43SOFRerURILFAFOsDYshbSTgo6pbgli6
z9CrYOL6xaX0H3mCsoczobECHFPMb66tvZz7u1INen7JYW1LZY1qMvqW1olx79fR
Wc2Hn7QJF6K9+YLbVAgHGj6Ybpma3kpRESrtvI+HYAddtF5uFNXMmQREw5dIniI6
KXahl1467KgwSljqBTWyZQRNIoa47by+9VsIod466P4TQvUTvvjbyDZTgmHb78IK
mJBk2XEUe3ytV4tLngah4m2EL1oqDsxMuWWaVmCKb6T+naXIVyFnmkB0BLGeq5sR
632Yc8BoQ1DTg37RInn5HrEw7LxDr0U6SM+RgzJVMCBpXljd3aY+Z0E4GpF7ybcY
nkLur8QbprDcFlcmUiAP/0jO9tahrkz1tqBGLqvEb20rWGATMPHZxzPpvRSnOG2v
fhLCSLpRQ5bEmLK/Vv1pHZb9icEJFs51LtCvB/BB6gGEtYANkJ7d+eEMnlWie/dE
JplPrRDgIJ4XrBVNNYT0lHjVSxrkexzUIITqSE7pvVwQf1Zs3zKrc7cQ9lQsTepn
v1emlLOAP8GlRf6LQjdyyoEWwDtEse2CJNIgHgWP6AJLdOYmLh9uB8yDKAVbm69+
fbZ3PHN5RzZSRv5nWjuHVDckImuvXBonLZ6w03oaAd8yvCM8AxLKnDitsB4nUErG
rCvPCRW06gnzonZK4YgzqtgzcmkLi7Vsb8sDtN+Pqb4W9INBHIp5dqRGDymnzfb7
kIzMMMoHCb1vzUSf+3sPagxhRg8GJ+6kJcwt+YVpAtzmHuywBEMmPM+pMedbKiXD
zshZ8AuSIyo0WapJuVnkA5HGL/pdOo4gSmJ3hvnM+/5sXL59AEaRGfrC2TfvCTo5
byZ3XcgT0R+aMJ6rapqmrKmNh5KdWvCV2Ik10dvAheYyPf/xKgvpR0bHNOwrTP5q
Bl/2mJgTP/7THrG4jkW0jfNbdjFgllg/tb5YRSjWhxQcaTyTgzmUvqXVQugI4WzU
8QQNLqPTQ1EsJCJJA1z/q6MdGopvtOBfTaoLj8uBvxt772PU7gUymKzJXsziD3+R
2rLq0kqNhlVVXlJsGI1yVodFH3dR16bevoQ/e9My+so/wXFm75Ka4GVuZFZUlLEn
/g2ZerydLnH3iI9aos77ty3WetRchz2wA/cZ3kO+n64oG+F+AhFXTenR6/RQmApg
PXCZHuu/eG4ZuhHnuh0sbx3VPGmWNkKZnfwJi1chuz9spWPRUbmMmneoKNdeexRg
lDAXCCQktu1toLODHIfo3VIE2ZOsiCSPZuexddhTVVwAsDDruYkkz5qFMt86i+Tm
Onnnt577UHh6JFvgnR6CjP/PuCXznkqzS5CG5W/467Jz4JpcGfvETlSU8c+MUpik
ghk6VYlVjO+EViRGP4bE/Zi8ZCnw+HqJ7tuf62+AH0vQM2QrNEq01owIuLXnbu2+
XkTDCHAIptwiMrgqxHA6vqmIMQwYkjWUn22F8B77M+1/n/D6p6tVmw0A7GdTEUe3
qnxJpxPP4yFu27fwTBcyWed7Qg7rptlIZ4xYssFNLZsj6zElI3s4Wt2gd8A7sXpO
WiTBmdhsglgR/X7l8KWpn+yWINm9fGxkx7MpSdYAvEngpTJpC5ZwCQhiOWFfFzjw
PQQaJhneS4aP9HTrhAFZEihwH7ObzbshF4uWJqwF4BU2n+5gSrClxUtSXWqh5PSR
+HXFsqYfMDwQY+TeDWLxmzjbDE0RVljLzbhO4HBvwr+XfGq+zri+MJYR32o4rjrn
dHjo24BiwzQOagU9RzQjeBLl403qnC5p03yKDvjj1NLByRMGpbj4kNppFscXLux8
zc1d9M6MvuOxOSHzX/GXmAqthLJMbSwdlpYQoTHGDpHlxV8vWO/tNNX8JWCqESZ0
0yR5vTj9UCnGAaS27k1kt/g/9+nAiY7Y9ZblQ/zvpmAGH5eBWxwLWIvhX+hzpTQY
8bR1YdRJeWHlU5PGKEGt1uS1nyxc8yJQrujzCnc3GbMFOxCXKAWIfpvLllnn6sCT
9XpOnhowtOBsclaaPN4bT5lyGAdVnDHAiTN2tgTOxSORMHjua43/G969Db7X87Ga
e9pi8di3+vkwX8e4k4Qfjft7IiMR+xdXWBJP53Dfr/KbWwxPM4tEQ8zEBehQT92L
i8V96AixVCcAuDx60XJLSw2ZXHLL9U6jTI5XTqRWUrtxWbY/Midyk6lA9+j8if7+
pqMytAst2I2d85NR2RyI2ll+SOhZCStpNKbwAFQY8OtbxIb5s2GkgZv9Qey7/1zg
JI+8WEzsYEdultu63jlGWrcX6ELADbEw/fr8d4zC8QORWLaLhS2+HBcENGp6aewu
1HnKbaJfgS02T+DvU0RD1UUzLpiu83kBUwoPG+88nZZDykwSc9GyiXNrH5hHxU4b
M1/YwM60NN2NQahFKWECME+Z3CNMJ/KlQB5GC0l6w8PegfacXdiIRJQzF6A1ZkT7
DftSq88Dz9FwRYETu7nlmjfOdPnSP+36DIuxeRjlYHDyiTwcfFONTCN7enHBwMIW
2hK+Oig6ByS7YCguj3FL+6Mpg3pnoSYgCBvF2S5xhMqFwiY21ZGQID0s5niKkXZt
0pR7WtsBaQIMJMgAgEfp6Ck8d1FYLkRawSA3vF6tWslV71h0EvwtST4YUZGdf8eh
rUsfUFShBBi8I+t3tD/AWYwZ8KlKiiMDci4vHRRsTM0w+Nb7E1f2Y9i4I1TfTGoH
ZtMMyDhQG5MKIwaVF3fgh8OpDqaZSa9s5jF+yvnH/7YI4sfjwEwyezg2cVOF9quG
QUWpLvT1j+vO5zaVVRKTy606iwE/nYxXvDIpOLqb4fNidfbuDUvFqi4tZetAQN6N
nQNqorRRV31AXpj4Dn194dn5wPi/aOQbWOHmOJX+YUHAWSHywoNl+nwubR2oZsx0
e+pN8yIcV8HE8JzK+0eD1tjO7SHyk8+RvsLbQoBR9TK+2eTX9Qs/rDFt6XyvSZ9n
taEBom2FigxNycrggiHTWIzCbHGPy0HJYAOeqwS8/w0WSeovPcg8H6LnWVbSr1SS
SblZQVAl4M2n3tZkBfNxNPNiZR0JZK+D/1FJeLlx34iqI2WZ/Go8AWFw/SVkGN/U
up6IxVgQhzPPAK3chdj8TnjAXCYeIIfAI9qtjQeJS2opGWJfm9x3dxoPgDbH92AN
0geaVTEQe6QIF5z7mYGLG2LmG0KOBz1ptt5udgY2tOgDbWu0z5MJLo0AOCZ1bwNZ
Hv4QfROKuuNbiujtMJWYH7m39lK2HNc6D5rp7TVbiT5ax3L6g3z9GBYEiSjyWsbF
iC4jAuRkZXRJRSXGj4YTgXAYqsEFZNYbn3770pGzrRqEEJleWIfleXJpM8ZF7bkQ
81wSBH/ZIOlivzVUgbjdnnOBeh1aB6gHu45WQZWq+udOUYXEVAccX0PxI0zoyydq
+Ejpl0of70wCW/8cWAHcrXRPRnYCcFa9QP/Bb64FsgbmgtZbEdZj3uX3y+20NtCP
S8GYzywAV0ze+S9Ma6nl1Mxt500IVCVN6pMfQJfNM3K14YlU3s8WiiGuKGbXjQs0
L9khezqHn9WpDJ+vK1+S6ssDYLVojJu6YjkKMgM1gg/0X6/XyFyHp9kah5C5mr0W
DSW4k6TpRH5adMSGMJZ3CRCNz0O5IjGo9h5yCf/NUYXU3tyL2D1Dq2Ejf1azV6dZ
cr8OCXDd0iDEFIAu9tIyguYiWjapCKU8poFc3bnzVPIuDB4XrbIRZ59XBl+hebTO
otlkAP54L6eeGF8o6Lqz/j+fXdxg9AyF6dOvKzBk0CnM3lkYs2xxgbWspYHbnNfT
2xnxgc+ACaR1RfORL1/+S6Gc3S3xXEndsDLdIyJdRzC5FS2iHj2wzfqGRZd72dNl
tEv7hMJFYEZHPjSaqlVWAR0WfrkdYT+zIvP0mN580LZ9NzScvsAwff2yeAfoi4/9
+0rqodWPBqitBECDRTiQxfOjK1NishqAsy1VGAz8zdCdrOT0L0gLat6vM7nF/rob
Y1lV7LxoZoQmANVYbAAOFzzZ1iydSCiTW4+yIhWDao0kWg2uaFZ+Poqle2fMzbgJ
nF1RkpG9QH115Kw6+OQY2HFzFK4d+wP3w5CD65/ojnYUK5Zw4+BL+C+xq33ksQS6
VttDLMK55F0kpg6kAK2Q7L6PKE5wUIohQID96FvhjxFQllWZvu9nvny0PhayLngB
O0ngXbDIhYy2JjjQwNQ/o1ddZ8ksFyXOgT00p7DRKzM/R6UPaqhzKm5ib9sJVkDg
dCEiPFeCjqo/ad/TADMOr5nYWupsB9/H6ELDk62WIIy84KyKUOEGOQuu6aDFumg3
+bEyCfUri240hQPV+Ehud79d7VZDOtwsqa0jhvOUJkdaEPzImnVtLotA7qUSFTsY
YuJpEL7laVnqXUJKSvclTA8sDFvBR9L7MOsKil5i5sRFbLpxAJOhB8z0dKDKP/xd
PqNFbR5zx6TKmxImOionyupYiyYA4yrl3YoXzfZiQTVvEDcILpKyK8XgMgGTsx83
9b47Rpub9+OTZ8j1kXB2PXgDNeq3CT0sEp5Op9y73eyaY7nlgdCZt9YKo+F4R/mC
8BtAjjpWWEAXk2llQXORP9y7L6VTShb2wpgcHxkDUYKrLzy3NjY+DDJyInRjWAn0
bsDgEyOSB9HDSBaocNpecYnJ7pI4DQQ2Ue/637J3zqa64TkD9q4RAOPQf3gie5uO
TzMtG/8rSw5WJzvHUh11xdAik/+DusFKIuoHgNSl+s91ETd6TOPFFhnbVHdDkAB6
qLw1gIZkmliCxZ4S1QDE9y5JfwEshkNgcbkS7hs8jdblJA3xaumOBgsvZI9aQdDv
t/t11mwcvtxFhvlINisPX9JSFYmJHalhyFV4Dhhmwgr1WUcdilGZRaNnQskucGG6
4SZq21PnrYeAgGiKc9wMc5FbGreC1zqAa040T9U03h0E2sKs5mA3NNMqRAhI0M1k
YRzOQ+djPdNkfnU6yKu8Qa4EDI38a6mz2nBw72A6uzUmSYv8SOnyuGYplpy0K1bx
XwsWq9EwyQ9+1cICcP4bYGTIfqiffIpb/gUk4ngTL9ZiepCOIO8o/Dte8QhK4OQg
x7nVNSrw+9XL9qFYGxarHNr+SO7GCU4D+l3Ydn0eBAOvvjyEGsXT1LxhTGvMmJPM
ppvy2UCDo9OzUSEmSp06RdlfvVjZOI3jBiL0ufFqb7uAAJ/IhfTLvqjFW6DaNMVY
CMca6E0byAl+Sbk0c+xcRwAejWkfpIe+ZUBL/PPenOPccXXk2ToHrxZJCCjMSsV8
MUdEr/YKSivGJdxWS8c7W4u9xDUJqXm8gjl0TJ5xSxjReHZFKr9oUNWGkSz4nise
OaoSzifMTeLQjefDHwUsao3KPGjRi2d8u0N8m9jerGir85Ng0NS2V7C/Z/mPNGMC
1iNgnhxInsOtD2V9f5MM46kRF+3eCfUo/sF0S/p36MLUrJXsyagB7QJdTt2DGvNI
NYEhtvV1azVzgrPqqleZn3ULydDbI1SaLv6M/qnaLgIVihVZ8//RLWxMpgt7vids
49odaDQCXW/TNWYAifAcyzXvhK3yKdPnL10sf2rutFaCJE7zg/FrsyjAMohIalr9
M0oISIbWW3l0At0M9uGEsQuBSSFoATME1My/4eTCND9LbNwMcAlZvEAMsdPW7aK8
Pu/Azsem+Usj1EYHSMIxs6WpF8TkugBuKfVydFCUR4lFFUiHiroGz5fwFrEP8PzX
qY2jjFEwHevxoIwfQOwkUFG+uHUi2ROzDt5wLG9VcuvO5LtXWlKe0v29AH/loBWM
CPvYRGhTcTCNOa69DO5q/GmORCyzpN454zusFi+635IJ/qqyIUL4/J1hjiJA1sF9
3dSrdc/OIxPQ2ydoqyHjnxkw5gpA9iqP1kZohwgUUN3+nGOrF0cLXw8SLbUs6o9D
wVQLfr8y4oUg+z/N5WBUy94/Bmj2+li3y43MPF15NI/H7SIfUED6xmugpHoeocQP
dtPgGkY6rvCyus/QRb9jfUIQWkvHApd0e5IRh7gviIE1uMeFNq7picZYkAgCrHGL
0SEvss79+/UNn3ECqE7p/WD4gmdPadGlqA2iFrya5P0IoClHQJbeVO8KcLJ1TbK3
8qfXteCub0pjt4gww4sK+SC2r5BLTAuifPFRNMw0x6BPpFtD8K7Lm3G2DrbpPwRh
2AbcOPhV7AtlDK4UU+kIpccSyTSsOBafGtpFpdLLtyiqNlLQ0ywWcFcPuQC0SORX
Dh4dZaWoYNk5H6XWmy5dDJgIohtYSPrBEnany+4HscflgYK5CIBFOmCQKdwzG8d3
R33yFFKe/ACBu/yVKz+u5UM6CalqOsifKXWQBoGWooFjx+B5nGGLewCHWwaA8/Kn
8tB08nArik8//7/kX9W9+RnEX01+Uj3v949/ey7IwHDBdsq5xW18N4PPravB2GwG
KEtDY+21xi9TjuIizMKE2s5Z0YiB2oBxFq0hvwS4ZepZhWhq48HENxmPBELoVUv1
DE/GhyjCyWknYA1+9XKhCEvPraaCInoiJJxjmHLcsuy914h9wffg0sAsGSI46tsj
uw3mQ6FP9LEPZW5M3/1p+BxwgkVCw1grAuyr5DfIX7FZ/+Yw7v92xFyvU3yGkIo0
Bz2/dxiZPp9eBaVH43IVcPnMMJ+nT1u2PMo6PEh3YRwCTQTme8X1vBqoQrCF72CX
Ry6rBPqFe+t6fOx73UHriU9w3zxiLHdz5BS8CttsBG8lV7T4k+hyCQHWFUlLgSuf
dbXoieK/POENiIdPDVv2NUX5oppGZbh3I7ExsUTR1l+XrzdR6i/N2W2P0zMbAGJ7
5PtzEjdueUXkZD/2BL3bCRywBxU9m0I63h6ISMMF6O7bhLAYv/M+UCEWHetJMdEN
NYmR1rDL+mMpp1EcUZuGkx47lTaD4lfeRapvfTi/2H8WdCn2tR1geFv+zyGmnCQ/
Tn0PPcw4lshSCfRDDa0YFKLLBteRLJ6/+LbW8rTG55aSMYKfCDfrjfIlpMvKaAeh
vftFqRb7bbVJ3mtQXmOTgMsk0yuHyfj6kLat5R/N/Jn9ayQWe70WgHHt0do+18AM
cB2Oq87F/6XmSCBN3yS3hwEwdq22bzZ+GZtC7juW2MBeCtBXGUyzn6D2WS81xVPo
UQkmliX32TDeOBf2Rt4ziQ/TaZ5dJpdp+rxZOX8m6q2V1QYA2Wu0r/qy6kwg8T0N
rLYERVX8cFFKhP9gep5/k7ZEOhi4sEKwEgsu7FIjqCZ8hCk3ldXsjFFPKfZ9x0bT
AWFSggcSidSQbwulWPJm9mwKGUrAX3sI+yk8Lst7IgQMfRkDa+P/NWwRx47HFVbf
PSKGFARPcSC8pj46Pbrn7P0GW2jWHwZBQL5ue/Xnk1l6O/eIjavYmk6VWz+w4CPC
bm3WXt4ewXodugqI6jZDSH4XwNdFuS0mw5wCO92CubBrNeMElEnK5GRQjfa6aOkH
dZR9VU/RA79taOjHtRajrvbf441jaH82SyltY0bPCYsOew23ZFSli8cGyDO21s7A
PT1deS7gUhldAFcX1GQjzrz4mNjFCnIbvJdRYSGA0PKrXzkMmxl6ox10bh8WfW0z
R/+dGhUPwBr0AJg9PGMA6wjzMWSoP5L81g8U1Q+1GqpgThppszn0GKKwmqxhqIxX
yY4C7RzcLYVviOMozWCIbkRZaDwOL9jD74pOADWC8WcvCbLXipD9NDkDQdiO0C+Y
jCZXqYzz6xvMgIPvjDSMKdm749SsnTM8ifI+IZPdJNCQefNqu55kDlvYP2biSrEh
TSM1txart4rEz58wyQMYeIgbFerjT5e4/jokf1uvUs0UiJZjjxizDi+mwHO0CqyZ
Q3X0l8REPcoRpk1dWAVCvI3UP7pYuqWKHGA+GOrM2U3NUIJnJSUO7irBLp8Ydnvf
0Mbbb/pam/vLSVhYMJ8I5wtVPaT1qBcGD9pGs9RuzzjesT0DJdyhBpHfBECbWznT
Dob2vlGui+RHHEDAGKVwNJJWVOWlXS9/SPdl/VC1Fx9UED/9A8DRcfRUZpODzYtf
aTCVaswFibdGOKrepMv4sgny5ubMsQLUJop6SYBwRvlKZnhtQceHN8HvQlQ/nUaO
XMdNDfA2Hgsc56Uso1TXMLkwxx5FTQLTNz2Mx6CmoF4MwM6SE+rLG9OimTcOSsCX
KYv+iVU4lYVo2NVMFA/DYBtf22Qy9iUze2AbNy1A+b6pNebQn+fu70MEBN1EnbaO
rgn6jUWlclsWWefQaAwX9lxfc7OzqLrWDhObUa9Qz2INO0Y28RjFC98FrDHrQFYx
yQiEWvTrKrQ3LLTKdDULsFMkCHs8yUyoOCaHuHODxMGau6dWY0D1F6w5SK3Qlg+C
DOvjmhnpbQ3PsP7UsjMDCzXNNtFnLT7eTv8HJIBw1USoYpiHzXFOb8Vt0Vdgdel2
cstCXaHj72K2hG8SWmW8tNAfYukwVzrDr/6O34ZiqROv8LfWWSQd6bQHHi6ts9La
SlFXC2aNvX+Mm6jkuxDgXd47uIGhr1nSP8MFUO5GW6d4kyWGHEpvdIxa4oOX3Inq
Pb8MgoSKtL3P4PHMaCTDaYW0ai4p92DqLYUyujTnCl5l5n4AC2lGedNYkA4T+bXA
vmVsg8gl/uLC/NOEJGXlER2aHvrT62LymvCrrmGZIBcEZ3hjQVAQXpHL+DqvJ3g0
rmTtLyVZp3wy9eG7NI3NTrMylbDHSzr3Esv4y8o+cS4JRGc1de+hjjSm1xLZIxQi
OoIw0VcH001RR+ap4MubrX63aF+8U0wVb7oicY8Zs7L9TT26bf2uNAnVYyJ4ITi1
aa6mS2DUv+mbYeTV0CMo3OaWl55sHVJQ9rkLMAR7yV9IxobfJgn5oQwnhjNZa3Ab
tICTh1AcE4sIVLFNjGrJsNZHxyM1DCeujJ4lyz8BHuZZpvbLoJFB513Ro3lh/Vxt
NGiyIzy+T7nyeLuI3GwXzxYr9D+/LvPy9WSV8xYY+oPYZlKkkzEJYvgORXLCX2Iv
tWuizLbuHfajIYmQlYudijlAFSmU175LazlDzKWyWUwgOoYoyzA1S+qhuUlP7m73
9v5jcNy2q1n/XClhyMK2LPgy5Fv7x+2LbiLcfI1o7BomO6djjqcd6/3z38iLfCbR
FKgF0jRJOXF7w3p24C0b6KAucrnOpbwbj+22UoE1bzuLm93KDU8sSR9pXLk5jeNj
DqiQTMRgxfAxq6FczmqEICHDdkEtZq+nH1qtrO9kJJA1MH/9HkhTkK48SV3CRg0N
FNxhdmPijVPebYA9jUDwV/Y2O96g6gbsx3CCEUvKFsIXLgNALqZdwgyRtz8Q9HGm
QBojbmbvchqXo15Tu4JsBSU7LN+bessP2wOVlOKlGGUVHbgktu4qVu/EIIEe+WLl
v/pqI7RzjWufyDfkJ8CXOCubsiyAlQ8JHIUpX8Y8tTTH/jsqyJOTLpHbGrY4vq3T
MTDQceEn0LtrNE5HrncY1ymDcPDUZDDtl/K2l/R1wp6o7runF/waHbnPQRSoT62Q
zsldK2cCQ9iBCegt+UgHpH92mtVZVbUpJif93j/5WJ6oq9/RN+Kn1tFahgJ0koao
2Xw60BqeowWgUCXpqGY8r6hgJAE1eHURyvpcVTl0kxSjKX2Ufj+6/5oBr/TXyAko
ptabrlfbqfYhdptpaUWiHbpex3PKjiPkLiMJvtXTq5GfgoZbylpiazsbC8MKRaEH
uEf6cSxl3GEodda51kchOBZNpxGGYdKu942JSeSPA+kl/mcko+6cb/gnn1PxOlPr
KSmdxjPJNPw1UrXCjY6fEf+nR+/qsdjcDs5pPwvuqVWOXVI60VINQuS72v+nb/NF
rOUvZFRE+03as9vW8JRVQsZM2SeBjF2pcEEM0YbQyjooVUqZrhQMRCxTWP0PSG2Y
SoBlkiTzXrTGDNWSwQfEZAc9zGv0+JmSbNAng/AbeoefJzoUClXuJxwM1RcQ3EHn
SiO0cDWqCpRvEKDicyz2zI2+aJmfiOUnZTsXqTgd8AgU4tiIBiO27BxEBPj6GsSj
acUoNlxs0uzvaZOLx55sH0ZOvMQbK+JdAsAI7fE0SHlhRPQVEzpv/PzbY1Wv5clm
8OYWDoZf7B4lo7rgyxXdFb9QHH2EGjf58DNTG6PUKnS7YfLgT4nvv8xZP/cL4Fqc
83okmLzVIjyWbUqCT4fUamxoVAIRYnbocvTeHABnkaui4euq9npG35TLRBwYucVG
qrlh/o617GsJaVCTmakKrBjcQL4vpj2SvE9qKuVtMxNsjwoxR7D7jVJQ70j/U+Ga
dK5EWCv1qF/oX5tjkrsDxQejnqdNoJ3nEcdo2lIfVLu2A57dq/bzA30Lt8cIqYf7
iW1yW5Wr+ihGyScwtQzkKoAwoHzADY0TVUQdCm9VfKgYRcF6tZpID5hFtaKYD1UH
LWxKvCELRzFCKBytq0vhXJIIPCbuVgKBPgs3wYz2wJDN5qqMu2vM9DDIct36W3aJ
FFKjxIFi9O55T/xVu537fY1wAXdc27T6E+emerd+PdV90hk8dJl9cKIJBgadvtZ5
eWFwteheKFwqNreW5vEoh48GR2j9Ddqgk03fssNZSbpYSlSexZDwLkrM6sGaRoVw
azxxUa4PeMb1tObnfsXNVvs9bDizIA2jEwbjzt4qG2X+FPbbWKiq387gfcDIlzDC
u4V0a38bWOK4YLAJk360QxdwUiS9Ihk9mxTvLPrVmfkx0GprAoguRd22UL1JyuNT
+TWvAKOd1RZ+NUKSNWfW153aGqzJ0hho9DV6XVqpU+kshAM+i/1xQVciOZmoNsMJ
0cK3rILejdDGFLL81MvC2OTdoazNshxq5kP6sT5IUkzgum7yTLZ6Gctt9qUupCSd
0MOYrs6OlNivxliAWj8XOBxRloDF/vmykrmI1MtjjlR5Vhw57goXYo1E5HrU71u4
RVikf7ID4T/hx9evxabq+p17EaWYx5vzxo5dDgP+NUzO+CsTKwy+DjqeMF3o9Zcx
Vf59PjyvemIsC/W8g0G0hQLfenYL7wjOdqMR3MVGXVpgZ3vqmlRz6o8PUJoE5GQf
QGF5wiFIqYw3QpyNJvs8LI1iLSbFhmzSVgJc8Ri+DsrFp92M2BIww8RhLlHH2n+g
qgxCy7sj/BEMUGH4CgKxhHTRiL9Iw99cs8iuuOHvtDlbWUUqdKsAtcBGMaUJRAI6
kPK3vHtB13PGK1AR4Y48Ymi2C6UP7D2chKGE8yyHFwlRUGMv29Fcnb8o661fObNL
Y32Q5dSeJrvkXykhq4t4jDRbdkMPVNjxVbB4TirjS4kAVm2ohAtokElijWHlx/PH
kbOSypXSzsRnB1VAufDV6t2ssKXCO7Ei+nqzzyMDsQBa5cEMcvhEal31XzaBjoNQ
/4XK8FfaHIJpsK3Fi+8rKWPr+AEIWk/+BupXRS49AyQypR/pA7k+5zwoGIQUrBc4
pPwHD8YYnCcV70fXiKUSQxd5N3Nd4KSeLACDrWvfiZRo8wKX17n4tQEwfThG9beo
Ge60xzoMnwf9UMygU06hHsCSXUuPNie3CLE6BQ7GUVjPlzXSTT/RNBOFSIbYyuAH
rLhCowKfY9AfcVamUuAFgw==
`protect END_PROTECTED

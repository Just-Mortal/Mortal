`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWGKJ1l7HLoS93uSuYcOadJeWzFSOJ3cgw1dX904x++utMmYes8P4hGeZhAjEp/m
5LozVXPID82lg17dj2N9ZAbT2Ww0XXPB87XtNohZSwiyRi/Dewg2Ao3IvqeKuHRi
Eiy82UFKuruPFc0OfPcYLM89+zFdEH9f7YTMsEY/ZUtZWqHuDqSgf2t0stQkVCSY
AvCd8VCU9YBAtcOgU+OlCXKjBlsYO9PDTYnZPsxQwhBEV/SIYYsDgb0opOD6dUfX
F3FYbllCsYR3fxBGnMBAYAsLZFgu4lQm0SM139B9Gh4gtQIe5pBxgwubsgKO49bM
iEvyZ7sDti9LGzipSsChzXNqQlydG/THVeH+0akhVZ+R2Cjqr4LMKauCOWVBtg+N
ff/XptE1qvTqe/qNbShS6QcmdC6yz1ik92qo4tSzuwUYbduJJmcbXCmnRNRYlV5d
1CiMMxldRJ5Xh9JWvTmvXyju4kO8Mm2FdvIv0KbpqeiO/z7+u8yCOJsi/Vwbm9gV
gLvM7vrVOt9bEpagyLYo0edttYLUbBp4xr+8qPolwI/bsBxKkFjHacyK+3/PVHnv
/AUBe0eLgTCp6+kQsscV84MAltJQ1UL/PuRcxst1pEVHllEM/uq7ObQ32ztl2esc
F9CRpS5BqqXx5d9iab1bygRpzwrKLdZ8HHRw9o6ahXaoFbwT9fUUdUAqcWQKD9QX
lQB0nF9o9rISmGebk8qeaufMgdHkJSoDYc2/KWSRT7tkNfgtUV1YL1cwp0O5I7vB
KjIMM33RRu8Bl5wvXnbfOY8sp92cGRaVjFXSWueD6fKWPwqW7hox6GLq3n/n9L9E
Bu7SvMAx3Nhr4ScFht7PBdiRngzaL4c3LQpnxY1rK/Y9pKjcEo3CIqo1HFYGjUsS
MxvJC34bDV7j5CGxUwcFZsxTmtjT1YwRXE3Zj4D6eXr07FfYNpYbkKzANU96TcHi
LbgL3jRw8JISjX6aXuJQQ4KWQUqyobMbCirEKBgYFpzcV0ALZTM6wOxzH881Mx8D
xqjvGUbTBywZE+HUm33rDdjwUsVv8WMgnv882JLG+OBX4x5FEgFMXp3r6+CB2Roj
XQrL0ryMJPVgz2Hq8THvfMYwxW0fm392Y8DO+yQQi64xo6QduN2ywnr9Bh0JsSz/
6TkDSPXfUfzEyFd5QxKFIj2TC5lEGuiioOEGHxzI7UmJ0s0z6mXPQ0nv22E0Smfx
0ViS89xWPsQqc6WgLLNFTlp6MfwHB3ERDpXQPn1aCWzfvZuBS+CgSydldNXKLkyT
1P2vTjkAmf9bdmvB/91iG5bvQC44deIqvWd3xpQBOm02/jyYmQAGSYf2EnILPa/Y
JaYGZFGxQ6/utRSFspbbK+7ZNfVXF/Q1RB17GPQsZFnsvIs/aO8C1MNBDypITJ+v
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VNaCy6ceH3cCyX7/Hd8oBVgJQxxc/xq4yfkOFAIltqfi1otFYods3FGPQ4Wtwo5h
gMhSdz1VB7yvwsyh+ium1qTR5ObTP5IVqT57QdcojxlKsjFq3bgZXliP9gSkCXPn
/XLn64nnYj2JHnuDS+ngk5EZ0FdGbADWu0Wsyxu+hfiLaltVKCeBysUvjMbgrh1d
DM547HyxHd+3wQpTswSasNuDe9Y32Oe5f9B8hrSItx4xbExedfpe1NEp4tChyhsB
9EtQGzjGNrsdK7P2zxjQqfxDBPpgS3iU+363QREjbtSczKLS/GCZEN4qzcCDbHQS
CaXCVIdNf1sYhrJ77ovXNNk8ZU8QnLsK9VQj5Tea/SUwXi+84m1gtAC3IRerUIbn
hGfOCBOAGCuvihVSTvZ612BHp4YxJ+Fpgu+vt7QPxIrOCe6gZHRxfyNSpvIlfHLf
m+KSP5aiWg93k526/WF3ZU0N7E9255S0q/RVFuYL2GOWwB0F59G32esaIu34AWBO
HVUMMMhjtwvwdoq+7qfgkmoRw2n4DXc5LVlCpEakiRwebdUsxcnsY1oyvAj+fjF0
9CJ1UZFpBKfQItdUPsvaodn9LxWn05ohANGICXLyZoLOdgFQD6U37/DcPzSVMxpM
LoSsT0o6eFdRkQ9Du9SCnVqPmGQEH194erh90fTQwJj1gc1uLx5rwLsNy9ZepHhh
kTPI35kvpbUxbmDcvmMhr2PFKn39axrAomnx3sLy/z9RhCM89py9QjAg58Yf3RBv
i9rT06W8qic7IFqG9mhPM374iXWhkk+vMPF9oaamIhvA4k0mpe6A4nhb58mJ76J4
YHXraQqdYimH0A+5XMqyS2QnfAb/dfoXYAixaKOnfHhjEc1sbIwbREATFpXBSElx
Nn64c3iDR0/0lzmOFOalnNm1hokEL/vMmm2w3gIgqmP1ELaQBzEGOiAhMt4wtI31
wbfJvrosHJQtch+Itr6R1gAFFpH0BdEtSZiynw5k2PRYuO8M696mnv9TjOE0MYPi
u6xGwex4+H4HkVgnT4f4pdGT5cmOTz3SMfEs3WH/1zI8+Rl3YzSb0M2kiBdDB23X
pkC1Ov3nq0g4na4noA55evy0JKTj0adOGwvESJe1ugPRHIBK2vmCFEvcg6IwjtHe
jfV3Q/8YqMmzgANOqCapThT0uIM+LFD4uSpTYpYtl8fZ9RN6oBhRYsCykHoM3cxD
85DrKtJPSQHvLatgphLSsIhaykkyrvIihOFT/PfgP3IDwsphp6TNntgp/f5/utTs
dvuX4tgl4JEJNkpF9dexeqg76wSAxkuCPg/I8jMppSJR6MG4k9lc+NwARkSrlDzA
3ZpPfiIiFLKl/IE9T2bAmA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RoMuEJ51doPWVeirwGKkBPBu27c+BK/o6jy83WYeM6pVaLYhVRiDUqQevK06ixx
PckJH0zI5AyPzwuHObY/Gb3jxY+sMow8MPVyicOEB0iL3PpZNImfimGD1lSGz2yP
Xwzpn8B2PJtWHeSjFhuRyDwNs3j21dsC553qqgoh4UXKt3R8v5UtuW8oqDvx7TTT
+BRekbpz/3/K5WPj5ZzAjaRO3Z0Rlz04gc1w9gkOEUxX/hKoEq2tDkUu+pakGRyy
fTFZ5r6nKdhkPfNmoWxaJAJQvxgkg2PIouiDtBSTvGSVdnF8m4XUPumVTEGb9/AP
AZwt1mBz9SroURYw8uOwqSZhPglLCLO3vH4fzY9Z44dvEzg21qi0IXxfEAXJUaI9
xQHR+0aIFw12IonYWja6trmQfHA3/0898TF5l1ArR+8wCUxT6JtUoorsRnTmoU14
w61l4F5A0EBWNNajnen7cb+sGyTz/b/mQe8C4N6C3l9zywhVor3D05bzIpN6DjKy
3sUd6bPn7/rOJWzWrfX7AkyB2GcaoKov+ZddDHa+DQCLZ5fN5lKbOdFqg4X61gDo
6LQDrBnQSH+839qLiW4o8VGxr5wGmUszsHUXIn2zgt9+1QqMpHWc3nVzdxZH42ZJ
YSh5JaTaEN7nvcCon96aUmOwJW9UZCxoYndRwDffwJR5bTNGOGjIe2S4dCLQjvrF
H5qoVcD713acsaGNlQoRMyE8QLC70Jm5IHim7VItxfY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FlgztLJIA/Bg4FB3pzkO7DOcvV/wLgvoDmCd8bYU090yqo/gMVx0jgKKnGG7blhS
sze2bq9rGTz4C2p4NnXSF2JkZ03xe8BFwy5f7P1bvxJK/jyGmOUNGvOOnfRyJi7m
/x8a/0kyHm5nGEOB6U+havjO9qllsJnS5ZqZHtkWx04ay60U+Qc2gIrEyDgRv0LB
+lNG4wEEDU+LEKxc5SIQRnr9kPlSl4JxcwO7+YiKQTlM5bE0f/IQS3dVW2gpZ3Wm
pgtZ1hbIJT8pMt3ajxznkVvj68CNG2//Bgg9E1QXLKEx/8ZR4eZZbApfPOmztJAw
dMOgGIuWZv6vKZJ7P2UHwGlJDW3VBcbe3fvLJmUFagQ9DiwuRmdPfAWWhaOrcRP+
Lr3ed33iH+YVch1GjUSpHaUEfWdLvQr0joDeiPb5NOeIZVm8c5mTjS9Z4SeDxOf2
kE05yxjwP15Zq8hN3hAysV3shL6M/lzprTRbQX3Q0DDxed9a1Jv4AKJjVQp8yL6j
n+TUEh57fOBGGZAl4bFmAupXsXgPn3iJ5JW43rKLC3NtfU82pg4fCHvqLJyDBhkA
6rZWyySgqkt8kBClQQq3Yurt5pdRKf0kfonsliFc0tLVF8seVUzKvEi7fL5BNSSx
bYJ3pJq5Qapo+vAvu/kg8ittlPzG2CFxRRtkxQn2qO6i2NTpNEvK9qTcbauPfQ6l
QPUaHuiUa6gfYD0Pvoq9PD4K0cKZ50fHkseNuLfTSBeLkIAOe95CJpZO268xSeT4
m4EmotcbysDNLORg8tB3ujzOy2sH6nxRFMnzLi3asGzykjp14a7dwrZlaZFq1K+q
KfVJyR8YXCMvm8f6GLirB83Ln+n0P0XPbYrKM1Pjn0WBjgh0lhnZnZlzSZok+e70
b/HdgFP7cUFKIFeHsa0jHhivhbs3gcGlvouyloT/+04GRle37rVne/VUOsYqvgO0
EbLQCv/jA82TYDKgcMwduOHPB4S4ZmcGkPHC1ZWCopgEhy7fHydc/jDC8OvgHemk
ZNRh5gvTIkisrzeDkSkv/kLF/KX97j9rGSXbyS/Xrlz3lc2SxaxRvKyQ2sglXL5R
f7s9ZoYe3tRFRytqdpDtkcULioYXq8a2dWIISAm7Fnj9Iw6loONlLyqVNhM7X3iP
hE+tTzq2NR2yJRL26jEwkzxFSjugMSv26qMK/oglNwxFdqQw9BbpMvtyI3McB99T
H3z20yM9rE0+JR/zNtw30yvB4fjBZtNADUk0DOLUVy3IkXVhaqoloXz0q9TI3Q3a
jKQDmC7yi2egCgDZ5A+wyFsIwFwlyx6MWNy3Difq4VLG7In6p7bhadrjGOoxBleF
Ab8FzmTKt01LlaoCsHnG3Ot6au7PnN/XeyiJ1HUwqO6U/FDm3Ebh0f0E99eOPv3m
LiWG/jujTVzr59TEooSIdQzSDxxEib2iRAOgHCHqiw0y6lppoFvVRi2rtzWKy3C4
`protect END_PROTECTED

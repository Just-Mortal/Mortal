`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmnlguIt1t9TfgsMiqZEHBvqnT/8yj1tQRWUhmQXpnSoOB/YKJgeamoHW2FTblSl
alphSafGAW/ZmEO4Fhm2dIijxFWmZabaMrRz2oHh2i7JIqRW2Xq681elpiWmJdnX
qtVk4/f+qRFJRFWp5lubfjLYhOsHZByBHiekinl/F0SOpxpJ7BYwvsp8L0zwh/aL
Tdle1m/JAlTqdgzunW4VVmoUaG2yVuTVb8FaOMlfXr4tuygSdXCSRkILf89EH6UU
HY+FdAdTgtnsB5GKjPs8pBdnHpFeKOexUvvG/Phck73ZYS91DuYVXozEBTOsKjJV
6RIIvjGXmFWjo1voh1pD1b6sozQs7TV5yJEIwEGyWXqj3qRigOJfTzf34xwKhycm
q1WvoXZsrEfwZ1o/F0jd8LcdeSRLzFphm0bvlB/V2KkdIBdPGC3HH+qb0QeftLdr
HCKo0f7eppR+E/rgEbHxxHyXU1S2lKQxjiYeF1Bqe5GPXmkIRj0joJPjPA3O2nbG
yKDEI7OrfmUjnuzx/lktel17Vz3bGVvmsZ4e9uQJETebqSKPOony+bs0LF09T5MX
SZITK9SHKMtmZCX1wwWjRSWm6kSyJTSYDS3VZ8NWnM+ROFxMGuaX55jRtZZbpvsX
m1lh6WoJUjjMBMN61py11I151K3tRm7uCepxJqjVmIzoQQsOzQclMOd/6J/Jg6NO
05zmO/2S/jlnpP4KKaZW6uSTy8t1He/e/U7dAJSWKSDrCj7sxkjpmUGLBhbJ/Zmd
dq+/dF1T8l+bo/M9vednd5sP+/4OTAuYHASFYLVEh7DWyN7xStnfxQGuoJaOyTn2
Ff1mfn518YYR3S9uj5TTDVn7aw2lX1l+JH/G/KS/p4TLcgdpvG7IukQQVVBhkpwl
PNK0Rqo//mCYLxLYdgUgt4hkeH6Ys8lrfwdVSiBJzx2LBqjHC7ivkxjpFyTne4p3
qvYT4Q+WF68F7DFv75i1DidAa2wUrMTYjuuKQtrxi4QqHp6P51lmVdyioSrbRxPI
nw/IYk8ZDt57imwWrLpcQzhgLKTWHKXF0MJXLR3ONIVLZ577Zn0myk+4naoqClWm
RTxkNWGr1Fnb1aXPxnb2KdmFxQu7jHTMNzA/7XM18SJjRtEsPuNAOeHNDxJnSokC
8mazdiQ55aH3t9CoVtb1Km4obSSoRjUZ50nmoH8KpISA5tPnYgmb8fJnbHAPuHpn
pIZsHinbhh9+wZ5O7HAlrKmcHGI5cqdp9PsC2NI9mTlidyx93j5Fe+lQNX5xI9CG
XJ24nyhycEAhSsWD6vpqJyBhJlhiKjEVKvKeex7d+YTDTgnxdFJOsc0dY0J7Hpux
ozmF3/3sMaufystys2nVL+ATaDKhSxEYu4eCfy8tEkF9eEDUCKzkOF9RpHKzinvS
DZsx5nD1FQb8tfO8SBgzI4+wHWs5VAk+xq3DHOKPA6+ynqDFlmKN+oaK3IL5io2j
68080mq+RRfHl+X0twjzxaA0V0NoGnp5xybLftUxgGJ7tdNC3Pr88GuX0iR1iNb3
mCk0cB5y50U/BxlPMFNrLgHfGlJjnIeZiUwQ2LPQmb/SRklyrzzgh28NH68L2dNn
ZrajFCfFkoUiWIRIM0kyV/fjteA4SbgASKiHswYnuhNDAoSOocNS9bFIVOYKhslc
OXStxE7bOAN6QS3F424VBpz1Meo3rvuV6hEq/4hC7rC1R9oFdlnH/ZKT1A+wMvQv
g6+3ZmKcMoCzUxpZQEEy57vTAEAXn57Iq9/XOgIN8QSAIkxPldDg6ovbTXqTnfv6
gsgiTAhw+Nb59Z36hzCP8Dk53TZLXRtvBwuHTakAthrOUpSGkyarzDGbWx/V5H6n
UjL3xe961vMf4+gTvODbAM/XKwSYJsapT5GF2MUu3G4BAFIWL0PdB8wfVprCbfZH
9rV1toCwRAAQv7vga4SyTOOgqpnwOQ4eHHzq86Bg2h/bWL+l4Fro1KdhYROK3c8I
CikDqY9sw2nCMyIuBTCXDu1YOreFnyrS7LD2zvZhBK4vSjst9CFRXpqCYFWcknq7
ReqrouWoIST6IYC2Z0Zb7uXzI/LnQ3nik7ddJVyMGj4a3YsUxgqUQineIcBWsWTn
jOvGKoV4uLSphFrY8zWmr9mhUEO3YP6YsJcMaql0m2HeMtRa0a+szYXeNfM2m4Mr
KgeDwEAkQfkq9fGUCCevI3j0ZsjUD/9BRgy9vH5dh//7nLLtk+XbFwKnQtcgGgOq
AJf+uE5yl2eah7/zjKeE+jGkkcMTSADFC8sh9Z5BLABiDH6z89gSch7FoiZIrN8V
9Ezjp3llhF7AyHp0oOXHWuwgvoE73xFYBmKIDXgF/9q5y2RWKm3j01tTvGv/vDW/
Bz5VIVFX8C4V7uSF8eKmliYQMPfotO0VTtPrnz5bM5nPMhligiYMmxNj26JOEC4z
qTnBtZvHkLrAlpreWgf166UW5eCJKoQtsFpqpXhI0sVryNOyCXA/nNH5jZj8eOC7
bvBDx3ATkmVX1EK9vAtqwvye3o9fCsFL91KCRi8iZ6j6LxH2FAHftRpXictb8kxd
9LtilNDHL2HAMeBGIGVtLHiwLkj+P56wsdzemVQnUMjvb9/nG37Jr1uMUZBnLDh6
xDzYVKcF2Ex/wTGx1Bu934qJlu5A/xZBZD+LUkcObpquGoZ7ueak3/s8SnYslQtJ
1/6nVpSOceO41dC6BkqVsvfooEo8s3vsNAFou0c8wzXhv/+3wppgscZwbQIwGWjF
2nLXM0CcsWv9O6rlEzPlVgN/hb7r+gy6AkCB9i57A2FBgLRkBqmphDxvTtH+pdKT
cIsU6V6Ih3eG+QSWmkKva4wE9HX09BXq9o8LaNasEL67ydzAQ5TmoZ/V9+VzjlxF
X1mga8aPu8yqpyi99fTaB7NdTe88oL+FaOqf6vFDhlUC4tNT6GGy0bOwo5IoYW/N
TA0Oec55cFpouP4chl8g6nYcYBK4+vt+gBv4GbeNDnc8HEZT11srxL46cGHCOaxa
7pt/Ojz9pkq4P9cwvvSdUfzcD6kgKpKFC30GlGGqh0HbZKjGm/A7VY5sy5fIe+N5
/SbBjMk3OObMK2V5WotsiMihGUaL2c4X2zDCtuVeEmvXS2S+Pzk+tt3ABLYJolnx
PKpD0aeh/2VisitnSiLduinVD6LC3JFar3ixGdx1HutPxFBqBHvo2HxW7obRDZeV
Vx1P2FG3aOEgL9ANWZ4LQC6j/9p7xo5mEY7tRbtOt5h4aGoUYFPUESXI5TlV4F4Q
ElEAxJXyNpYPB8rHLZ5Ik2ToasA8WCslcWus0+H5LR+3gMDrAehjCA7FZOcz1oTE
Ok/gdgJDvsgONR29PCpaP9yhYyrpEV4xHWrd+IRz4AhQnIK4LvNrNQqQATc4WkCD
IOjca9QZXFOAOnShOk7RsgVupTj6vSfwIjhwR1tZb/SqcSQ4snqe1EkMnTSvD8sK
eNSnf9SByF06DQzzYxETs5k2Djp7EoIwduoDIXAzJqVFEco8lnAhnqKIb8m9GnZS
dH56pbgZmQJdrIP4WK1/YJIuHyH5pWwwP5LjxRdiMJc2s+7TZfSDUoeiW3DO+hkN
TlRQCLOjMJuqewUt/vnqF/Ufs9mWByycZgaQdSl/EqtgdxEoWUvXZbx0Z6rF04kg
toWdsgq/PzQd4BZgeRmaMxdmukT5fRiJ0Vx2l0CslpEDE+UEcAbBp4TB3KODbTMV
8QZG0lYzAoTTXH/EYIoip8w+3c7kq7A702hhAzxzmZkGiCOCSZCC1J3f8d4iqrsE
rX/RFjJZEHaikZuX3BBXPYNMBToqO0xR6l05Zr6RY6RVS+ePsesu6yyyhBqZ88PK
+jeADHUitJ2pcqHCNbmcTuQPZ1ak7VPwWDEwOpHDRRAkJvg8wNpdbn4iV4ktyVDQ
NQExa3qFOe1PUiHLwea7jtWgB+IQjoEPK6ELGfK40KQY6Ril6MznILb9jYfpGoC7
bYo+oh74hgW67nZZqJKlnNBjv5eDOYMbDVN9hoCL0iGTOwwxqHBou/h1L0jVhsUF
KOZRK8HMmlqYoY9pZPOkGOS6sakvoQDJzoRFVeIueLpWpBPca5XtSjpv2UXmPGS7
bc10kFXr9E/8QFputb9VwmL8f5ajF56JBoUiu9x7zZgjZxmwGLUGUbK9ym0KBCTQ
GQvVrKBWKxead2AqpWlg0L4qe47KU6Z9UIO3PS26Pbw+9MkyW/EeoptEcNYRebrc
oRl5Cqwiq1NsTU2w6FY1lnL6XkiUa4xE2XzrYmq60xGrAoNvXbm4Ew40PR+dCmBn
3gnPY6IcWxkC28jCYrlQOxWEuaULWTQNC8x10BTWbG7unpDafiNbZkjfmMtnuyA/
V3r7Qh0KS1fkW4l1DZTNmSsAqvRH+dyHJInxUzCqVa2ZOM9YEP2F/9NyNaqAmtTF
CSt+dR5kdUePAi9eqWcAxWQTIms//ySbhgfTAWzYqc8+X6ngnHP94//FUL0hmTqx
6YjXQqmSSzhYvimNYfhJxsNALdYBhl6BAJd4538JdNOw8TNham99iS208pv52jnJ
+oG2Om037KsSgbJVNDpUrkYDosyHrrIvtSdeJ2oX6XPfUNC1d1CnvwtRk2g3EAbV
SDjAYznapiGv4xiAtra4wulgDtmvkoZfNPEEaAILdLhzkaj8rQ7J9Ijxn4yIugrp
+06zmL6okDuzz02qGdqagBfYLmfR1bivtnk7PJZkzdAY0F2UiSFsFm+9qnF0YYCj
sAQ0wY+I8whdWmfv1taLheJopiaxtcmuGH+zfpLHKneJHjMBm/4EJduQcnIahEa0
LPAjiAn1wS6x8k6Z3Ay0V6Tswx4c0bCIbfshAUfiWbG4gfLhFqIZmzxHUAB2Jb0P
uvGX32WM9yeVJxoc7DxbfFNojGLMT41CtZ67sNNCZ6Gg3Gp7kyEQ6xQVrSMPtt9/
xcuM5bDfWpOJN3DbIhgUB6471HQdHngnChojhU0S5yxCcqIqN9iU/73Vl2Q4qGhP
JA2I2GPasmiE/XXwiyhGXkfKPW3uQKKNwuR+C1Dz4ajL24uv6UCyJ5kZdX6/EHSq
0h5cbSlji5mlUGrzqLKBy3o1f9dLP3iL7F1wCPqDBJdNoPm3BaC81yDWBsmwWSGA
df9D7ecrUXb3Vkv7J/ag4HmJGJE6dSszNspZy72Vij2cukTM30+DxLbZl83yr96W
KjHyVTrdjgEdU9DuSF6ndPTjdnZvyQmYHRetOesWaZiqTpfforbKsj2IjVMpUg2g
QzyyCD4p4Q3//whYwkIEgDH2BVeB1bW1befosPy+fdmnZJquIiGhX+IbtPUVzxE2
Imr3bD8H+OIBzgN57GQNI7ZpbX4u5vL5TpSJfNs3tNGFl0LBz92uWmeEnDqcbSG0
4D3pKxxHhgLOkou1bhsopPyZuSnN+CDGQ14YWjai1vpF5uHOObjppL/d1qlwdjwD
cdWCRn6y3/1ZTs5LcpMC+cZ9VBnaRbq0xvRVY7NSjhJY7tZQshmHdOiQy82rgWe6
pMqDkHmiJJybsOxvHjm/VM7zzgsKL/aTObJZogDRhMwfyOvoLX3gNjDYIBjo10V2
xOWTZrN6+w2ROF3uWUnm5HwstowNMxQH0hFjVxZoQtKVDlpgxwxcAslSMqcjJgnM
O5U+DM73hRDdNC9xftKJ6MVce0o4I7jE/M6ajinNlHf49r22CZLAzapzAtqdK8md
TkVGRoheO0ubmueMiiXfFsJmXfSm+3paHVCbeFZKckev2+5EJvib3YexpFaVa9BC
WX5L1SchLNn5vW70Jt0KnnwHYzAdOZYJT7TWg88mL8Y1zsjMfO58zVq91moPxK4g
FVymmCXbynjFGJqBQXyU+tnBDXh3V80MgUTAii+tD826YZc6Mn02rgRC6vi+ZXZQ
eYSl3ZxD2wzYb+n1YeTYOl/ei/VZ4ufcw5YBNS3z0NlENlKMl5tGDKoZmR09SQja
OGngi5xU6jenOzLKQ0LGTrw3GLfPf2bZf32ODLqRmkYYFLzvI0MA1SpyeL3icY/r
pJh+KfCFOSYh95iufQsLOLxc+C13knXlUou0eGlU+tu+hVsP0VLPRSmC3X6UahDW
PSOKFDpMYLEx2Hp9mNlBo042rpD8DDvidfKfPuodLut4HLpKrsPhdu74McO+BDxB
KZXz3cDLbZm5EOogB7qhzlXgVnGzkEkkk/4B9Hx3h/45YNduwnEi/0sXo1mGrmpc
ZMBnAv6jjqP3TZKY1eeLhIvIMgcmlZqCCuwJa4sEd9hroY2zxbcswMqusHSBuKjh
Fw/LDIKLDFiJCl/ulbXNgwn2omcMQx3xD2rqSEO5aPw5c7e3SoPx4OxHUSWbc+h5
ZVYzK1raQZ5wzt95RSIxf6OA4Cq5BWejOv6UoI0+ISZgvvvqKUs2sGnIKLIdb0hP
gxhdoZA8UnysyrfzsU2fNp7YmV009cIkda7W3oY7cxfWlhuHNehRn13UUsJYTTpC
Pm3c2Lbxn8CoXYQlidNJTgKUZ1b2p9lLlwLkKWSjopVUJ33q68UyeLNyB/iAl2qI
`protect END_PROTECTED

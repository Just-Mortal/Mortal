`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9j/hwZlHY2lJrGQqNXVsoUKuwtwrmH0Q3y0kaYjYGkUs2Z2aRM9KOhQafhsmzP0I
+1e6LV+4+2Nyy9MtoSB2sDLnCwz4VgBPKUQmL5DpCpti4eUYe5auH8ZlLPhxk94C
du4oY6bjo92IpepV/bnGh9tRjO2qinrLUkI1KdeGjBHIfi0oouE2Axcf3lG2D0tY
ydbspOt9Kgu2DfjUhYVTrQfNljosUhh2k3ekskzTudTdo+Aas/Vsi4twjhlOAipG
yC4lMZ8i3NyKtvQV6gjoytioUGu4z0U3eU6lw3RFYOWRmlX4ZZDna91lOpbSHbxq
UOgHKNpA3+VLzrcM122Y2pBFeQPSIp88bdhcnNOsfSVoafKsZD6dNvfAqm0MD4Vh
OVUgxy57zA6xtXUCsSiay+PDIqxybG1wdtKAbYbuW4vpjRt6UoIkeqIHuEpyFNFj
EqNZKeQ/LkbGsE4LfHRFbgzLyxiMv7bCFgbX1gb0JQ8tqSQY8aOPuKtunRPKB1XT
88OHJZEUg89/Oib+E1BrNYy2wRy/zy2BLvRSgRZGGONsQaqCi/9XNeEPwoFStTXv
2fKaxi+MXuZNrIFpZdEgeARqGa3RrW4kuWATWpG0uRfM7hPA3cXWDiW0XQY78JRS
3uAV/Pwxem2Bj77B3MqiMhvap0OgHmyO+ezUt771Zq/cWsqi5ZsBRifXrwnAN14d
zJSEAAMSzxuZKIvOHUdQa5RjENjq8VOhW6eRA1MyQvNVAuobyMKFqIMhHGI7abyP
gXjSUc+X1gAv7Wd03+xIbAXvMTtjL2NBEo9ykD2o6QQWTQprfGaJWuJDPl+GfNrZ
sw1EreC9mil6SklyRceGBPJgXL80PA++sSoW5ARKMLvZ2dxmI4Uevh1Zx6cH+KD6
+Tk/QddtG7JjpOxh5DK6Yp75pH+Is0bY+HaVM9yUBX2yWnBt3mCOghfGCxmVUR/4
NOlqeyWttdNUrr7dBTqNKDCaPxEnT5DZuU+wtK97OanE4NJ65IS3IhWUBXgFJVQe
qyIQUlf87JJhKj5O69KsOR9VgQ2rI/BEtZBxprOgov/SVb8iHwNeGJJcMyIB8zxM
1E0ENQ1GvMUADO0s5EAFehxBNzAFa4seI1ENm6sYS/kzNoVaMXl4QTeEmxFnuFHt
Rc9KCl+qmBgliVsEOUXYZzDI7D1C614q+y2DDc2Ys2g67Uma5YnAXCeFzzPC3JS4
J5axSkvzbcmKBppD4GWU3Ui2wRrjmxGikv6J+DViErBUjl7wJI9mLZOh389OkhI9
TMBtuwFgv+VksHjShhoK8j8gUpq/RBU3smK23PVulSIIlcJgeBiWMzWU7UsivHUI
D7oiKuLZkfeJuAzBcEZYXjYJNaS4jGUQcSNkKAt5mtEuZKO6pHyX2lxjRqkNfOYv
192aaVz6DGP8VVjL2EmaSMyuLtdMJmi1JdqTbh//0wdoGOkqrV/F9P4KKkupSpVs
kQRe0cOAT/PJpcvTBqOH3I3S86L8NCC9ZllfdJ3XYwZguvIpbz6/xAcIPCqqq3b2
grxeVo9rA1uMxWx5SoR2N5abgDzXmcNTTXDgbzcaFiDEYhCvxQ5QuDIWHiiyVQWa
Rv/tgTh0qWsdHXVAG5xBV1eLmUV7GACYHQ80+tD2r/GyOZNIjIK6Pd7BYYXrSiOU
1wQROGeIET7AWozGXbW2KE5IY5JyPIEsxzwEudq2rAZOpuuGq98MQKMe4SqxY5lN
4O0x5r5sQ/z5zGCJsf78J1sXJx9RgL32WXC4c6P4QY8=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tmYJPn9JVCkb0bW7PNtnmDyfCBJPWWUC9obp8B4H3Ae5yac8MY13n8EkP8O/m20I
zPS0yKTG0FS+rxDvGyNCgH3bBV4Y1EOysr8MODc90CKGmpM5UZ0Fg2w131BO4nLn
pQpFT0ImdmuRfZTaI7hg2b9Ey2Aq9xp8Z9Cuxc3Pa8Cr2Y3N2Y95ONq7soEMHw7B
aTRsBJDqAciu+ddWQgDzjfe9gnDV/jKBQXGpUrPQmM0nSF5mlPEqNsN2KiRGEpQx
NnUBtMCbGB9jGyu7xvY39onukrPTDlEfVNuxbj1ljx/J3k1agpnEzLDAiyT+CoKe
dT0MQX/p+Lo0nQpZEdNlUY1oeM7eSeSEEnaJ14hAVASq8U5NHKRI0OcLGIWZqmAK
XX5qsqcCb2Hz5jn9bsf9S/qL2xiWmSXYz28GQetbJcerpJKa+L9bv/tFTWTAhmHn
bmMPpl4N8U5CEEhT3pry6aO4zU4FJEfibP/cufwr/J7jvmK1HAXoY0+IY1vKTBoB
IOpn2c4/qH4MI6GA9//Qi/xuJCvC4pNwtOgAz5YY/LfBZncXILg8SOT1CHmPvzBd
jDnJTR+qBHdAi2sN+NOb8qfvdBaDZGybMa2zq1r3aet3gvSGu5aKsH/xmMFRcT2g
P6dV+yjtjiejbkIpqsa/iydRBlAxN7fYydPWD4HbrUCfzpeZd4xU6PVfUvhGU7E1
8tJNCjjptNaVdNIVkE9xvRA4wX1T4XBF59T6uW1kq5hBZ8Xg5YKMWFtim1o8QxSM
HveaUAtkqxs8bcFLB1xG5wN5r1SEkergczkEp///h0ozjG/gYw4iQjlsWZ4Ch9ID
88fFhfyz+ic5ejZh8fsvnqnQoMT1+unvjWHNYfxzBSjsJkcX6ZwQSxSDrGTnVY1u
0PYbLA1JYSysPiWucbx3wg3gIXbJIuDAT2IhXTNQMtImF4InthoGqMLxbs4ZqROG
qOEQhTWbpYkrRoBJ6vm0dOKJ3GnjR+QwQpUIXJ3BdX3jIrHSvHh2eaU3XRHHYGCD
j96JDtFVG0EhTaHWKUBJ3mAG+4ilwwKrvJ6gUNX0U/PrqKzJkssLFvaM9pP+mU+R
evt1GpYQZQOflqUqCMqM/8+Kpg98uMUZbQK71bSA+7olM22K+olLLORKHd09J4ug
SCF3XB3EpXzVIOa1q4DWLx/n7snsPBw120hF5s73zJl+LfzzitVlrFx9DzRM5YiP
jdfdrG0ZwF3Mt6jzKEHQ64GYEeZtYjllAqnrh1ozuDjUS+4atp8pmog51rUK7eUd
n3gWz/Gpso4uKxgCH08Tz7Hez011KDMAHaRJUcCOnb289n/x1EGuv11wj3FV0Pli
EfBh+7SqgxfQI1pWSHfWhgRWSxzW1sYx1WIjva76aiOopdk5eqpJMLR13K5AR+Ay
edrNXkRSx8jtNqvFIefVrP1rqJNyjGZFuib7P2sgB6XGd4tqt/qXcYGNeVgeCm9U
WcxpfudnFxryPo3fNT9mn6IEHdPDhOQJi4orU2A3/36+ps7f9ZbXGWhErKihfqoo
qriwLXZ74ZM8F9xPFrPDOL+4YjgNKSdJFiih+YB8kB9kygyS3Q7LJ6pxO4UH5t01
RIlQBIxk6lQI5UQvhPyaT1z/L6AIGmsk75k8v2lpXcY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YedYLVXuWv8q/1iOe6yy4IyupTryASYc8bEcviL5al4l8oAN4vh6HZXhYIZcTXP+
cfQ5W7p8EaRbDd7TxTGBrn447Isi5JvgXBSKACGQm1f/5Ns+ILtpCVVrFBaZ6hY7
oCwld4R9TLOBEj0lIy4UEJSFQxWtoeQsbDdnpTssIkm3CuFzmPmcHSxl/WI4GPJz
TZtMSCn6/DUsTxyPzyQJQymJ+aqGsEEDjzPiCz5yOKEeC5eYELhl7jx9ArvG6YK6
sQM8iAyWnWmv0QapVI6tUjR6ywv7//K6L3KpanWLirVsjVCzhTkcDfcgSYawwM1B
xwQO2RPg582MVn+mEAudxGGWIknbp/5NTgYCjbA0KVk1XrzdwGLw0vjKFc7ZAPcb
OU23Bp3UYJjiDNYhgDlRB/N/XvPmAUdbSNiQjv0lL3dSo+e1Nl4pRsNbYOYhVpLe
4vbJz+cwFWAPvxs4u1FFmCvgQ8ja195s34JG06Ka97B8esjg2sIaJX6PlYc4q0y4
qCSWMOe4nIPaj16/issp897swrVgSwaVHEroP7iS+IewsvNmiEeiEoKRF/9jSID6
0oF8bJOU6J/XsaqLsZWp8CQ9aEmSLufskYM4Y/Sdg8zBMmJa7wURUtmMJZ+h4ohM
vmrAexQODKH3EBkSNNv97fcDQLdUAyx0umVpHMBxparNcPeQpCqVEtV3EHq0uCYt
ehphfWTXAdPuHBJKLDMHrVtHzkfUY1FESC57KHJmcpUiZdmsS9pnKA/rp73U6R2f
xrcoPrbtP0TzqNJadSonomHsFIrr8yBujccg3oq+qwFWJTL3kowHmpEEOErCV6/U
jttQ+Adik6RSWSQZObVPthp2cPcg19oe+iE3GcSMXfXeUJb2rFrr/vg3feoUzpax
6XzE38+aOIKOQRJL6lkxzCH6YKXfjTnde2JUglZVkTS4BhkhzV3tMPb3OPYnepJR
XQH9ZehRHkYOQJJ+UBDCHkyvVMn/cLKm4tISmrCeObl1o0c8Xc8TK/djUgnw+KPr
t7Ov2DCzZc9V5NhfLsWRmF6LLykq9WuOj3MI3lwWIXb4lcKjeTPNkRcYVECzZzvV
qOTFCuaIPC/fH6AtAKBC3Lu+COIEQ4q8qnXAa80uON7J645rJW80iFWPVxQBZxDX
gr4AzlbzNXtuWV4WBZRAS2edkaezyfTAwXZkaXnA+znJBgvDgCnJFlLcBq65lL8f
9F3Jg2qbdxPTRsEH6nD6nQRecoK6nGSClYZxwOkKuTL/TVW45xSb/3UuQc6lOkFo
4Kut+affMhCBgGrP9ivTZVDhMmaF8MoE08KMuRDFvEuNtVIh2QOtU3JVRICwgrOj
mg0ZtXJwaQwSDDwyXwFKCamsE7P0U7Vz5FuOraUfvWy+5HGfEMp+SZcSe2VVShEU
PcYL9fyNdsHGqgqvnrDI5IBubFN8Rx5qLrspoMYcwYI=
`protect END_PROTECTED

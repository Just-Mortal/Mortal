`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mbtib8o3+1JGFSNg2MxXBK07vLf3TxKSH9OjST7AyGrhx3uP0eZ81rNNsxijCDzI
1mV7MLKULtV67dCgWBW8vwUa7KWrXhfpcjkHlHGeLeTUM+8hJqVyVpcbOdxQ3gpM
n0SAEYRu1RqavDaJX/WlypOas9vcERI06FW63k3g3XtNlgdhJc1a7eldF9b2epbh
fQkp2uRDCA9I526SRPzGJBRzUpH4Jb2P8dBBTCCPHVoQXLxb9JoywU+chqr64bcz
dTUBFXtz3iSgO62wFhSHjKBuxb42OHibhxXP7nY5us5ChBZeCZ39aw3nauvqVwqd
heZb4sujjsT60AnEN8ziwRc8Lyko1Dr5Z6eYp6tI/S++xOTnMsWRCvcI7BZ+Wsdq
wQWfUqmYqKF6NZIQZIqhvvRQiQlMQ36AxlIUdHF8fBiBNIwc4aZATZl3NuZC1QC2
UJ9t0wm7lpR/AIn9+byI9w==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rr0odYnbydFQryCwEgUv2vMQG6qUFjoZi46N7nbsW7N0DrygzYe80nemAyKGCJms
67FzG/8v/yT0jBtcrjrj+yBO2EEHILaeZgJVA9H4hgWaRZm4f6S19EevJAqFdL9c
WLiKdcrn5rxfWwFxqtQiiA9L5KrHPwSM7084tsLrR/uriGdMlc2rX00yOjOeQOZn
QvxURKBWm3MzRTys04BYS6SK114tqHh8vPp0D3uO4UZGAB0XAM+UDgvryfkRghjj
+xlxcZ3Kvfvgn6Ne0aVo8f4/Wq+kyPv5ZFPmkZwPUXT39g9Onz01TI2nP+nc1rnj
qlXBfOjDxdy0/uHXzZ+jXfA5pOi/0snJm4s4nrduCBRLNQNIFvcNXt6OIhNtohTw
Se3LxaviDR7hF3XB/7juvM6ouNhboZJv8yjtVU+ll+bdNkWWk8jbkjfzz5ycEvE1
azkygFXsQ87CXQnBy3mNj/GGEz9yQoZMkFT/cZS0sCDU5GSEzrTwo9+szbWdBFkd
PvDlnciken8nEEGhUWcyBzCNtBaxZ7o0x7YvftSYFwcftfbJqpmP2j4r3J5fn9UI
UvFVmtkcVlPS7YmCgUb0xwqhsC1wdYgtOsBtH4wwbgRsEGg3V/+Br7mz61eKJeIi
NIWHSv9w+rIO1yUlOpgQEhomfqqWoEl/W7uzAhud6iUQl9A73CKpHQOL9t0Ozj45
DNtYKm7l2q3wbOHZI+9PuM7if5uS+X0EZ0iVBr+ge1iCt+M2844ze+oiYnl+v6hM
oz6g+5p3SJgSYIpf1Otbuy9bHFdYJxIXtDGIgQFkhbLeHL26TQOEZ5pi/gfbn2TK
Ho5Vog/To1r2TtpjXcKzAxOD3EMNVVzecaLyCnRzPUy2V32xkmwH3ry5etOsPKCL
frF012ssQdYSqy7HXYtCADBxInAHrrodzHO2p5sLz7SXBkzu4im/U0eO0VoLp8Vd
kj0NotAdc3gMGQIxRj2L4BFWwLPPvo3Bb7DzOGOQtuTwx+rlzOOafp4xrTcDjPQ4
1jk6b3/NJsHKlgQRNMFri4hXYJts8MAsi76bGOrrAaWqyMFQX3qA0Cq/yEupNUN2
17UQpeggkg3fTC/6p4IyQLe/jaORc4Cdv1tDq8b03OkvLJEujgpi827vPLwjlglU
Sov0ldTUElZ0lZQZq5HeWCQy3pucc6FQAq8t16HmZZhsTZjLFjtLI+KUZ8Cvq5z3
z6aXg+sQ1cYjGgPsmJ7kv3muRDfg+avearh0u4PrtJrSs/LWdOy+eXBYU4ODp02d
bfJH/IEnfbYGFyGTjpnlCk3SEzwMYF8F5oFEJE72bS+xMe4PguymZHHRJi5Q97LV
xeQaQx7X6Wp6EzQc1giLLQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xH/0cwkkDaxBfr+C4YmTQVrpxhnu3hOa0qiqpJlDiVdTvy/YRrcTLPvn3hmwu2Sq
CU9+94AGuiRKiY7K+Q21uiNKpxo6lEQ9u8gxcuiBX9s6xZWVizhdB0T+06Q5dMs/
M5XXPL4VffKN7DHCV/aI39XU0vmZv/m7CiahSvx19eswx/MEGKKJmBdM/NIwy2EL
CpgtbwoV24n15eKXyfiEpCxM/DyMl/ar+J/ZbUcP7+ys364v6dOpbyMeCrr5i+GZ
WmjMHIzs6/+MLc4q+LuZkc5jJzYfSDc/fuy6izIyBqrrP0sakTJGieKImL+X6R1/
0UYsEb7/zJmqmY6kq5dRt4cD9vHHXOECPXNTkKq5Uw4WAKWwn+M22iSrc+vahu7V
04RYystRIhkYGfZ88HmrdzW3BCm+OmKH5XG4k6PQTPSMaTdK4TVBwe2StyXqYwIa
`protect END_PROTECTED

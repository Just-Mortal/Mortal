`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVCMOiVejKHfcRQi+QgZ5x8LcLcI1CD+ufExf/lRELa6kKHykAQVfBuvtHZhCH8S
92n+i5tlmTRpLo16Yh0fGss0d0lLqdaOuy144J0SwLCi4qSriDoik4uvYRkQAg96
D0QTwPkMWehZtPGs4aF1Zw8ViK9RoETVDbRLCos3rf2mRaeLyxAoqP4K/YnBCkbR
sl8r2H2aNorQVDU9aOGL5FYqwYORtm+ebav1u58FGChGjeqWDQyWatmu+xTgGNyH
7XrTBByvlsfLbmTNpNeYGimbBX9rUaPqJOZM9oFnolTc3ZnhPpHLd6kuXUOI7f3Q
d55XPa2x8LGAEIfRNPsHM9z/stopuxwKmlw1TgmLO9eeUfH1YIbFEK1JAJjzyAmo
ckjGUReOAhSX3kYE6trLgZn7JtGxk+di9hyBRSkQADSNv9lafs+uA7qTIct/fAFB
rflfzI+K4e96QIfqjS7MT3Zl1A7HBjDvQ2jt2HELUqVpzS3I/HkYJ2cF5H+0pO07
hgTpc8IIwhkBunpy4g/v2377O8KL6HmHYrEOVgEwWKDB5gjgXE7QRjRU8CJki4MX
DqEcnLE+RAmIpXSo+q0gzcxHW6/ZqWSjlFpl8vqnuCa+izhOONk73MriOEEbLOgH
kYZCRVtoMA3i8T/7ICMF2AUPFfVkrtseP/XKXmyno4onKrG3gFm5yMcD/Iqmrsjr
J8OTtB33xXjcuqxwCb3nIuSs6I0e7CLF+GhuuXA2hjquu+e9eMvBad2wXCeIpXF0
o9nXgTG/p51l+0qno6RloKZmD/slUr4llcOQzHZOB2p2dSrWfFPyO4dcx1qAwP7Q
PmsYXZ/pHQNiDNtlp595L4O7jiwJaFmardMjFyRVv5hMdm8kZsV/XrrsgiVRb2dt
zc8O0z8vx57uJs+hM5Y/fLMXGZF1kWzzjNdfzrUbgiiQ97lghk7HXVnY27Rv7l8s
0WRM1AlyyzDBjDYdJMWcpMVgC79mqVur5TI9Iwr96ElcP1x4HSspNccYv+fDQc+D
FruIpD+aDI1CTgoXJ7JZFKjqgtgVWI6L3rFwQdcte+CkXpCKbX3lEJfAzJ2zfpVs
s4l3ZgwLgvtIc+B42voG7HeT/oLam0wBqbDlKEQT+aog5uYDXZ5xtMgnGf51FtA9
c+wka9XYYqpxsGkgeYRVsdmmUuL2hh6s7k+sBD7Oaz9b9TM/ojluZFOsUR5Mjcde
Amiw43yfXSoMz+Pr1vbHD4Wop0oWYqlRf/5u/+Ljbg8ERy7SL1aabQFK5JOdkRry
+pMWp+i9uj8OSMz5w6VGBVMfQePGZwu/Ux8SWv33x6GuhAYOCVsW5H9i3o4OI4WT
7XUEY4atpx3l4BJRDgYnZGSwIuMsPgRuahgfYwqjANoPcpMWTPoGxyTCgzJQK/6N
nElqiMtVK2WRbvfhhmxK9bxhEY3k8B/bvJBxpFDbOJqeb2lu3NvdWzFecTdB5ykT
KP+VdQ5C/96UvLJ+IC8MWCZ7VgbKF8YGAyYky3F7Flp8maNmIrEYcgCLUjC74sGe
08CsPmRuYCrTi6PbQfDsKobqrJrwVh3fNVMCMvvoMqfE+O1XNbWJfYp501RuEVgj
TIZJEyC7YmZiAqvjqlc+0R6vbNy86ToUFnhQtaMN36RSZ3CPEpcBib9SmqER8e2q
lZNVq0W9WtDtSLnLFEWVPBt1Znpl+rB+KOlA0j6JQw1CGSx+UMMpVKxN8jOm8oMt
J85W72EclQFKF9Jv4JISAT9BHri7NaWfwml8rv/aWzppZMJ3jWZ0BY2Vz+bKAckh
mUKdDq/yHIOK+GYHFxbnlOyp8GyTM53nBEKKWl7pNgn1UyK+c13axHGXdb0hR+lT
bJ2HZrJ1vSCt8Oq2HcKN1Yuxaa/6AnY3x2W98cLobvSflnf1GH6bsDqLZsviSLcR
w1k2uFFeGhw5/o+IfqRDK0ceh9spLG1+YrzYUFHm43ZaBQaTUssZ8vNJt3ePvPUR
QGzHtabHlViPETz2Vv0YrYxvr67s3HwpEVHSXleToFjxWheXwc4ob0GhYRTcyhjn
0tSp0szvC1JA5bX1j3vdwksS1nh3CfTQiRl/QUp7w/LIf6ilKU/FQtD9LozLRJtl
dHO16mYoQMgsOkO1v8SRSNELzEZv1Ebt+UYpCmfAT2Y7m685vYyKvzuyAcaGlQTN
QDj/Lk7StzR6zib3DLLV5lgV8WsEGV6Ph6EQQ6oQjT8xh5SBrCtCNilZ/ihB5k+R
z1Xw/e79/OetxHxoYBVsKCcYrlLWWoHi3IPEBbS0X5/djX2kO0PjBXnq+/LBWIl5
GmKCdabCSK6HA35AW4Iedk6vhi8SxDfYhP4Ne9irxcuvXECbgB2AHN/1FPlsBR7v
BoI+wPQZoZZCX/lekS2eHlYp+JEwtsT2lgF3mvIwIYWn+7+uhOtDm/1ApLQqXqRK
tSmDjCIoE60XwUpcl1zY65+CLEv8vr0GGEEcvJs425HpgOUKHbxMQLLECexcBnEy
UfqXyKSfQGaMS2gBwYGsoRV/LtxlXI+aNC5OtNbAnaqPgq0jdCM6xzTTKBVEVLKg
g7J5NN8bOZrcpik4DTVjiF2/7MQ3PhAC7HYiIJH2cB5oZGDnI2jIi6w2yBUBVhod
jOgL9B+Lb070P7WCh1+beImUhp6jzhIiLdEucAbCHkIGWrR6IzyUPNCSzay5ozhM
kQxYonqQounqDekT1vt8wp+7Qme93AytO1aolXDN794xG3jEAsXiBlj1uRUoWfMu
T7dB2+w/H8JMkvLrjLCI1jMaz1Q0RCfI4ILZoxdFK47OQs9MFu+eTw5qPtXmleHl
tcLWwA7bRnlCU8K3kbvysd0CvsVOxEHHMXSU5TociZphXHWybX8+ZL6C/AsaN4jR
3MckOp+vYi1UME9YZps9OFkidCX0tniXH58YsHB9B9axOvEu0lCbt4f5Co0DI+K6
htr62EF3ZL/q/RWnFmD8walCPZMvNjyPUBsXrf2PHdpXRDFygMZ/NIhUHulnIrFN
twN3dsR8HuPRsM5TQxr5E71DRInAkg+fNJz3u2q3MgLCl4T/Xsu3dLgbDu8VgqUP
1Or7R+6G8hvO4Cso/kRb9DIEl8JnZhRpPugXsvKize2S/Orag6Uk92pQ6zfTWBTJ
lGe1YnsvEML78m49XPPoKTPi3NZOArwC1z46Y8P86fgBpUReW3UeSCvw+hu+c1P2
x1DAjzv9FBOwEHOEI+NpS3Br48rR+UkCZw0puE+IXzrKBHP4XzR8acypOUC4x1oK
wwwS9GRyUeGvUUkVy62cHhPh5RZH5+a5yAaUjeS5KxjNIIL1P58wVOMri6GZxAwZ
h4HOhkW5PSgTI6HFpkLM1GJiIB3QrQRn6GY6OSzwEo9zlb3b9foM+fukK7g3z6b6
kzcxO/725EPk2pu3YEVLE2P1Yb1nBAcMs/p8z5Ux0xOTeYGV3aVSJvTMsILGrMO0
JI1ETALWwEP9GRiZSUL+r3nRlDB7RapUzbxJXMtH4bLtCxZZM5UE699jg/Oiopys
CFYdbTG/NQMpNgSAq+GIFaJw+1+aoh4JGESJkf/FEN5XtbXwvOH+e7Tde+rlFCVS
bL3MhGAieeXSrsjrqKwmHsejYtMSPLeXs7upGs7dyjeqh5vHVsgGbKWjyNsr1Q+f
enmTAhHFY9f0Ct4x7AuPOeZ+ID4WYJhHxR6/NUJlaQGkB2r2qifzpBkEEPSVsq7d
LLdF2brYjsMw6uQSz+WYghDutw325QWb/IcQ6HCQvsZuhim9JcaDv9Zq6dD6/jJH
BPTZ7dcWSxlSRVXd9wOaKZ+zAaZkoiTCN3O1P8c0dPjvTnI9g+IfIj3IQf9mh9QX
JSIM/jvhxzQK6UcGtLJe4OKd6k4pabI8JzjqjAtpjtRcrjk5VGm7g81x+8AJcrdw
PO/kjXXBv9g9vXgHPxsc4HxD7MCK0VrWFbdnY1oj9p16xXjLWjjS01bLs3sasjhR
Q0ZdhzR0YB/yqg/vHzdmBbs7o9vB4seBOq+cOyAzbxCRxfVoYEAr/LrIBjsXxW1m
bcOSJh2r/TjVJyQBALJjVS5asoPAUHfT5Egv1yXc6ZATJoyJ3u3M+TCxNt5LsoI9
NSl3HMagctSE3QRil+z5j4BaSYkjamwhTS+eeBFiXSvVX8EQuLbXccKp2+qF8iJD
2GVn1AGl+mGSiE/QvzlBh1kFjiI03v9mB4UuNvdNbEaUFfHgOXYt14M9TMIMqhK6
b+hHIcL28+9LivaBL6BGRHO6BxF66LSHNC2KHQFekxn/TDiZZYizbvLpohYMb2cx
TZassI1tuK2p7oxRb8Ec+RBogiogrJKqMjPXf8z305oPreYCh310MxteN+xp1x34
JEOGsowejso6Bl4+XMdjCFwfgI8Dho1zOsNg5fpghFbJPYCd45ecgPMbRMMVlRsb
z3SF6Esf6y7tNSguTGBFubr00KXLq7w0rLFJj4D0dp9pOyuUDEg30d4+z/HeeRS3
y5wRTcGq26r2LHwpOjPFj/Hsr7Ugx/UK9fwQBbiMetYNboG4DC3Wcm+vQET512uQ
lkxaHVoixiu5YaF42ZDDkOrayI3trRpCphtfiQizlTTriCRj3mDnJleVAuPnij/y
oW8Td9SqVmTPZIKvVyYScM0YFwtcymX12Dkhj9ydowTWbdsZbF7IJ/qolNQsYSnR
MQGkBmWhIPnWao5K9ab4oonsKl/uSEkRh4W3VlNnI2He6goqvGZ/5gy5TepmVceu
CZCl6K1DGNPMHHhGnYrmmEGf1QzThOG7S6LQQFFxgqJVPFjU1nmfFFK49Js+l/om
w8jPyg09fYSTaNyzX/3rFNKHuaOdN1rSttLeM/5eBJQWc0Lwh2JSRHuV0GyV93SO
WfspQuBSA1ICwJBakY7UIlV3cGypEwc30pf6b8ZWC5GjWlF0NdjYzH5zZS51FgUN
c3priDzD2OUZvYwbnKoLuL5vs7IKJhWjU0dowvncwIQzaTQ8e3w6Gv/O7gAbXcqZ
f7Rpp86EqZGsmx0PDWSGVadFdFyq8fz5jEBFZPfJsBtskys7O8Tfliu/YC4r7JkR
C6ramVdzrex079qhrHdYg8N5+oV6Lc3gSGbn+IrlOJ98RBXWZE1q5wAvvWKCGHaq
MbSaa8C2L2+zfnfC9XJ9c0RWDcIvl6CRPYsQlR6OpBn47Uo0iBMlrgtyESd8okvn
C5t9DFxEHsQSVBCxVysYzUXwMQEFeWzLfwHOx//aJ5XH2xm5Tyaaa60R7llsUM31
tDqF+37Y+zEoY1aiJGJyYv8sE5N4j5ZYmhlfKEON00qpnSvEZvHqI5lg0uky+2zJ
kF08Ya/BpoSTDdIffBHg0u41gnuOoFgKD/ka/9tly4Uc8rtyFbDBXfgKhqjP7vJ8
cRP1Xef8IG0AaMQXiWJs839SQ+vaan7JyqzdT02P4+FCr74mn9s5cmXvqQe+eSLP
iSxAv34a9OE8Y909492jhXEhynT2dupyR6F4T7BADHImntn90dp/Knpgji9qyrXV
v4IemkAZd/WeOCjKyb2UygiObku60vVn+GsjDnmObwth1aF6FtG9HSK0CMLDpjGA
Et9n+wMtNvRdWxiFklRV/MCLNxF/XLE8PIJXy3mexHackuuwz/uiWKt0+3mNy+fE
4UKBt93r1kObPl7pIrYopEzq7Fs3GTLrxddZaFVLqkvOBqHk21j49VYpagAFO88+
FF6e/b4p5etY/0ssaPBAJW9QviQbDHeRRS1j1RRvR03/SF2FAC0BmlFiDFidzSfo
KKB0l3diQLvfNvTsUFUVF05sVs1v61AHS/9pZ6bz1V3Sk4j2LgQvuhz2ADxSrBz+
olBnARd4Fs3IWfPfqrFCsjSrIKU12bir06KamPmsvcRb/E51wGZL5jjDWawhppGQ
sI5NF8weNUKhbOZPK+UBl95a2N91XReFUNex55kFYxpq92EODBiy2u3ZaK3f8IAA
N1D7CE/BF5TQQCxyw7+620DSR/R5wA14EIdZ4SNLzfsjWs7SGjhXgZ7ijVBJ7vbN
JlwLXTZKxLGJkxtp7hZxpGHBwhbNxqRpk8y4Ng89TbasPlgCEmRrWD1jGuewBrin
KDrZF/OstFK5jLNDBW1iJyu8aCxXw5iy5WNHG0N4mNt76v8wMdDM4Aa1BF0nk8rh
IIoftVcOnDSs+XnbvwEw/XuS3HQX9N4MbMpeqiTZnSlKY8bLk5/f94eBxj8Y7tn7
kHnwVIUtyibwX2mpaXkFLlgqaH3SwbNXBnklwl97XhoQL/QAIT6eGGEl5z62TE9O
1tILyDQbg9FTN0o85SvVH1QdOgu4dfd1R14Ue4MPjRz4s6dGfmXJLVuiJ/H/XZNe
h/8YaeA/yHvzIoROwqIbQSS1MzKSMHt997M6R7HOB7C+33otCyVF+gHR2tDM+lfo
bdYXTnP6o4Y28ay9mSwJXhKwADPyxfl6DlbIb9zzCQCAa63/CHc6srhMKwLCtYPt
GlEib7KtF5N+7gEk7LziNYID+UOzlXwrGeGaXr1uWkcfTAem3bsJ+08RFU3IxKoG
GLNrWwDMc2o/q5G35utYMyPbxfSC6ehuovKUDbGC4J5G5jn0SsrnFmsbkeOEJ4md
z+441d77FduoNjC2e9XFcE72SswLa3NyfNgRDG22wv4KKyRYPFP6mslMDajyteQJ
n56qSB7s1lvqm9jAfJx2sgRbzXtKc10d46+45cvxtoWddL1J0SH6MEC12AVOJeZT
6NLpscYBF5If3P+TBgaN/gPbrzakRlq1UezAiBRgY+OLOSpE6CfW4bW3XSTK8BiY
7UIrpZNkoIujSKzHMqyTj0V4tIUAcEwd4T1Xhx341pssSO/XpuUCNBFXxq4cp8J7
xIrPj+VZ1wz4TW04ES5zsLHv/pmEw4+SPjgPmfXMZybJjjsSWkhHKak7qnKEpQDM
8GR/nCAs6Sf0owCvRXwjtV1l/W7ORu3WtAvJCw0wBo6pXUYKlzxPgPHOquc8deHF
cMnceOY/IhaxYIiFkONhajiuE6qgra9Nv3a5ahHRpHsu8DNeiWMMb7L6uNp9RhjH
yUl5hiZWILdXDW/xoWyRqoaZS6ESyKpgE1xjo4UFgykU++bxpA/Xe6SbwSzev4Jw
1QJqPOEBTxBMa+jo+ee3WxAmQv05V48c9gFgZIpPNALzEsLb54Bttl1aBYFkc4dY
Qna5SFxKkO3RCkonXAUA1QLmxA0/0dcobxCZzLRMGCPtjsWn+1m8UQMvQUEb5sX4
Yu2pj83SvwVKQOVsHvgim8PzH17wD4PcStVm9MfRAhwPxVc0VPxyjdb+vpecRc2L
4IZrESTFUUZKj2MUYrc/WS2hsykUdjdhh61b+KWmGViw9guGCyk07dgJmPhCqcSj
bGMyqrG+yCLCWhOsdW0bA34mNXc0Uj2qNs/ksIpE7IAUaynbNrrO4/TWQ8fnfh8/
JpvLXXAqtahcYeJxqluWThIFit9FL3GzF2qgJ8XLJHRzePIzPvKfvGiX1Qaa43ey
n8AdC/50orpIArrfUJ3TbEbvPOn/sgpgTmfPhcvSCjvLffcYUdHTC2L5MVchHR6O
u+urxhs+O24GWt12S1E/KnKQwyd2kjWlfC/aBevNXOlxUtjsMfSoFZZJ1u8R9URx
RSsSDif2ZWPOrqE+hNqDFzhIZ1vdf/KUQZM24dDpb/zSRlyldJLCZ/Jw7MbUWGRP
y7puIHAzKsFuJYZ6EgI0SbIpeO/DGHKmEHfuTQzXqs1FYHhe4M+JDor1JFQuPa7M
VZHJWZmKXNsBob/K81QX21hIY5gKXhJj5qOeyzpOBsC9d2gE643f1xYQ8X0snoLk
tygsnHGRNy1oThyZkqVmFEHM/uD/zDwSEGPZVxiOocA8/FWZOVi+Puv8xkCtbCHK
eeK88Md6CajJ/J0ttZgMjLdphTVIy6N0YZpZ1VImpXep83cEjS4AkvxzjI2NfK5Z
Gn4B1SLeijq0zVbwwz7DapoezkP2aTm3+6nbWtk66G4irecafBy71Ce5TFrAbxGa
mgdnJkFX4sxxHo5UlwjTjJ9xZycWUK3oJDTHjr2hEy8pMBJ0luwd0Kpn526I+SJV
9lqGiaOr8FM0LJruWiOLZMQRECrhBYP0gGvCbFjrEBntgLq3so7VKome+IrJy4Gc
O+SpVktW7yZYh0byldsGk3flpJMkqkCcMqvniCS40Dr2E8EAWMbu9ULd7FBXvAEz
rTJsM4uOHGMFxQW4tibCxhAwvWba/fCtnU8zKxHmHFTN17GegXZZhbK/CdAWVDDZ
x0N0XzSGbLh/ribh1ZPBWYWBqFbtcFYriA4dPDBRpnrZRniZY1oxQ/sRKrtCdIUS
0ZjfYDd0sGDgud2cp1q9CewOZ094b0wD22A9TkapVsLbzPt7Zul3TcBTXio16OWT
fslMcRWVjI3C/MWDhMInCpeE8zfNB/lx/vw2tLap6MZ4QtG+DdCLaQdnEfa3OT7C
15hJ4DzAI5fd+VMmOd1Kq8/GFmh5Ej3I2YtjFfSuAUAEsM3vFvbzvy2VBkAehhX/
q35e30r/WRuyA2uSNgz3tJwzhoX9/9yumGP2wlfVfxfGBMG7bC3PFsI+HrFim/ck
bKZKDgl21s2dbpyOTxQ3kuQ/aQJN8GfD0AI+Yz2pJo+r1y4PK5iCaBvDbwTxJdNa
8bCcVaKPMowLzfZZLzAUqe57wU//8emrYuKUylXCbGPdxfbT88paeYcYd9B1poAV
yvvfTf1DnPS4tffUdvKlmI48cVkBGwY5+lASGBWuTTvaEsjqhK7z98Qe/d6NPL9T
69K4Z2YL/uYCkZ8VKPDLVTMHudhhLQkuoufUVdreznjDT0uiL9wWFE5wtcDWC7kq
o1MGz9xpC/D02hlVF5XAGF3uwf2EvO4rY/Ko/9cM6xJmUzHLVgFn8QBeyjP1kIrV
NT0k2kZDEf40i7QyMMYdcaIaV+lHiQpD//HsXZVLvTrtoOAcV3f5XH9gfyqNj0E5
uBfvgli1UG147C5bvhiCcjQIve23khpul8n59IykM1Ia8gbjjZ8oKCzM5mAu9/xe
vx4ypU2rj3nTwu0ydEqceNqH2Z3aWP1qnId86cyh8/xnHywj3sC8egczZJZdoF4c
+OHrhIf0vdPwGmHXXd5uoOQzXPAoOXFL1QnBiIkAmsDhQcvJ4Az1EgWCoAxBotYM
n+/BRBAfcRNIkG+LDGUYcfXUX3wcTT+fZgJkAqMDV4WG4hVFFCWtPnC0DNdhNZLm
AtNItIk5jhcDKC6+yWtCqwbERHQQNT1tfBVw1qd5o1au02smzwcQrWXJOj2SxmY6
l43JdTPK+gGayn9nTbNgfrV9A6nyadcydZr+xiCPnFJi9FGtTemb1k81k+bAm+Cm
L3VtGdzWs9Z4LWLf8a66oclwGddlKJ13GxPJiTEfXdb2sATAydphX5v4zKj2Puy6
/i4GxIHSBTK2URwQQC1GHJPB3nJr4UaPO/USp/TmCKvJ64a19M0/agljhAzfx73M
x6R2d68/ZUAvy8xF/Kjz8Q==
`protect END_PROTECTED

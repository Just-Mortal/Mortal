`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0HRcr5hUR7woyxx1qz/hAoQX375x92J/gaZx45A3d+N9Ak/znKLSbIvHp/w4iC/c
WMcSiqKnL+eTd7wNerV/k8ljfs2AbetcEYL7h3lPy1zBkMrULkD3g+hF+7VMXCTS
w3+kws57HIAcPjuD1hTHINC88TlhUK00hRammIIeMu2Tt0VLgfJYXdbL1sp00wKC
1828GnyxkVO+HHWol/CttL/Ac5/aHpKl4jh3ft6EBic9IKS8Fhox6+2Uysm1AnD8
/epK9jufvbiv50gaw55XyvXZnwpFXJ+LLfXaUxVApFew4sMqEvGg1YgSDpJfrDA5
HIrzJSVhLDGlX6NKLcVdHAsBqnhl1LPMIErmCAaUErhOURBHc9QgHGIYJabNKI0t
G/LxUAGvp+W1qaiGr9X6eZmAF7N6DLtjoSn7HtVqMFupI57gncn6CpSdGhJ2gf9r
FmTGX0utpJBT/tdgAX2oM5u/cf/8f/ntIk+jNFDzoyiM0eOZOYgW+kl1yRLyo8Lf
nFGKThCKjhyYaIKMufytVIxzTQgi0YHWmybeaEJkfVv4XzDkZJNVHeTJOLyn8L7I
ZX6MipePg0/uFL8rXubg0m089tXwMkYnEeD6g6IMi/xKbxILJguX8MlPO3lg6XSl
W3GMGPUZUiaxs/Q5baAWIowbkEj0LyxVXvFAMkVrELKb9hvs8go1wZoJ0jjAK3yL
u9CYa5ZZRli81MmjzEtbEM0kzgdJ/GYV2QnsnnIOGcivn4c1CmN0q3C/3cPB28lo
/5yfjBMtV7uZ/YH0AWhMzn1Mx3+B0kODF84mDVHTPacST948yxfvmERESn8x7Lpg
FX8sjH/ArC/wPY/MkKyFdp6k0129QhMNbZj+oaBcBCcmnMy4bkSNcArepkRs0Qia
uHNXiEezCTFFqB+CeZov9I4jivNNDFgTgvvQtWg+/7sokecwvQM92YeEFmVFKUCe
8KHTtNY/XvyrHkhZNbz3RTZ/xZUwsIy2YSdwejlm6sFAiVShJgTslUTDi7v1LO1R
+C5HcDD6TxHsPBxdM3+bxZPnouZRXD9E59ZweZCb7dJphHcoKxvjKCa1Rslab4Qp
Bhi6jWqyY7p3KOs/JWHjJpwo3ZVAedlEgcV8V+kFazbzMR43OMsOK++bL+CqDRNT
fFNFfQFJu8FIFmRfOJ7so5iSFwKGkEtFBpmHKSSypFbTV77dQ5s2Nr3LZ4vnXdG8
BvdgoBzYmM9z6svHqHVt0r2WYWg6AUXEV4McCtJGvYj3S4SMLNUKYU0p7Iilat9V
Ce0Fy/qxLYCZh8J6CU61m3j60crPrmSsfJ9zg2QyDffb6zb6xEl1Wz+GeqdB+hgQ
BFc97fASRVVZ4H1OGYyjEUwODxndzje4YBxMT2KmTcUr9DVQ+gv6782DCyvhj5V5
+uDF62coh1TyHjyZoL9K6YpAeGCZbvQR6If2CengnEjcrVIekbklFta9vdq7oPXz
P3APssQjkEGXQ/u5DKGXAQ1u+nmVdjVk/bY9nIiTlJdbyqc1Mv4PEWZhmgQijdbL
RdxBygc51+zRjqX9Y28z7NIL9s/BLsnBNKd7y9x1MqANPMNsFXDtt6VM+K/R/8Jo
vlzU67xKJmzbVpmETjqqlVgXrdV1Mhrp5mpw+E5hGKD3hS0oZHtUJ8V4FFZVyS/m
wpxExBSi8WOoXjSKk4eav5Ggb3Gy4vK13N2dbCzMewjfA2LEYyUQ/q+5qyeWtJz8
H6dp6cgLe8hh5RNGiKkCRDy57yB1qfrsUslGz99P/RYrKdA5e8Kw0J5awdrZhuVP
TQ7PQg9foK3ryoAw0KVBbIXGVINvxHvsAgLxUwuWLUHZJcGnG7L0dleg8+7UD6hW
9sK7i4WC9iliXYXbjFlGfnWcVJVD8Uy+Z1F9klkNR72p75HuTMO2ZtlNMObh237Z
cUp9y5LbPBxqECpcYShCPLdUiam004k6Eqyd27cOaYa5p/LbE43r6ugR+pyWHuDd
XNRzVMDBWpUOq3HFrDfPHf2lMToN4U53dmOJaWbRCMvJR4jKkPtazvgpW/mXBxDY
OC3nFVgUxOtDaMnAxObbiH49PnOvjhIXSOAZrp6rJbhMZowYaJf/j+eCAXYDEEqT
30c/wMNPk7ZQPmlnHvV5KSs5iLv287oBPXKSNX2lu2dpnnnqlr/Xiv8f2uqDvfbC
FV03G79YJJ5lxXRcNTWWjFeV6n5dNtegtj84jLGzZw+DcPk2n2pMVhcBh7uyMi5C
DciW27bDEAreasU/Tbup0l5zKAfiRQBa5GKedaHc/aYtL1kBVaIYWaoAk7InbtY5
vDO5UUUQU6qOJ+QIT53lGPgI0Kopn1CMnLTeyMsKvQrPEOiYi8XkTzOFLIbWygBZ
hebnrPsfjPBfDB/6pvZJMbiivMuW6P4Axj2G1E+ZlShU+Eifh1eTf0fTKZ2toKtE
rf54bkK0KQ2BTuUxojbpwJun0P5gOZc/Es0sOofGiIRgBowc00e2GgrabCEaq7o3
nwYE71zzbrHxyPIjhyIyvdZdM+Zwk3W3iZdWi1kI5JmDhGNVNfqiV7tLffEH4Zud
Bs2VbxaOxnp5sdYNwDYCWmA8WK6lupXO8VlDcJLLJX+qfaBdYawiFfhjgu5Vwg6O
sKwNprm8FwlBghu5sNZoN0VZU5//9h29sMdyz1hJhhComRVoIV+vdytA9LduHlqY
6DA45hu+PVtjwv4oiazo7QswLOZI7RYnfNiEzJ/6tWa9mBV1Tvh5ReCKcDTgqENS
kW1gysZ1lNn8+Ibt266FsvBBkbbFq0yx3eKD0FbI9595yHI58fqyZGtZSLiY/0f1
YRwcs1kS/9SWP8q12fBnQ885r6zn0umCP3AzhsX82Y71jk6Va1X4BPcQ5ykgxCZ4
7dv3Ywwa/CQFWja5m6L12tTBVmKcEaWutnrWXb1Fye5I4IC/2QrxPRTWvt6+f6xk
q3eOYCVc0fWegR/TmdT+1gFfuSrjn05IILw+ECh79KiQSsyQE27GMYccaDxPr2Zv
AnA1i8w+hJCGLho2UJAmpCze8HL2/15EpTUt48/5GukEWBl2l8XRd11fJMKBejTQ
qsuu6mjuwtNF5J09s/NX5cZVyC9QEbLt/s+T6jzSzfl+wsJUvAl5kyxj4QuADMnC
qCGDhntS/A/7ILdv7fu8KhcWsQ2mkmAA5aQGdEBqABnKXMmbAOyrk7lQcYHyMIqJ
7MNn4CRequ4QtxvZupbpffi/HbN/9LedP10vN6j2h35LFdDE4nqDtp6Redu5hjWE
y7noRoR0oEWpP3qsp+4HBH0ok7tRtQq4llzs40yLdOavMm/a4YEmMY8vNPTieKX8
ExfqGmBHFj8c1vvpnxPvoOR5QNCMnSaGcP4qjI/Ox1Hmu/dM/CFBY7+/ClPlg34a
nDe1PW1Tv0jHQIu5B96lx86jSd0RzvRHKXX988qyVKxwi/T5zRGeq4MxyLXOYfyB
4mm/6OtlLcQn3fBUR2OXg1vWC8NiLR3FTdpBjWbxF0/Olx6ZrZZ5XtVwnjR7Np1V
Rpihg/vS8JpWO2LChLICx07F25bzg6lq/TFxYFU8VO/4ctgrZ5gAn+y6rbIw3cKM
BlPfg0Xxxx+ftNJadsLtA4lY+THXnZs9mSPnllMWt9kNGS3Y2Je8e1XpgOzCF9qy
/g0ryGGN/QfNP3IFQ12HgvmAGHU9S972UbYEvaJ0EuTQzJvd36Ho7AWNGnSVrXrl
uf7b5sKxKokjbYxuX9t7sI/mORJsplI0qejPZxpOiJbOMkFVH6OJcIjOZ+h5xT2y
JcQjBqb2nRJaNYkC+huLIo6+ZpYagBKvYE/YUHqavArPzWd3w2YJ0H7stKKy5cSH
qsmBtTP0pojufte8RvfrAg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0e7f7tPBhKG8WOYaGiCvR3JBnDUBG3HjrhN+luaKoelBMlJrpXhRWQ2OciyyisqL
jcSUxbXxZZSC3cQ6e9nh7fH8KE3BWz2d+whWblxGXZ8EempdqioL1K5xBhMm/l0W
C89S6ySaPK6I2856O9kWKhYkt3OYOL75RoxjB4VLRYflnCIJzWgzgbRc4xYzu58R
D24TMV+UYP6a+oy5Cvv92V638d4CtGT7kUPITbP0kDPdEejKa3CJ/ENGHORF2/dn
vlDOyQ+3jQ5BK37j1oGQeWvxbZCUMrx1ElIc5hja6rpE52ykIIck7DdFx1548lMz
qsgJUlEvAozKAQxIjMZYpHddkshNWrrEpxGf+QBMJYSvmwcG4DXHg9loE1Aj2bnY
EMKh8CQRCmwPyNAFYJORAmcxLSzKewyfKU3xI4jOEkT3v/tvzM85aCHpzfkM6701
NYhf8Ob8iRQjqfR7LM3qPNiywjUhw4i1pa6NzbSurvBHu2/cijB9RNFN82L7bzjr
fCDmNCK1FrsxjsL/xldTRUqjNltxBeYXTYP7oepFz803OTigECVTPjIb537y/SQz
oW+CZpXGttD7jSrD8l7/8/4nWQqEva7myoyCqNw/vAC/LKqORPoA042ZUYWlrYDl
xPEphR39MiJuXnABfzOuj7mfX6BNti9+N3UKwuBIlrsnFai6y7JkydlANmTcE5vB
YTi6ijLlFa5ozxZ3G/FbHjtnlD4eDOO/TKAgyJR0A60D0br5V5wzOHs0LPjDnV/2
JvLX+45KhTwfnEO7Fq2tjiGI2xmkB3vLDaCwuUxKOt1pStoQ1SWo0PoH1BtxeG3N
YdSwC56YGyvwC9A6MQFvB83AYP805LSmxZnmgsu4xI2es+NbgCGQYUo+lCkRlG4k
CcpO6UIGQJC+8qk6FY3UgrQHH59nmM7JCuH+gEwSVgkNI8CL39Sbx33w3VBPkKi5
nlOLHsc4j37PpJ627DOutOKRykTbczJtc5fRjm07auyyHE31/BFax+xMbZyVHV0s
jKVgsnIGZjXUB/sEKlMCgz9YcvXR5I2i82vZPj96nn7FbgL7JJLsXTuuR/Q3nzol
a2Y9mUzD1XMYRGZOeFQJfhzc62yiGmRbcIdjP4aNwY1L0JDQX6djITwyp0ls4bXW
4lqT8p4ZfK9H+AbhpuTmoB+Oa9v1zaWPFxNK10k2fSETSVITdGGoQ2Yctidp6V+d
kFHbWquec7lb+upvh2NxEA7aY2lggI7XEvRNAqgHJzXs47Go5cP06gWgQwDe2aNa
ImP5YGcYLt1GloN7Z+AeRumRiUsSMIh5a0Q/XwC5pkz8ADgK9JLSl2kJPRA4Utto
DKOHz7YCOHFpXJ7bdj7O67UdayF9z2Y20A5zluQTFxVbJFUGQM+aG7VeWXzy5U4E
rLA12RqHRwlFKeIeB4cnhZe4e9tpfured0K69fC21NH02SvZO9DZU1oPJLPZ4740
lcn4Ty6jU2w5mSWLKV4IKqpD2e6P69z2FF3mBGzvP3KKyONTLnTFgSmlWvbraHjb
nkRvzCEQee3ahpM9YRFXGeL8wDGDDKfZtQTs3vvrIggSDAU0ANEpx73IXMzlj0hn
yv67qUfOADco1N6HoMty+1WkrmChXYuWdM0hlDY+gc1inEa1n0ZMHflq/+DFMtYg
8EtkfcY4Qd0M+alyjhKdBM3MH9Ebw7Jmst0ghZlippNxbASLKMvz+kiazdvv5Xmo
PB4GaK3hOpMzad3Y5HerUM/esRR+xumUV0xOXfLZdsqw/gnReTglc7T4xvfaPbj0
Cz8JGmrEwz/rmiGfwEGt3W3oBaj6FjBua3hISFdYO9PSFW7feGQ9UkLYtI9EpsGo
806J5iD6SEidl28arLzjewnqS/FT5OhMSNivU+NhAVuzOJs2jdnmHGnxOR64HgJe
rG+OF78U4y4wcjQyUMjewKMuQH2Y5+qt4weUk/PcXlyD7SZpbnMI/JGEQUENl71o
/+9r39GzKsEoPaqd3bvY1Zl0FzjFocl7/IHBfISnrvvpsGNjOtI7fzVFw3Lb4zOL
zaZkj0uYc2tLvR0dI9ZkSH+5yy8fcf2kDgMFMJMeHNtjquaTKU9VBgzkXZNFZkTU
+2iFMa7NXQe5IZe11RaXCrJYgp5agDyi3Kaeg2mA4pSp3TBjt6+U9JXCSJBFZLO4
UTqPURU3N80hZIbEM04LMPvYtiLQxQvwBHtEmqlIhsZ01qakWpmH0sD14KK9ACAF
Ea/B6Ex1iNeIQW6T+sfls2jIX8cYWD6Maj2kMvN289Q05KC8Ph0C6Bq49gqS+7RM
K6Ns70Z7QobDbJ215Of7p1sBlTDo5TplBonhN/C6ZtyFK4EDF/xkc/Erp95juwYi
jUWfBftNBQQtlJzg+nyNOmhjKdNczod/9HhK+7+yqbeT44zVIMHeQP0UDMNIt1IQ
5DOmuYIpmBnOxWgmCdAv8XiD7U4KTzOL3MJyHBsS/FBBOuxYYXt8A/SUfqShFn1e
XhR6toJvq/8bVtTr34UHGbO+CI7Afp4vgO4RXxXWoezIwGNseTartpvMmOSb4K+m
kdmhxqq7rnTBWbSkGlL4n22wcjpw4qTZBrjjM5Arg4WXxHUIYRX3B1q+2nSy8TFM
IEx7vzxK+MFOvtjR438D0Rr88XrhFkaOpZDafvHg9p0jP0iPuQuRv0/IQ3EsysB6
zqbpfQMkc40ohveuTEZRwUNs0zIPQTOsQPbaw1+mvuKPeO6H2BjvsLB24ug3jDym
/QF3DeSEl48dBgb/XT3x4D4tuUzV3qpbMM4PKhx1YQPfhLKoBp155h9BAcFUGhx3
B/7YQYbrR6mH9ID43TusWRGE/bgw+op/5ccigNBmN66IZbnarCAF9mqBcZZc1+by
AwWLS2NOBaTlQHtxcMEvbLpQYqSEusbQF2gRiIIZGVRkwAY9Qp26a/wBgzhDlI9C
fHVrojik1MMxX2I9oNFQlP5U2BJ8k1TPDTJb+k86u9eC7XfOcwNsRdl9FigyuxbI
YIJUe0jpjYQdoqJRStvxF7XEkl5w94Bph4m13l58lbZ03qJGjc/zyNJ4mtXr5y9c
fXA4Q90SChG05WyMTJODDAOmZQ3D52YkArNiZqPdFLXSz5utoborjvhvCT86ATRA
Sbh5+T8rsL8/82sSWn1K9zzMur/xM1sCEH7VSxnaEcN6Eih9ZQAVkQZNmkXs5HwT
sAx1KrK/lOXQfJtIw8R2urycxI7XPCFzkYMmqogjreIYaFE6Wo+Lss9wno0U0KjF
JgpxtE6VHFhKfojab68dbDlnFhTDWz+YSWJMenZwW/kM9132WsHzCfubGNyRIuvr
uvUamKBvl36zzmG04DuWJJqe+e9alMRUm6SBXatTQmdKXK0NajYdMuFuOiKqrRzX
Pv2vNu86IHz2HsZ8po3mCW7YP9lWGMIpezte8jSYSmwRDPGZE+VR18NdhkFImEv0
L7Jziboph41A//7NfrVAMonvvmKRc1eKBhnQM7e/kPssGQC7a5kmrk4IApO5I7Hy
54Xyt8vNmxiUmaPdmCJrDSMQd9KQcM8usDS1yPAu2TJM5Mstwgo4nSG4LqzrSLK4
LZUZsb/dTatogfSfB1gdWETPZ1LUIoc+I7U7/RPSJe+UvngmDzXFW/rONi6ctzVW
h4PYQXltX0WvtkyWuD8c0e2TsfGPMrIeyY2tNybOLKDM0FtiS/d3hTSB3x0kgCvS
FMLXks3cuKBPqVZPBwzuYf9AHLPryN3YVL0PaeYwO4D8b6g5EOjR+WwXq4xhJHCv
k1tHBK6uvIqY36m8yd/0bXjBBNwoVGrEwQuKHqo6rwahsgjsiz//hXlpGC0ETf0y
ZjvTPyO75vtY+D7XtmylZCdBor89PYD2jrISeYzKXsp6WsTJL6Py93qmf9FIyCyO
vdWVGfaCaW0paeH8e36Eqo+ebMoK9KeOy/iF6dcaafgguAQnhIBGr5W9KrTt//JP
Su1eZPJ2paO24h2UqJgiWH0jp1NjzdH6M2WrNh+xAXUR5fJtMDsrxZOQmMyfCVQf
BMBV5ztGQVQlyQ0+wZrRSEpQB6SPidj343iILMuY8xFrs3j6mDNgFVUm6Wz896dS
nq6s8jzeL0IFy6133TljQ/WQlnbIeglj4CfcuJn6jNc3uI6Dpgpxt7pxxlq6f5DF
zOejZ6go5Nb81DbhHKQtUW4s/AeAfad6qO+HClV6HfQZcogNEIDbmXRqKbn36Unj
9Pjx7DAKXzI77pETW5woado9LJaFiX8StgfrnncM6HSziRigZMu7JhNgISWikwEb
HpjDRjvygawRbsc8dlih5GVMUDmU2rhEOB6kZswuutCDE3ffXLTrgeFDymfJ6zDh
1ih/Jmcs+q3B5RV6lirgNxdMGWrAY0YR5GO59FeBxv3JEtUUp/zUi/zzhgL/FFDV
W/RwI26JthTHPv+2tRTaBegwuX+vgFjWGe4384+eEpzUoRHB3fpuYvIOeM7Met7i
EEC552v47huHkVSE9iPmA/Umm27Pj4DlklAVSymNj5/tAyy26w61uQK2hGibVZGn
VSBoF0yU60lXa2jGd+rYTYwR5OGncqgHhbLuC7r6MVLmUiznFqFoZwkAXVnjNg8E
HQHU4pargGWupSC6RTECGgsxaCf97QbO4iOIk+tDwaauCaVQdWKqN4QFEojeO3VQ
FkgkWsXJeaYvQAsQ2Eq/VOkf+HKGkURhQAQ/9IwHohQHKkj5mSAGQ5+WrPtAzTtP
f3uwj6yw6yL3kS/C5S0exFe/GwoFhYCgt3pRWjwOI8OTC0/eObX2T/m4ofyIzaYf
vrTy830acFi3GRMuU9X+za+DIw9esMK4+vsmBhxv2NbFuGB4Chq2xp877RyVS+jR
lPmGIGlp4Cgz50h0De5aoPLQPqHERTnrXBi+rSa6KUNufb7IgerEO1CKZRZur/Ia
HsMlOcVLr90j4Gp3RXUWxnQa3i3MExcU8W+OBcXpKXQUUOdsR2QeTiLBTRSd4H2L
qPcfxpws4jhTDXHQLH9I+diFBDC+pvFjOtA4C12tNL9xdatyu+mmyffZeUDVyjrz
wGNvNeamPhVf3zHoGHa+6VhStIHqklGNkn9pz5yUTTkUlPkUWWoiiKjHkvYSvn7i
aSG2Zn9pULu3qA794JLBGXrqwv0xck1QiQUyXS8nwOW+F2Cmlcq0s/606fA9/U5D
9+tPuoysykr5gYb4o0XzHPadwo6iZMVoPj6eNuRpUQ5E4vO2lXBj2GnPcgt8zrMQ
pl/6wicPbbADAJPE9FWnEBtz17gU9XqlWzggtIuO19MrjudWmaF2xPx+EH0fkUpQ
0hLKUcnns5ZkHhEQqXLsluR+vnEFZOg3gDkVXsMWgcUKzaxSBWT8yZf7XFPrgsGV
MWBuBbkMJ/npMydkZASRensKkg+oNmOd7/X80yD3iTfLrhLddqIqrKL9YtUgGwu0
qLL+uel3DfS6JYEHCcIS12NshjiUtxY1ub3qLLiigOaxQ/XsQttYlxMpoTKLJscr
A684xG7M03GxS7yPsVSghEpmw1oOfBbD5IfSAStfkR3gy3zfQi84XwL1dTN09P3l
MHCl62OfDrmLTN20j1z7h3mmfUkjanJVzVG76psM+J+ixbSSji7vBqY/n/L5c7Hx
o+xo3K1XofWDPALNdbMIRdh2vkPojLoUnbGHO3FJ4MGyvFbaCge3Nogw/TU7ot3D
Y6dzMKc9Ozwlz6hSGqwseGUaQ7OROAmKLRZ+0pO7yqFb+JqHEbvcXjE3dKGH0Xt5
RV86khxOKJtXUmgsYBaV7wThu7NRtMHSUGEZ4BLHNgsyqXmXfznzkoMlOiRko3WE
9q+1V6KiH+rUsI4hHsSvVzXtHJgYM3c63N5jUzJxXmzXodnokQqp8yGmPIuGN982
t19Ps8l8y5asbhqAwXhhn8NfrkJ2JqsRfrMlWVqQSbRfqkna8Ctr0JwzWjsXHhn7
VxWAvRAdODBO7x0GuHT+lMrEB5bO9cFltxDOg67NTqy0fPSe7ql0OZBYUcjBLzoz
XZtnjNJSSDZfEbHbhvzqsV9Fj7Sq9XEaKIGIenfSqkjTrVRECG9rpI9vGybdd01v
XvFipO73lC/DVkMfjSzr56QMUXek7EpHUTS8Q2Q/kPRkejdFWvxyPKZ3hSEajko/
m5nCKzUBUJ2IFOW8Ycv92I1IMT4a46Jz1FZrb39g/ndyoqRwP04wnPk9LrrdVbRe
Raq/oNmrQ4n6//71CJvFXKpBuiC51Tf88zi4wvTCOiJiyhfsQIA+SRsePn5+VmWo
ycW32dadlFQM9r4CAHVYhhv3meplwc/8bfPhMwsSvKH+AydEFXVtAhY9itOvOzxq
Wrmy3r0qGZ8R2rfVBM7XPvBLO+v36Di5kk5fPNKYtB9V+1+edYMOUXyB+DLw1EMv
ncxIkJur1DJJVw+bPLJLYteQtMCEFdk/EqQWFVp6gB+1mSJPhco8hQLGjLJkr4Lv
Un9Wfd3vu4kCuWxeBIyPtxTQQod2PgcT6plYwFO9v2Ycaf6pbBzvr2AdeDPOF9vk
dSK5bHQd6M7EKxOYvtLN56Ssz3LRL/x5z1J1LU0zs8s8gEV8qd5kMneBVFE0ming
ff8n3dWL5xecdvI0Ct3UMFxTrAQRar8HDEzfEKk27RmWFHQOYfBXliKU0LRstTnY
M1N/M7TqfxNWntLN1r9zs1PAO9t5Em+WucjsMt+NKeweCA8rrGX4yg2SA81leK9n
KGxZJWCxEHfnEIxBr66J/HOgU+lMT99bj5q+3elXFbyBCdQ8Gn/mW03P9pta8icj
LY0VY9CLQyio3Qv36Rw5Rcm8xh4uNuqaAu6j+UUQLU1py5q60gw9WVSJemWSrCpi
0BekPJd9mV4OAqxgGXwYnOQWaSxa0ZkWvt8weqidngOOqd1TJ2Xc6Ttx24o++Cu0
CbNgL/YrTxc+1/Q7FzC8LWBPRJWzw+wluweUbOTe5sLifqZ6HyBduJFU9oIOzl1Z
18MrvKt7U8sqGtQ9F29G12shrpBCSJyKmOMqZ6uho8/2SBGFTU2j9I4/OYP441cN
JybQPZFnoiUsAgWCHqHy7HPJthLSGsr6zA5P8qNuzlYHyNo3Fz1yjnZseQbJikbq
msUuzMqXiku2Z6JAE/6wJLEsq0n1VbQpv2+QbpgaCO177hnAMBsTR0ljD9lDmNh+
IFc7UKoPQZBespfkD45LRmUaz0AIhiHLEZTRgIS7xPoC+VAVYp3faXG0TX/KpRFz
v7JhvzA3lPJ1v19E7nB72cEBC7Q1X5ybAz4ZWO0v6gbfp8T71PqMW9n4smdy0whq
95aUukPO4vnCw19/TbkaLtpr/a+MudLoodO0jgGvFSGQPACkQMVnSgSK+sVJ0+vO
0jSsB/0Xh5PnLh/Jvo4QMbz7gFqvIx1hwy1dSKAALwTV1ZW+Qns8VUYGO0cFi178
MCpY6dRshqxcpQ63hd/vyXLOHLv2qZsr3IVZKUuV8/BUOCYRpNro94Ti52MB5Z6E
X4gi8amk2WKAZLVt2vJ86tcWko8tfEh80jZPg830DwgjdEc/6/RY24vovfi6YuM9
us4FzJyP2mI8/MaMq/ZGnDCFcacp025ba1NvXXXr+QthWmNmLFsemmyz9+ri4jTA
tw1T1XrhtQAxD60DJWLVbZpkWGk0n96WL/3x7yG3rqMggKczwlI7rv5oMZF/9vnt
J00B58caDzqcGYfegE56yk9sF7LEeJgpTLG3SvJ+f8QXLUQS/xp0Xz3T5jfph/TM
nelH4CsfYr+h747XBwO/V8xvNI2GCAU7U/bMp3yzTS3pCN61HuXpkAJBEax5Y/RT
+HAJkz26+xatxQt0x5NzXRE9lX3AOqEzP5CK9/x582LeGCUptqttdK3tsKUO+/KL
f8lyYzTPhpNRoFDErw782PMcPtJj/aoKKdIbQLiQ+86tBm4BQvK5+Ctvu/DIO9E+
W7kkzIor2uWC4Rtult+iMbwtOMlhBUvudEVQ101EiwQYX+QLd5yjHXhWnNZZaaFa
cDngkEZDQINf5v7VMX15qSzwBN0xxLgn5WVjA/B/JCGgzrKUUoeLX/f5zR5NCOtg
vZvhGmRFO+gOGkG02eM0F5r3CaKJkCSupKQjijJ8zJV13P7otdLYkzUuVqIlRwaz
9sAE0YDYAUOhsixVEgRZn5wTgb/7PvYIAEpmE+DclAc=
`protect END_PROTECTED

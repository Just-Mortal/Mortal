`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p/AsmnPM0NHKOwvI6i40lvfr+NA1nAvkXHxopoLXoJzrG4mOhwtW6+ReBgN1aGc5
wgNuUypoRBRNcevpFTuY2U0399hRVNTvqlv7SfXAiu3D/1bJAtTQDxzlaZtPdYOS
Jc70JNB9EM0qKcNtjE7B8w9wXhrhbzrusV4Emx8HukfF7GVKw7OCS7dUG9Xxr5NA
rdw6rQW+tWUcJd5ijKdFBmKEhArrin9pyaFR+If4GgrYkb0giN2IJGZIBCftg3Ho
TU6hecMWNyoslOgG7YftcqRQrh7pRLpWGr4XXm2hjO79+PGYoi0jrcrnjJirYSw4
tUJI3x85PsCtv5uk0pJrqZlaWPumsUYuiB0RsyWVGXwkzwElksah4bTbA4asvIVz
npvzZi+z2W/YGhH3utB6ur0R2eHBP4VmcmfCeQz/pd2vj9xfAqHEdyqTQ2mIdDQ6
jfQimOplmxah9ACWlqoSI9j4en3+gBh6qesCWAH41iy43qQfsiFEmDVbpPACh5sL
vMOxvTYVKzy/pfxLb7VFOsrrZPf6oqGOhVpM1k+EOmcPU3WuiIHSXvm1JP+O0Xfc
Vl8AeDrfgQS5nrRbkb5ApX6U3G0pkR1+uSjsT61bJQN9Pu/m9Wl1CkvcnNcUTaKo
/YeQVyuyuco4m1/UrDl7KIEE0sVVPMzg185ODSq3s7Uj+DbZH5e8nBHQtYTElWS1
iMFYY3RrRY2C3q4zlC/CO+8t/Zn7n85tffOFM5z3bvaOV30IUIBzzBfu9yjAMhRs
zb4wcNDSeW+c7jzjcMFT4EDyellpRFJ1tLFT2MNQUX0O9jRc2zzKmtOYlLZHDiIf
FYAnl7ab0jEyq8XXJ8Ozz9Wwy+rT8q731TGrJwLL+KAdvN2SvvGbKMP3OX+0qMFO
JBJobwHQgTV2wjWY+79qtyhWdHxGZISxCa+Q4ZEtn1owAHovyAzh3vGgAujjVtY7
emScdrKOMDo6wH+ebSfmAkZ4peitVFiY2SBizkzasVfmqFE8ZFZNiYw3tzKrTcyL
bxIe/SOiTCzF10M+3S4pkaLNecIdAiaxdmbqoZQFHJkRJeOw30zn5cWyr1Vo7ndH
`protect END_PROTECTED

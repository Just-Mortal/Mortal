`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BArvwlNG3RpRolGN/fDntsYOgby2gzP9WCwcRvAvke2CVMXK5MnFreUTZ7tZ0f//
7MiawkdBZOiwfWSCNzuaKncaQbbwhwEDf7sgWMhJe2GvMG3a06YOqMTv+T9gLuMj
4eWUERLAucwv9XtKQwetuF7ZAuwlJxyFPTICnr/HyeQIpzlmV2oOZtJTONIC8uZ6
Nk3kUfMfMar0DZ9vC9UyX0couyOQu/apxc2rmurfkqWJTKUhnhcCgYwx5Jdgi8Ca
xZtURlzaqr49/XCyGa9Q3REk5rbhAQ5lBwMPd0DKkS9+ZvyFr9fmNF7HUF/p1sk9
xIGHlGnJKjNqJ0HA0xNPQFZHNMnkB1cPeo7ojd7CMFWCKj2Uf+pAAOLz4UwO9JhW
pgizotgSAaACZXjjZbDKmbCV9XgOR1oZnlC1E3vCJzBbuwRB3TyFi3jRJJet7Zyr
hSxTGekAxVHtChtmyBUWQCulaluHuKqRjjY283sc3s+9yLRPXbxjkdoCoiBxP5k6
5GW0RBdgV2I+NXoADZLCMFpwT1CpELEafyXIZgj6x8npqSKDpv9OzLw1TpX6GCj+
XBYqj9PrdAh9fdM5Uu+z8nRfmQU2RfKeveHsvpV0T4fktFlN0BPGiytYciueP7Nz
aP4wCH95oYKr6hXC9DmztBCwqNJnqurGn/63jkGDAbGLIbkYHLeoWeXKHFyRi2AN
rfhO8WmUXzZTiZDTV8aL7k76ljEZwdZ60oJRicw4YskO0NVN59zQyH2gD+/YBH9C
W+nTDhkGYxPieY9+jx/mW+Z595tPAeSfgliyYv/pMwQh6QyeaKpjtsQNEL8dtJ5k
zxlpdqxS5qN+h4yCaP79k6zIBHbUOBkOUsInCTpqyGVqI9wATB0hS60EIjRZEgYD
tsg3GQfNSQQbuLMfjLUNpJoAZQqOs598s4o9es39bYs22UWAbWQZr4EesVijDOyt
jagy1nd5q4nNDPfcBg35iFsbVpcI3vIdrGCCE/QCxfTboekEhHkQcE20R4kjarEX
jQtWg2Na2fUneHIYYQR07PyKqExytiBZQo+Er3z/KFKp8Y64AgFg/8RJZzbYwady
gN8wwa2CFmb2axiVYgy99z3wc2JXLJUN98N52Io3n2o0YZdscXm5HXaB55wf4ENM
AkoSuNKPcGJbuR6ucN9Jzfted7yaf577FG2TIA/Qkq+k9XQ8cjJNy01ObYf0KtMC
qfsr+f3K5sWmFl1gX9Zf5APBYkWY15CeGB5wMJ3AyNT/bN9JQwcFwGbQ9wjrzV5u
W6J6KHhs9j4uw+sl+eDzlM5f9AgprrQZz+poam/VSTEAESSqivTvIPoqECiELJHR
CwXR/6Pw1IUyuSeggyPBp+f5c0ErC6yxDfad1M1sbqW1/iQnL2y3oTVJnQU1FFnq
3/9Vm5wzYiNY96aHT4aqcl+fIcEe7QygLMuaZFVuL5KNaAVqrF/C3CpNJK1T1f8j
PrEWIQuwJqLxiH2U1CQIjC2CwL8YYsAfeyK9Knt+xECbXazNoutQR/wJxj4CEmsD
lSXNfLp0mtHnqxET0EV4gJMjm4/QKw7OSlLXzF8B6rPFi5PGa22LcPeXASfOCBv9
btTWmlugjgVw431M+LROnCpXBRL0Fo61bXf/MNC8zl7L3ZWDWc0Z6kN+K6bE0gWD
xxRmEmYeq6HOzAA2SJx8ZSi/TDXHl3oarAtyNif9VdsssM+G1atKUPwKcnP/7/W/
fgorNknpj3d2xpeMZkQDqK+mM/TRgR1/Kpa+6EcqLI71YLunoaJjqs40RxES11F1
dGesAduNr/zwh/uLEybSBWhqV7ug0cFeNgxdZJsAYBeEqljNZGEQ1pdJ0C1Fd2to
paGiGAXzfCI9pYYkTGKGUAR3VDpYjLpSs0H5VzZRzXQ9n2/Q2Nb17Ik93TfWw2d1
6Qa1a99XgfE8/rtxg89QAsR7fXZ8lAZA80/9/zVDcBTVYs0rbA9roDFn3coiOyBg
aVF6MLqafYCOXMz3LqUxsnlkVu0NBTYiljfJtEoI0vlxbis5vfA0bsU/eJTY0HeZ
xEmkFwMJkiXdFueD6qXclvfXLg/BMEYG84vp01wt1ncu4SwJKMH+eRp+/WiU5h4X
Yxk9rRU4cx5ylIp5PoIn8hu+J4eMIFEyG54/1thmI95cNAxqECm/xvePe49tXkFD
ST/729bOxaiaRUANHFOOSot034Tlhrk8+ngwSSdvc1EsDuK/N1LE5FglxamJaOFv
H0IQfxyWcMVA0jywqUiW12UhEvJ+3UmDSsReLFUWmiTPJLi4tG9IMb5hWaugWNyb
CEaq2mpW2xr+bx0nbsrLtGeXuba3ta8yVILr/+z9qWTpjyW/lfZ6VX9/3hbb5wsK
nkJ9lAscZiBtVhskFArpVBMsZirKGfrLYVIIEToa43zoRD+0DWcSIMNjQ6MENN03
A4gcwUwZRoOn7rEQez2pD9ohqJ6Isfltdg+ceUF5ivSa0CIpIYs11buafpRSHctK
B4Yy8vesctG0Fu7+P/dDFwJvxh4iC4Sl+2+cdGRWZkhbhx/SreJmSNYy8iFpeu97
jQntfx3KmOIllikapmw37IcIHo2jQkrGWCefp4ETrgSrLyNLvbt61IxtATVSXj1t
5oW3sjjJKnX3PQlWciK37Y4q2ZdMuKlMx6GuUbupq0gIJscDmKpUIdfe+zDMrF3e
r4bia1U646QUgp9YaGYMwDUJdqAVidRwT0qaj7wVyzTL7qa+RjaPemW17RVlkqDh
78uySOwACvDtoMAqZjYNI9dh5aiLwENK3qjaKkZ4vUG7YTI9PO5PpCP5D7i72HJD
dwI48pUnIs3X9+ODAhadhnNujcvOSQO8US4vdX7ekKNzUwDzKBCfIFyENEMh7jhX
DzvLXIhWkJc3y8YMoZV5nn4CgDit0RmlsJ1hFLoNRDbQzscX8D+xbXGXr25J+DXv
V+RZ1o8s+0lWVoer5eYlxtDX74Zys6qE4amePFVdOUy6epL+zMdkcTfc7SpAzHD/
5UI/gqwQ3My7AW8bizyuLdq/BtTf5s0Gm/6V2WaciXSODWMfDmrW6Tr6w0NRcb0+
Wiz0d+rsznnwB1oUxdjsa5fEiZEztVpM8nSBrlJ4N+G3ueyEkibZgJslSnA+VcqA
q81XMO2quFJr5VzlYNmsQEOlLKMFZr8GKBAEk+9cn6U+YAf9bq/WzM6DScc4lU+h
oZQRftaITybfvNKLh2xXNkXFN0YvPKg/OT5kj1LiiVFGpRL1koRD8Od6afsIgN/G
oOqsp3DOqu86WwCe8+bZUKl7x7GsQ/wLltX56OovcC7fszC/hYLAR6R1FJB0/r/g
Cl6VUbvWl76IxdPmXTvoAW7sYALWMqg4rMPGSkd7FHkYgv27a1YBFpY31Ey4K9UF
FYv0m5bqM1WqGJxoPFcehToLJxXEMLvfCsdqv3vvInizI2uc7otLuwzzPSgV90bM
4RU5U7QrckqNeu1QmcjAR6VdsX4kEAk6lstKZP9K2pndkF0+//DElfcx4OtMFUDE
NCWyUUnxGfKU/J7mdNJ6jDrtzD+qZtMoDs9nDR0+Cp6lrA/+voSNESOO5qm4fQAD
vgXkm4jni6wHf3MefR9k2RgOX+MRz7brxD+9ynbw5PLPlFq/1UKBZbvMp6UDk9BE
9ti5BAxv3rImbfRZu+JnsfuibuRnVlnROsqSDzo/zEIlr810rBZgn6YIbOhDmpvv
hG4fm+9sYJ6ff8Zc+9UuGgjCk0PUTHZS8Nmrr0Xq4dRi1qQoGkA+qAcf39LT9TYN
ZQWPzpSDJv20xlDbmPfNBhnR3vxe1HKIKQiWrsd+DU4w/coyt6lq08oVukK+nYnQ
oDn3WOi0/sJQm+97PFeOrHqctBL7RYD319Qgk7F1QBZqlAOSKGgI973fsGK2wcAY
vNrk8AYKamLQZImZ5ZDSoy5rWmwpZaV7fzfAh8okokoTglxW6HJmuS1fpQoGq93T
tDg3iAdicpXwsnpT0zTCiE8tOS1Mrrx2+ccGE1YvQHRm2HO9xBc83Nfqp9Q6PKq3
xHgoanBBuX2V2XFvraPtZSBRDPRpwKBlEXXznXZIcFSiONOKoiTpnS5eYtLpyj/P
/D8HO9etAakbZm98Cc4AuWRWHV/YBAhio7wFvVRTi4l/Ahe3N/oWFVc5tLupZYP0
76n+E+6fN2JKvUvHwxjb6oKlz3kl45r5vLs/3Crbb5V+b933E0S4U4gFaSXRRC4c
Fo3zOzQyN7cnBVS+Aw8ri8QHUZHB59I6n/i4pxYSAnQK7ECYd/S+/11RMB3UKKP6
oSlfmvOcAgI6vb2M8u6rFCttk8h8oAZppVTq3vU641twf17O8hwV5/rIfVZ5VmWO
QlNunvQ/UHhT/BtFIt1acwK5InhupLfCtipCii0cd0AryTmacXSHX6VO2OLZVWlT
93X9YcQKNEzyNGnkZObW1tU8HgXVfhOnLv4oKM6rwh9EwktNMvUxetikhQKJpJex
yoI1bq0eC8ncbCJs1GzflY2ThRQzrH0D5XJ0BatLXNQN8Kb1XARuzVULo2VO7yFw
/W+chcpXvwEYSroaRmkOaGnLeSt9R3l9N1zszUUykzXwk2cd3a5/dSgBB66/AaC/
Z97Q0nFpSjvkSRfybCbhfUVoc83t+OTXm+XR0lrClpryqRV8z/rUPPpYKXRaFsS5
N0OI1EInWdZGXDSnOlUEFmhnYQRy7rCIC/L0SpgyozuF3kYBPdOO2VKpHDi/2svo
op1/d/BCs97WDKLk4IxR/eNI4tr+I/xtHhxb4J+s3d/i4phNfYIHEKRbnPzZ5Jp5
DYbJL8IT86AGX5Ygt2Hc0LXq96cdz1yv1PYtMHvD2BS1r7o2r4k7j2mIa7j3rdDz
a9Hm8biM1UufEyS8hmpHqAFwG2Vn0TSac/p1ZuebesV/845cCwQc4bVrPQRpyQIo
6CwW4XaTfN/A5gqFB+GTqODy5ymGk4/G5/7CpCA73i8Zblqz7V8J+Y8+vldynvGm
C7ISlQ0I/4Q9PVPeoWFkYt6gNJrrqXgIj/X+kbL++DKE9Zgz6Xps0PRfqyXG149D
ZRxxFr3vCk9j40AULS5N3/3nIvOna/09+h0/u1PYHtVtSe73mwrzNEUpAVFAKdxW
xnxJjaVXzkKpARNaluECdZJlZQHnCHCXv+rT0vGTg/45LdnNRX6AaoxVRdFp0NfE
lRth3AgSUVtdMmpAqJuJBqemLi4p2uxyFoEpdADqRbmLmscCguyphnvgcedZRvSR
Xy9a/Fv99tuqS6B3P+NSQy7p+7KYmC7et2x2fojv9JiL491XrJtxqpLYi5SNmb5Q
gd2st7/BlNtzPJ39gubLo32V5cfZQFQQlTwbkDHpiuqfQJ3Lm7j0Tj470RpAe/au
+RB23ITvQouuDwcdcqNGZxR31n2hirHr9w3S0Wfxt/AKmlxGzbAugVPWl4ZN0Qx6
NrGNNzpTmj3me8jcdz6az6/WJEd+OHBC3vTKwddcUdWMU700dGUyWuCVp2gpG87o
CRNq3GJuRI1WSinYEZNGSuWqQo7+Unttzx69L3BrCb1PEiV9/PUfzRhC3MJ+FuO2
xBFgARjeQnNqQFxNYcwYV5yqzMwVtMZg9IYcYmnoKwsNi5LlOA2bCPmbtaiXyM3Z
+7C024N7mlbngXno76RQJFhm1zguZDUsbDq/M001K5LGPOLG1zONTC7JIOKL5WL5
C96uspsBb55gl9wyW4ZWj/CdlCqfUR/gO+5pvA7QVG6+zxA1RJyLp7KO+6WLUYtt
0HLNxz+kum8PDz5qvV0c5s2ePc1hzRzXDZMkRq0AM6tfyVzt/FxqtEJ/KYuamr8p
2arQUctCwMTgO8p9NTub6ueIRL2BqxC1IMvGeG4OJSyGx/+FnF9MiZjVKKB0K3sy
+NgOEIM8QG0uj4BpDnWly5kbD4ZKABEpqnbOcdkJtlMMzhn+LiGKmlljrE8DDu/q
cBCboC3C2Kyb68EBKiFtedQXJl0aBTg0kObTWSuaPYQVGc7G+7Edl+RK/zYSwQVC
RhlZfnoDIbOPAFFtErT0fcmySp67Vfx+gRMAWX3S3gHUIvemRbb9gRkupoE+Vb80
wvC2uhYvk0LBCDC+2uWT1ORKdcP0v8HV6JZABH7/6tDHSjbYe/nQNnA6EQtowJ56
HLn89i9906EzwrAtFQJC0GRB4ID5/xA0L4vuydpbWZC3LNXq8N+ZKNHoG4dJHgQg
5hxoqE3UjO3XNBmRFTxD07jk6DGPLTOVpQuhl6/Hd1jQ6Zz53o+SWJyrTeuooPvm
dXzU9TsnpXlLhBf3tvCUUDJgKiN5/ea0UICCFZIs+04mb9v2zotoN5qo/9XCvpNg
rABoYkKQZdX6iCruMpRa1yM5XiSzeWIouwaPHqrUazTmwJDRrr6WmH9uUI8RuBkW
vMXDRc7ON6YhKmgq82ya3y8BVR2xYG93g7RpumBSG/uFEIXDowP2MlNXBMTZ9Z1H
xNkpwiudxV8hMDT9HMmKvL47uvrodiowXWd7Acrj8HcfbTP/xXdD1D8aPVSGybtn
Y3gJiKj7tOq/Nll/RfVTg1DRDXqDyODtaH4puPfwDz+LLcdEcxG14tB//B8sRR4T
LfK0mcN6EcuVZohwSF5rjkXyFmMhGNB+Spcm2L9FntAMaP0/Ur6qv7siZ8e0IFdZ
FBnA0GhqjN+czavx+u8KOQ1ZmFRigtDiNkbDBEIIzPrRmNDCHYhYoSxIKEIm/06Q
ywGywvjdWt1IsQfY4atUQfPTuGWFCJBt1wbpBFO94zL073TxTcKV1mkIcPX6UGGx
GtcxRe7L39dkfiFjju/9HrlMtREx4WtRrkFaqGGJetLgG1jz6rOfHKt0Rfnz3XJ1
iJiU7RqoUSZBwR0ZCCizoRSc9pTKOV+c6I/dKHETYCu8A5g6lFrTuUVFhSK25FsB
11Z9CpSMx0TQLSZpHBRRYohNQdj6mwa8u9VgrdSGwecbHqJh/LJWms093H8bAPfs
EDvo/9pwdCFzc8QK1VovU//XEWoBccdl8LZFfMJ38P0F4sb1cxs2Neq3XYVZO07b
FkjCH6mK41JChfnTyzZYulwgHa0JFq2iuKeNevCuvzOMwgGsbpYd6bxQKrlIDs7G
SwsHo56SXZ/pwVhixxyNfgqvgiwcisCCgjORILadyJCDkeMuOXYHrl9FjCfXyt5J
azSfUajHRQezUIbLIRXXftpZxKDjqabki97JaoISsMP47Q7Lhj2PZWl8psr2wk4P
Yu0FAYOe9lRLqFHE69fWnOK2hJMqiVAJpFfBTz74ohSKXd8ryRHHcuLBGPntGDdM
tJK8ufDHta41pygXdaeHamjjbbmtRfRuPPK/61MU62ZUT0WIx+mxCeh/2fXkHRnj
x8lInxjiim+0Mc3xEVxmhxu5UR6GYDrPw6E9vGPGfGxUJ+Oq0WUlY4MOAvmDhb0i
t+ZHbhFu3qeUzWOUpHcJcb/dO6cjzn1UN6XQ4dNeM1jHzvES3m2Bemt1YHqUEIhL
fC3uxgyT9HIAYrQEsR2mHkOYY+xgTT/58Eedu3RFQey2BjyME+7SnYJ5TrPfuPb4
wnvgzMYQ4e3lE0VCtn14hWwEZ/vlFFv/NvA+syh3sXXFWnd3diYqGPGaqbTnZol2
Xn5CoIInvrbEmg6dgT5l2VsBYa7+IPDXiFRVKenP/WQr+krbqjvd7+WT2EyTEnfl
y7j7WyWhbKVkhtjkA7Tw2DAOYFMxcLgLCFiXg/fqKp0MlRTCXhzUXyEvna6fYna6
Y9rtpI46wH/K0L0y7OHuHtFUVfLjlKEYRMzsG57kUWcv45vo/Cav5NpoVsM6oCUF
7XKdigafPhr3MCPQ/GHTYiZmcgtgU7CRqvyBvpZ0KeNDHrikexc4upVDKgoDO522
QwLLqSeFoOQmPJy1DJ/zKdpjBfpHtOHtgIERezrp8plQbZcb/WzNzxCKAH4aGhLY
C8pC9S+WO7wCDVym12630/meBEtjsnq1m1pSMAoNNfGZ1/6uMgQnnnlZ47KRZbIU
Nl/QjDyBAhlC6Gnn9Q6PCFZRiD+LRwyAYM4TiaIJpFHOlaqErBWSxrTHXHvVa3UG
CCpHRirqPcvq6K3Qcx2+GXj0HTFVvMm4PcankGSX9IZsBhPM8E/thPXmUnmVn02S
6JJ4scLjRFOwEXy3iFMpgJ4wd3qIuFqC7WApAZKVIcFZGyHssAguMmDGV2B/l26a
wW20iZdCufvlLyh3sfFy+9lkwjn+cvMl9y8A+6ujm/5mwS40MNtzzqfAgSTxoKws
FMewz1daPptVHqeuBRBOWbxy9U0CiVV3U+3l5+E8OrcIb/L/kXqh2LbWa+PD3mYL
fhB42DSsBxFJoq/t3KSrGPKrZyM/wPh3NsfcAgtIRrsudQSkwovU6Ig2m7Km7NXA
LQuFVxdulT7M24WHTtou36w2n6KqgZW4Yatsto/PHsFj8wFaU+8Mc2sVKVN/2nQN
nQqLZthwgeCNTA79dK1pEac49A2ygLLm8mGuOpC8PD6KdfBQw4AwPwL5bFyq43Rg
JzUlts6HbE8qTUFee3dtna16oATwLmRsRzG9afuaZ1r2CWO48PvGzKZmXHddga+M
qvRIfCHiGK4hKPX5J+fU+uGzzyJK2099Pi7RLUEzVyeR3epOt8lqMP/X65nHcYbn
akwF7zrTps97uD3978xIg+u1WK8wQ7VZbP4mAeFUtM5qQrX06wmZECZlnpnfkZt8
XCUXer2b1AL62MX2bV/8NSTulh5HAOjtzt+gKKg0D/G3l70zNMOAIo/NEUmkiOcb
InHaJB3keyWwIe0vk8KvLGIFWrwlML1oW9lQXIN3vmwTU0jnQup5b0+4TtjguZFI
PI5rlbYvBRvYHUGF5uaZHyzI3PK1tRF4Tt56Qqmzq3jXEoqg4RgiBozWe0c8Q8Fh
qxQ99oAVl11fZJZ5HJGhBhrUwNzuxsJAzfM8j7A8gzm783DiR2xXVn1U/029r2bh
zQpfFWqeGR1y8EZ+rWXUfE846QKw+uM54GK3NzP+cmgIpp93zgLg3Tn1XeKRAwd+
4L3EUgPriBCY5N1C0TFCKVUAbrRH2bwLImxvwnsUfXLqzYCvfGZPC/gEOTtahv7o
ZD3vieILbsxeyE/RCGz8qgTLl9YvFgQwD4eKsLagYVPYk4Rxuvp/rrn2MovehVEL
giL1/JO9JjPDog1N1QCaxrNkhXdHvDR0HWb9n+yY6NDQ8T22eRepGNz9FyUK2uvw
whW9Z/fik4YHVNvkBFyu3kNaS5zs1KGobsCeP4RXx73sTYGs68suIuIwaXkVZP0Z
/SCeIp1iJwp1lulSUrZs0RNU9oQMaRb3K3tT/5sVeKFZ1F3ssp9EBrXirIDN8KEn
axgUiqo55u86qltXZTb8j8cmGXaslpIDjI7fiZfoHsdFlXOKkoDW6/jTDeNwtHek
ZGeooLCfHoeH7OP5gkwS/HZG9QaoEsHQ4N42m2YYs5PgpmsPVsYZaDyxVV/F2FU9
ehINpHg4G0wfNGIyWz1Od98TGkqf2f/cFwf7miwl/25p2/DQMsv55ghZ/vVS4g3z
pGSSZu6fTvkQr8HilAJO8ZGOORm9ujc//aYLsGH0FOSQYmAlOdNoZxhop8DwgBOv
KfC1e8goHfJSmNuA/yYKv0t+8IkMN/Ctjczb6XMp6XWnroX5TxyLPs+cnUMmINCd
hos9Odf9CHxJh8Jz0ijvUAEofhEp7CkO8cbdKSRgCGup8xtzuhMHCjxHciEQ7+PU
AMuzlZoWHs7wZeZlVriSPWCiFes1vFz6aqG+CujaUPUywyxnmYEB30LSotpiMYCN
C0dlSd0rljZpdh2BRbl0bypjS76l5rO/KfRINemKclCX2o4qNiFhe0+X5rxvis1g
cTv6YP1uWu7lSQZEreVSaDzED/nRT133vz/VU6XUuthtpO5gteGNqYhenG3sDMdP
i1muOkbOJxzOJwIRvtQzGsMu+//SS0/KnjYKBSwdtbKIzvE6d0GJJSxui5c/+b0o
7tQJ7WzWdiprCyKFEZW6OuJJFSLHOcju8zE4Y/hyPFJsuzJ1xg5Ahvk5D6+NCdNm
DUddhWT+938dG/bUTCIGfDxhYstMayGzmarjvqZMnNiOb6jZOifu8VspIzexRC6v
jr+7vPOaeWb1hMUvZKKrAe7jjoYrDYv9m4I/UnLE2WPVuclyO71C0HhcGCNyWMXb
NUOiPAdVTKZWUqcK7DXpsbLQ/kgnKictxRBqJz5T+KlDr1WQiUNng9Yi6NZcaGBM
iv3znX1Nbz0cu5MuWqghCfgrOTv32FgqAMnzqRP6MZgTFEXRsrYQ2VTL6bIezaz0
fPvf2EEU5Jk6DesD11XsKCQLASipSt/WCvzmMjbpzvGOpDEP7KzB6tQxxm6lrHLE
opvf3vrk8zL4kl8G84UxJ9zC4WidWAXhR0r9Nt4EC3ZGlF/80PFfNSKNW0sK9J0+
ScXFIjQ+CLNfrbsW39xGM669aAGOTFKVdQIg8hO+3Xo952fcZ96aDmm11bAmT/bi
LTZpn+POcszrNe5qNVIDCCGM7Hxx1j+ZfiEQeOATPUDm13a+JBG499NIyXZFNDM4
+HPk1MFzUtri8C67Q1p7HoSecNE/aeZV2hFiH9Q1xPqqChHHZdBTUpw/dn0vbmYJ
4/0zhLqtgb2XLGKlsbnzGLjAFQFNR6p7VHLhoNnA5NO6q7XKM8lOENBHUfe6Kzpq
W1SDIVeCCEosY78FskjmNfYMZ2UrVjPW3tz/K6N6+o/Qn+RJmfFzZ8DPd+CiZ4wO
gisfchV3gwtKGg2K7leovSTswkcR28L6uQynoGLtr2KdJaaRUx1srahyvigcWX0c
P2TQrD9Ps/6luihdlAbe+Cs/KNx+gmsoR5f8LG7VkCybSyO1XxM1NeFXZc9F7OpH
AYJUksrAla12kIdhr75FrPcFBQDevqte943LEgDmSbk7ztLIWfOTD8Gd2AGTvGUv
Va/xXBELrYXZX6UqRoVMm53PNoKq52dxdbjzLMkhqNFBkHd8PWF6YGeMcn15IfKI
NaemsOvu9Tu/p6esvCn6PovajhH6QRR4vZpVc+tHpjJTe4vZ546/bY5egYgxbC0T
R947eJ1LxXI/TpczGeWnx2A1krSkaa0ANu5g35KKsD1zTE4ZYTaQ632Y7hNLZqoN
8gMdAHm3znDSX1NHjnKHnMgjL48AiBwyCYrvQVyhqzB8aqD34kzjxxEwN4DrRJmY
eTqxCw/KJDWY85aioli02wENSEG4Gze2amgYsguSOhR2yQk04NOggH6VoelOCjVQ
E/Em+Yx2p1jEpyThSckwXLH2nMMLNsE5gE5TujhZr1rrCxWAt6NvidZq1KONecjW
b5BH4Wysx8CV4hoLm7UJyQOA3z4UNuRFINolweb+VmT4tWUkZxx3A+59wbVVeXH6
T/BXuyYSJ3nrsOrF788eJPLYrSTd5+p7fYq2uBccjoSZkgkKrSR6Y1w0hMc2Hezm
TGzBuAIgmkVYY55x9SS7Dvl7ec41fZWH8xzKVf6nY4DQ7hOGhv2LqsfFkE1ELn8H
x+52ZzXyqwNqlLrCQMJ0k5JgXwKe814YaoFLcUKs6q/khMHzriLq7WyCyqMYOMHj
juxnvGr9+fmo3izbl+beV7tCkBMWiZvjAQlHdAyO/uzpf+G0gYf/VdDa0oZ1EN8j
GAi8Q8tPuJZU3OHWbSL95aEbWXYD4TJZ9/16FO/srNN5LrUm2BcMKwVK/DCzxZVy
+MNDPAJ+o+PaBhJy/Lm+mGpq0v+OZeHz0c9JjpqlzrGMXtch6tSp2iRHavrcymfI
ACrokat6MN6D7RPr1mT3Uo0CoTd4WOrJFrbm5gbPtxECJotT1Mba4Ad6oXVemuEi
XtTa5U4IHxtve3nvOnVwk8TXzOj+JSzKCCNLInNqWxw/Mc9gKdQzDAZh19MBY3hG
y1yTNiQXXXru6NbV8UuOzXn6SeJq59zimFPzSk/CjErNJRJm8aiE1yT+Scjw6T9a
4YtaDCVSnoN9XHAzbK0Pd102S+j3ZHoc3abP3jgYqDZIRVjRN49ObI2oo578HZk5
sLh+MW5oBZaXW3At1ggK5IuhpRxqxv24lvcPvVvRSR6BCUqf7dLFN56zHqWIXR+4
O+TXrmzJjYOKQDN9gp5fBL+aw4qOUQ4VHVDjAY+7QMRwzA/xGUoqBgoYHzU+3+9v
ClF0qTy8I1v4TxCHKGwn41RzSMqYgYIjXgbeBF3LG2Bj9ztmkcXJ8qqIdAJpK1Ba
1Rm7nPjRxXEalwmFHQxxROU3kH/qyPnhcBbxZentSqyhhE61hNGrNZYa49qFeBxq
wdK2+B2b2bs9bFXg4ZS7tnvFlmqWJlvJHkDgU2N+RXxXtRyD4pAqTsHdol5ieaNU
aUEA8PUBlCujgLBObDSLbi37/gcMgKUVtxsaT8ZSbFM+EIAY84u64SiD0GMk5n29
1TVlVSRDKdDWVdnK2sJY8suwzLQcadxRSSDDhm95Co5NmEOd35S5baZVmnxiz7/c
QZT+w/Ar25dp0miCqb66FADhZusdNYCEBIkGjmvPaTkZsJsMskjCU5C/ub/SlxBq
3MliGXwXSKYdlPbZVaZiVk0SE4H7O7KHbsdGjJwZJGi3d9ZxgVaVRwyxuwVE/pSx
Jqb5DsTiCciBScrXloI5+OwcQh8RfSCVVoFmEW0vUcUSSRDH4F6+Ww2IHasHnisB
YcaTD76frvASr8EJOkPqex5eo4gRdCqR7aihNXUMO7uEnp7ZmrbdAbsztdMa9kAx
mOrqbU5OqpZTuA+5HHyjPAX3JNtF0Kth3nXSRhjzFSUZ6n7ZckEBrdh4yrzIf9BA
H/VBmJZGta/HdqCkuBeZKPIjUmzYq/YUDrA9/8ElaDDC9eD4HuG5rM2cZqX2tfJZ
50Sm6oueLyUjXO55L4nlfKCOT/TmHXr0uqdOE3CCLwKXvHJAF3Ys3hODip2KFV5J
a3e7yRto0cuJM6TtlIqSG3usihWLsWGha/GMA7OQEDSNa8+lxDZfqm+IIJS/29DM
dtV5O+4vYJieyA7uyUZ4ZTOKKG0vBzbRQMLm0FYRhhh23y6wBKTgI+QlBPF6y6UQ
CAGskPaOpzVxlzjzHOKrTnvHxzhP1JbC0eN9Ahe0lKW9hEE4AJ7PMlReUFnwkmfN
LV87r58d2o/80jYeSF0EqQf6U9yKx3QWd93sQeFfYf6dGiP27AIIk87uKFRWYQuV
M1Vi456GfsuBfW+dQqatEhwg2wKCiRAPJougmiuBusjijDcBS+AzMD8gFrYBS0FD
5JL6YZeNdx9dE9/DKnVrQtlFfEqDIKCVoM5b9ms4ma5d/sXY7oYLO6pX4lStr7xH
bRhYK2V8XO5k+fLz71/poCzS/aIMj/1iaBu5TPjB/zofW3GQhKtpxGAljNozsrD+
G6cOAsyXojalPPkrWr/8XXWadIQxt3sRSgihbCFtl80G31g4PRvVKpVmrZaCZDZ6
sojSphV43QP5Y/ZZp4NkZsRHJ+b6pXiyTatitvNcrp9RJLAgUndgrXOquq3K8m+R
hZrA4+Um5CQ8zRjDyjucZ/2Dd3DceXFc9MIxCq8yZAqmKLsvlDV/ORxVo1mzFthP
goWsJUqlzosVsePkawOrIFrDeMmDBBRQB/ht5wkDNjtiLHLDBGAirRE5Atby0/nB
V7NATMD0KyHqBroocE7WqU2Wwn7o9mhtqED7LGtNnItpacwASW4h2Nudb+Q6XSVv
0REEs5/J8vM6RBuJ008JjuTaUtBODi8VCvpXBPC/gmm9R/5AzLALKwDsf/1HLqtO
vpOzkjv8a1dAbAVc0PDPA0yjfRRtYmXCB4dkHscxxG7tWw+ciybj43jsOn2vAq7o
7lQ3tXuyeP4zSXjnoxN2CTikPKvEQ6ce5nIC+DZfzmEg0A2YyiS7ZPu2fYz9mLBR
rqCbGZuNPB8VqT1kl8BO06GV9mOjYDdk+1VSnvM9pNjrZtjtgLtl5nrr0pofNWyo
/8RAlbHV6TdRxwoqtXJ8dgbKCHBXYkyItdriDRf9j2gxEkNsirSfdgyJ1LHxVuTT
6W2rZKFW+EHh3gbPOsU7PRUJlATZpXS+unHdqWk1jh+eMDOeGntf9XQZ3jx0D1XI
RapIfil15KJaYyskUkl4FT4KVIkwqteYA0SgTNexi3hTdS20X6tF6Un1S3CKvGv0
f2V8va3ESHe5DtgaPr16KtvQY8eAzvT3lg9aZHNI5G88ypHauHDLaNaKQbg0X15+
WbT2lOy6VLisZeV7Nv8Nwdb6TpF50Q6D4j1hkTY8/PJ8q0I1K+M7114kxcZXsi+L
1rlun/PqSjI1pAGen1XYwbiW/H1NIzCPmvLbInxCTCtXrDI3YREzJnMnUpYxIdkj
uq+VNrNEROduk1pE5qkFgJLoGrDiQ3ut9+zfoKongpsCdH/QvQTVz/dITV4mmt2X
KQaOu1TlDDfTOLbr769bRLxduJ6/Q3j+EwyxszT290woPPXcHNiv9rkM3gSCH6Ga
EnSZATNpHPbIXn1ShpLxRNAwxPp1cygzA/VzktK3Howlu8krU4X7D6MpqqPKnY3s
5zu8QXh+2rSsnQqz8IU4SX3LbTiQ8uOQw27OHoNq39ZSQ7yTjlb3VAzEdrLcrt6j
vdZCmZhHnd5NepgAr9xY0pX82N7Jgy2moN5Z1LvXhBzNkjj+NwYOr2HjERF2eXhK
gHPjYTsasV8VKghsRfx8hB2L9zkwz3eYhbZXOuejRubFEn1nkawcm0qBunD7uzU4
Og+KQRQRgWolsohAm8ga6xRzqOwKET5R1lbUusxfNilyzibPNWWh4OKzujcygEvW
IPXMGuQYhlDNEg0lKXUIhTDDZoYA+IybCwZT5Y0Y0EiUv30QIctdQHjE1GsD43Qi
jtd3L6WxhktrSgmXqqrrC3bl87jGifaY8dDHT9iqZxJEq4rAWDIA3bJFt4Vp0Z+w
v8l74ZvJ0jyKinafE3ao8g67jGFMYYDj2Q71JoXhpli2v8O51GdmYlYoTp1Vemjv
pBp2w1Y/UlCSk3ny1yS1wttKWxui0+5QGj//NalgExxH3zMLEcuDqxpi8lDtuFBl
ZoVLa1jK1ufELxojxe5NGhVsUZMtIjj7+tJmQDFSKhhKRNDIeHK4BbEHYxi6O26s
OAPXksC89LCy9UY5O/3XUYC7onk9/toIm9YQh/fd1mSHMflzmWDEqthsrjKhDQ8a
QkMM8EBMXVSxDGLB1ZVH+PU6mXcfScya0VqMbWKX9maKL51QsL/3pEQLWUflM/at
uoPetvGUTwgY8m6+8uwdXjmN1/vnd2QfMCTVDp5IHSbq5YCM8d5LhNA9kTjQ2dc3
YNyGaEL/Y6Vwvdr7IXQwWc7q5eProZD5o9X/EEEPm7bWhWUEotdVgVxXrQtygxIb
ybXvu0YeyX5Xx060R0jCCNkuqOfTvCx7+p0RSZfbUgwh5iqnmB4C9Z3No2bLT10t
Uq+VZrZLDsNL22MsMJoHeA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zhc44gNZEZzjuDVVFQZYCfXoaGhBXDgARsboJExX04xTgB336APFEjNWgtXDb2A
5Jw1ohpLO9f/Vn4iCumBZ05iwgGjN11pfS1fawIYQsajNosfuH/RrDkwMqu1l4zz
FVJxnSE+SqguscgHS+AF13w53hIuivzjfWwmEyy+B684bWT/mNipIqYAJoble3yY
Gdmpw7H+kFegyAtqD4ndc1/LdaIF9uuDhjjaE7R/FfSj9wZ/8864pjNUGfri88T2
wXPGJv7Qg9TszE/kgna/pLyypUDvEHl4aXyVg8DObdp4ZglbHtwc+q6BBIVCAIwF
9TmnDbkH30g4cUHZRiTFv6M8qKMLMmyPYTDGafNFaato9tADGQs+DDhnGxaJu0Vq
kAB2EieH98X3e2ARMPZvr5apeJPnDHRKXTF0PGJfgrXnpLyZqpqJ/y25EiH2Q4gT
NamlX5pAL/vehCuWSfFstTR/uadA6Hgo+SnrBvIfCwb7Z5mYp+SNdwlQ54bj8+mF
FLmgKciIqPLwcrwwMsr4+H6O978MgArWmc7bX4+ZiU45t6XgQlceNic2VJzieJ8r
+YSPpgziIpU9K3NL7CMraG9I6bxX/3aV1EqHON2adEUig5aqnWEbgkYR2Hd5q4It
EnrOzc14SasEz/n3sHQrpLDSQYN2iXK2FQxVYnEVhXu2vc1ahS6WgaRWQGQKaZZQ
ha4pKFZQ8tOh/1xqjF1hcdafd5U3mUL3os5vA4q+LiIu56Eff/4UeakM/oC3aWdE
3Oj13RYfG6P1NT3YPQDtNYn9zAHcmJwRT/k7es9gy2AcfMwpr4QxOPfDYGksUg3F
kqcPCh8eMYo6+8eXnqNaSEuWX+qCYsryDwDGr2imbcSN6w5v2NWkTeIS8zhI/+O3
hU0Q0LkZfk9jE2n1U3vLvRH/u498qhO9MzO2bueqscI5VouN2n4fAG05WGams6pP
yoHEvPf2UKeXfi+fEuauFGOWoJSNyU8+IwHg2GiaSOP4ryVYTOeXsE407HQV67yp
JMfLt4ZVbkKV0XG+rpCxX7n2YoYjlqbhfmm/t9I0hvaEdYnU8SNVyJQo2UjDOnB1
Sy3ekP8onySUnWfJaDL+KntG3m45VQXpZEf6/yfVg4o=
`protect END_PROTECTED

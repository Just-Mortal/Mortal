`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LLOFV+c4PAqmiCMtkYl+7BPDFvrzoiQLeo+X1FlefcP3x3VLJZk2tcnzkSdcueZz
OMGTuq9emdag5Mj4ChJKB1MBonZSHFrvLCwL5rdxzZSAxCwNuOXqU2cOvkCjLrqw
oSKlQ8nO1rOac3rlEfg/1A8TjjAcww5+N20HEKKSAUJPHiImZtzbVFzwX28I2wWa
Mrf448Esgfv/oiYj1fS2ojddFRk3Ou1yLGL5+uI8DwCfcHZR8zGqZfz/w8Z1CIDM
3a4d/jy/2s8T6JFQL7NOgI6vxjMtG9MR6zBPl8ZgJrz9qlUu4BQ4x//VWVjV4w2y
npqvyYsEEw1qeTH4Rvj++/5BnIAsqs0G73pJqEng872FGx3M5zpCfzcenBZYYw5K
Gg64rSvSYy7nQdJfKxeMEk56rGnLbeHUg6yLTNeqLCZyTT3z7EYl4fsBKZlRMkxU
RnPIVrVc88noEJT5wrI3cDh/138RdzgjrheQNxSXIbkNo8g0Dcwm4SgOYu+nPqQ0
ai10Uuscr4XQbsDue+wV5F8WarOuYp0XnkHk8YhM2Bqvw/455mLDLU6r9QVQ5ENC
0T+qBpo9kTNnd7KNrqdZacDEDYPBCIxWvr6DkF7IxpFfZSgLqbxWZMzF/YqMKopY
eGXHAQ/4nPmouUNS3DiKzEO+3UrHNgzI8ekhC5kHJX6+8IDi2Vy9eBMIJblw9bnB
s2iXv5gxENGEgKnfx53PLNqAXPukvE882laD/5g4W9Vkh4m3FtfNyFzHABhBNyZY
OpLeeG1TUSasFGyDmxUQMDHiVPHaD+071Cd6e+1OvfnM/fRdZ4Xukl+N7FQYs74h
VN9W/r/BDWLoL7rE728SJi0Deif7VRm3Dc7ZUfMeSVHFsKDyoc7fxaUQ1MWLRToP
67Fyjz8UBp5HE/mq8u84FY+1jS+XA+ZptWFt6mRqqSQ9TJn8G4tUuy/9kDKyOcJg
8aHkZmH2nM8653pE6lWghFQOfyzT9s8Da0ipHx6XRgU2rNUTfnuzrcJTg9w4pwGb
WLZ4tAt/Is51IiSQJNqDqmFZ+sWhW8lzI+objJKDswEJ+zwrBwLB4bZNbWAjH5v8
mlD0mDR4/ae5jizqW8amt8sGv13egghK5gKHSjcm3erEb6bjMpzMo2et2CiToxk6
FQw6MMD4Ud+18esa9PUrWhReqvHQod8jwVNMRL6IsyYfK8quCgmS+TO6X+k9Cwoq
Cc5hs3SZKRHg6YJXJx5F8eqWdpkbW7CH9k36HNP7ZL550ABNZgtXsSHpI+AEuro1
Xn8m2FBqqEk0kxJ/4MnOb1b/F0y/xA1zsZQhm0mC3Rwi66x49bhfAo09ubEBYIYX
YzjEAtQnGB8Q0CYc9FGllhzgZMkTFDtk0ORpMrnuPTI+h7e3vezY/qXGN1Hhnmrq
6GUNdv1eCTarLM9MHLE01kg7rngjx16N5ipb1vKlSpI=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DsBdSSHZ7HnpdCH87Jmb2X+30EAx5RBcRJi7vbirINFPNOmQOoRK31X8sF431r9n
q6Sj5+eW2FUsAzB9Ha3K+5LnKeuaq6AVUMdXciPHbSOtJynaBkzVPe7J2C7bdsMe
3aacWX2IhwWhdU+NBGA8mJqdLCas6U+tT0yGcv4bl6GrrxQKyCuhAaL0LIdJ3NzD
m1NU4Ql7Cre8vSOLouRu3oDW5RsMHyz50y8AYRU2b/0CNCoP86z6uZrPUPMHGewE
FXUeYnH2wOPmIIeMKU2+yjosFONOw8zeFX5hM8BS1f5WkD4WKLrQYx6u/M9NahZw
Qd7TKDwNz43D0hG0Up2JfjoWOPacSVnMQabELGq86j7LhVh1M4l3ceuM0/fYSbvZ
6smFkEt89WmAqKzMoHNxXCT8Qwb1OQQ1ioZ04GyTnGdpPVoXVzhcYdiu1NIU305f
beZD3Oo2ssk0Mtb+U+djTA6wsC7yGpQkZ7eS2WGXq483UTwRO5ItizaLvYEUcPYh
bkWm1tiCus1ONr+H02mB2FHpiuHuRcOfGXMg20MFfUqsjQpFhWrUN8doVVqLAnfQ
lUIhJMlucyXe/qXj6EIzSohneP1c5FQuoIePSiwi9SS5KU3qClUcRBveLlezEcpV
CsErPZgQ+0eR3YsDxNnrmnScXA1es2Lgr3MgM2Ujm1YbnAvqSbXnA1OAcMmYzhDG
5V0xOwEsPrsOcLPAnlHgsPE2dfkrH4zJinlF5RExX8oqhpegbVqOmb8oW5dXouWT
kulJvvhH5/L2/u5vMfIRmrRn9uW8dh8VtdosZ5xSe/oPyuCRmWf+RgqgytSgBC5F
c+RnjHzAIlm2mp0w8OiiEX2OYhpyxCux0msTA5b3doS3U1/L/s2DWsSzrJBF+M67
1M1Hf3Ti6wtfapP+1Qkt5mxBV57c6rIZuxhrS5P7RFCbgOECq1KCjFDM3z+gXsup
IZ/eAuJqNzS6ghTrffbzb0O6r3YwGzMn+vn/HQuTmbP+clQ28bV1HLAf4HBg8i0U
PutTf3NoZKU6ft8CjQcWFTyMT+pF85oFotAQVLPLB9AHhlRrh0zHmu06JRKLvmlN
qPzgOTyM43n+hwyEc0xoFpUr3axhPIE9m3iY4rmLl6JJXsiYp/S3XJFYWEn8xpq9
PqhYIKQzcrdpCIUTk7yr7vXS9uCsc6zfN39RsWth0HbzqjTrb33535rKkYVnUMg0
YXtqS7MPW6D4MBTX1hP/4dL70H1j1LtdasqGEPUHTSeF+tkC3w5ydl7H91lzcnH1
hap/70Dyk66QE+sziWGFvZhHS3ot+DTQsR43x9m2yutVoFNlykdEjV+A1+evpBB7
91dge76t8ffYH+ufgyypjdCwCaVoUvlkwfNnn1ZgN1StvsUdfXer1lA3nywDvG3C
HHl5t+L/lvKjWRO+Ta5RzPz8tK37+u2PPTy5qSLJvuCvbnW9N1opHxY/cB5y/TyC
i0o21BU2idsAAsiV7sZ1tnobFNLLC7f7choC0j4QYvPrSMuKoU0oIteX90yRKN03
/sP2tuOr+7IeUW31uDJtWJU2FQtpZPPi1llTrHu71oS/kXXgHwv4oh9nUhpPQDRK
TCDDRBTJ+UuxpV5NsxgJpnxsnY0vAJO/ewuZ0gxzOSaaHo1pHfoiSRW/6OyFA2dP
QOU5hjFsAuzqbfJe25Zh9Cwm9PFFq9fa+40McMDduVumORGJErC8TNj5+y2CUwyW
VNv83/a19aL37UxorHR4xfbZxB2i9Eiuf5u+ZmDamXloH4JIJZ/jVkNRbJTZ9u5z
rWr44lJc53nUq/jGkVTI9CYfE3wIE/synU+pUQSEVxOwTxQcDmAQ7grLhI+8Bcsx
zUbnYbf+We1MMngTc3DdWsrHqb2mKHchOtINUgv80IftSPbQYDpHFQK2xgQIPwpF
FmtiHUIsAfwyY+yFxnFHq8sMv9sm+uR1EYJix5T90nEa+boBpkdCZ+2GI9V4+pp/
i9k5dWQ1VRIVUTdzJP6hL/tzbYl2aT+WG1OitavZnMaCwU8uPGKOjAAc+Dv5myci
Yi8uALJMguz4PKK845tx2UEH2JYctApofPp4X698NleFTY6F2VjnfgtVFzRdVaLu
3Q0frlQB+lv+EowcZQxVeNn2s/pxIo2rKif+lRC8B41b2uhNcSuYFSc/G+SQe6zb
HTFzFEb8WJR64mAv7H9sz/D/zuBKml1CS3yA06g6TLNslmovJqGKq2NVnbg3ZwIX
LrjAeCAX7FzDlasKWC7CfVQbzZQGs4/owikTwxDnL4kjbT80udg9vONu6Z/AgPWf
yIOEJuKUMVB+PXcuAgMVwLMino8L8l62fYceiZ500h+G+p3V483Sl/znCQnf3Jhw
he1SmBqQs3gr7sNUeCpn6TywMnrwOI5V0a8Vs4V/NwUUVB0R+F+xVoUAxiXEE1nN
4xdtuM1uMMuaQBRhptlsDdIBPHEqKGru9cxPkVG/BdR0f204EXU6LmpF/M1X8fSk
6dQv4aKE9Td0f31jnbz04THNpen1Z2vpuYQJVOW2zdGyhvfeVncSThXHfsYtJBZS
K3kurvMjrl3OhWConwppAzwlB9roTFSrIgRIsoNKfQlaERzk/TD3acG65EggX0M+
WrsiU1LMXpqkWE1yB7Y8Ud/9w9xro+9i5CY1Sl8AxZMBdh2ocrUeL1s3kp6kFufj
gOtsonR6WoPQ35klpU0Us/1sVS6KEcf3HfBkCiMzIillQqQ9PMOuSAhG0OKXNU7E
Lk8qYfnvrEC0JStDTi2Pt/uLbyELYdJ7p4VdesK6PJqcnG17nFOXzxMPQ7P3A8/5
hwGQ71wSv0BQOcqwa1fMNYJG2kIE63u9Z6UUIX0k2N0w2AGKENGIg/Dz6ziwMZnW
fdDMQh/GfcbJ/IP5LTV4NlLhiHKwG2A7Ln64iDFm+tnIhr1fSI/YKSlzp6RhRXW7
oY+zRj1gHSnMrNe3fsCut2KkDzYYXPofOnQPu3Hh0vyj7IzGL3hTd5PHGgpzCXkJ
RDFtfgD7u3Wp2swp1LDQyROWR2XgfTSJLm9+kz066TsDkFZTAyIPHWFmsQSGcCPa
OgK59ZIxBlUQi6RDLFywb1IX5BQ+jsEJGzDMeqc4N80LkGZvZDePEREPTEY4Ol+V
ye7UerQMJwgzrbXFrE8xRcvKLS98IQ03CPY+vlS2KVPXDFvHBBNJi9HwtHEuFjcE
MuZ8iELb6McoX/7qAXY1Cg3nVkQZtxff2vLHUO1R1oQnVLgkNvrS4WIOxDHXTC2X
FyLEyEhXb02u6pXRdKGTj+av2vn+GMPAc7Rl8i9HbevaZe26KYOX6LyY8Ob2fnW1
iT66VApeUarQhjyG4BOO67WOs86g4PwyZnjS9MUkeSizlYMEVYXRMlFwHCrjvw3M
0UjCH2Hw0aaBce8jfsOHS6iHKkFD8isaMbMP63AXmirc6wzsFN9NJilT9Jad/uei
CvLZVrMGsrYoDA1mKZW4HFxzG/MIfYrB4clcZOux/oBB8Gyv7k63NaUkdzD0ys4K
1xs5gkMb/2bOiGwNQZOSPOo1b6y3vkvOJIQLbNT0wJi7WdaF8lpM0D/1y9VUTTgN
tKzIofWFvAKF9HoT4TMB8z26UEL1xT6BnJxFD46rBotaX7gSSzvW321/UKw/3E7M
LjTNKziy4F53PDjZUflKCcYmi6Cb39tvqBH5cMN25cBHAozJn+YnwLU9tzZzHlPT
s56PIi9zCOICyZnhAGuefDs53CXCni9lFiSVDIGE9olKuIrNxSNO3Nl82vwRvMLC
II/mM0YGuiVbB/Or1f6/XdzXvai/BNdDskS16WKM2TbCGm2EQ5O/k0Alu0skVP7z
RJ23Y6aIabS48wqSmLNXG4fqhOqKSykU4OMk2d6OHj2oyUIg12Ql1seitKRhOMuJ
I6ZtmHkssxIj6l9jZ1hKovMEceOrPnC99de0CBmsRdeP0HSqKJ8DtQyDaGftynZA
C4tIO7FZbFC2Q7vaUrMF1E5h9fe4GUKBS3SITHjGiwHah8E/2oOHBbcxbJ5lIHA6
URwSp3x4+fqExU4g8UOtwsLhIe43U70t/nGgVhQGngvdq6AQqrtczhZzIeZqtCHH
gZTNyzvCGFQHnJ/MKnVC9IUIxrmWt7CFGHH9jKK9DlX2eucu8FtMNhVNf44z+czp
8p23YQiiwR39WV4LwwQwL6F5r70fNF+wifsAU8Voi/xN6DWXyWD1zLUNZk/+udjd
Jip51zs6224NZrQPYPoANo7XUcfBR/BUoktdNrJQwkq/sZGiDRqAtrQrrpuqAbzD
5kxCd51rnHjddXpaty7cfl6AS0czSmHxjkJJaxpyrwdpA4DSlxU60k8dLG6DYiBN
FMDO7YVaaYQn/WBUmJu4V2QEdCDuyxFJHZsXzEUyE+ROWu+ISFXzb5rYA1BOXP97
oi6H5Jh3cg4fo0GVnNr5tK4JSQz5obwJQZ/Px+CyBNAE6ZEzRlDlgEn+KdN+mOLL
NJ2YPahV1p8sE7b28WhU8BNpU/TzduSrgtk7yq3mcqpVryiBVmjw/9R4CrjL3QF8
8mzrUANinjFQT+Lrftlf/Zd519KZS74ci1s07vRV6ofc53EOurYNzwTsBYHTh1fu
6rLVaNF/xbFvsnbF7RzyHoSivqZnFevjuHNr+Fm56KrxVpYcmdjRvYGvu9/Nu4xO
/RWoL5t1JAPVZ4Nr8m47Vr8hP0JI7Ib4ledpSy93OF5A6Iayjw2nWVCpZpfk9UlZ
Xl0NinAyczPTPCmOWxGif52FzaTfhkJs3SWzPHIQHtwgq2ySefRHq+AEPw3JikhY
3yTriAspmf2cmBI/kXJJ2RmfdJgf6KnjUrEgPDhAxP2h+LVHwNWv3NL3/UfBDP0l
3E1go0nysIQGzwGviaEfvihbmPD/FmtOHABd+yNzlntkMo1VKP/09zDQrNoCQRPh
1jVHr+Ni8QUiIlQ5L5Qy2r8lQzMXgTDM/+L2s4BcpwdDyxSV/kNDKdho0Btyyb/k
BTZALN2aUyC4ZWp/Upp7MAY20v2ABM3nSd0WBajRW3zgWCZvk6p7HK+AbC+3ysjG
Bq5iNoWMEKxZsXplNL385xWGzc4DGq1gifpFkxX0bHaeZPx3BeD+iFjI30BSQutC
8eaAVS6Izm5mFGJY/V8hjVuQzlcHt0/mAoBgHlAN73aMnuZjltP8ffzOPRg8hhHZ
+L79NSF0xlasy3gvd4QZuitrOxsvleZUDaiShLHeiRq6k6cqwd3s54OnPMhlQg5I
j9xJwHHBexz7+n44YK+f9BOs2s0rNIXdCnWWpcsguYjnGORDkui3HYYn3eXcpe3w
YDsicdA6IzsOB7qoVqL2bx8VTDayllqFgpbIQ1zulDJE9H73ZNfN1v1OPaWnlmRy
ymoIGN3MNe7VmDs+t7kvKOM3Tfz78qT1hhYC3osfxlu6z5ganPs/EVMWacFQ9BrF
Sa7o4sIToXMttIYgN5/8cdpyXtQu5hGfU8HkrbXp3xpHygdY+lqDY53mncQKaSmf
aIJKo6tLlP5erbnXMTDFIAO48YfoTyVAlRDHy+x+ucguCl1UjR+xOHpu9efKSdeM
HW0ErjRD+Q+bjCWpwI+5R9XODdw3K9Nu4GGgcXnM/eAK8NP2KUh3GKIlAuLkIXQ9
mRZ5kaZ1FNnhoseHI+e+NTG6W5Mr+CWgvj5qfAWAxJYfD8Sp2QhIUDNCTtLTMRvM
J6w4XwbQpYr2qwG0J9reOKciT8SjocreVnqjDxsJBFudS8C4Vx9Xd0E+sBIYnmTv
kfwt9yx11r6aHiCY5WIxg5v5et5NhjQiO16pyg+TlLwCjfsO45CS8HVgSiW/z+Sp
IdBC6BaJ/EHfTad8DBtU16mOX3WYSrIWN8tpNCwlDhk=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kv4GCNDibOGW14S5KZEkMqAj+Irul/jGVAtfvX3G1vZI/QctGM8ee0fhnFBzPx66
yrTMxFX1nmyVSsicp5tYxngm6NRp0MgHslFJkEsdCj+VS+ZfDpoPc56rNX0IdP4o
KFYnysljKphVc+IUvR5MVHgFEF4mhEN/sNsbUXKk9LCP0/2/IPAk1zSoDorGelPK
0vWH5WNF8EpAQHVRubdbvKWfC3kEj3DddlbVEh41hhb9wMwmeUmMZ+QHfjrM4eQ8
kK6shuaVmHxPj0AM9s+bEoqJIYNOxNSOeaz/hPGTb2KQ/E02mmTpe91MkFRhY4nN
aQtHJ3ZK5hcJpQx8gOVrd3xV62dIiWnOvT3r5HXAv0KZUCGzVg8pqo0EYQc5YSZ2
WHvrwaB5CkmMkWwr1tJbUJxQeArp4HQyGZykllueAH/BBpVKyLVfBTmcLY0LV+mW
qJZ/SD9tXvlJQvP8WgUGr7YaYnaudjQqpBVz1HvW43a5EYqOMKe/iRFTjxMtVmXo
LqwtO1pYnoPNDwa5BLkCNiXDNTYVwPZVpmYFxIWgJbth+Xhq53ck6n4wP9OqBECS
vMsHwUKSOWKN5S2hJOV0DHdhHgvuePZYV+YJOhGS7efK4vcLBGv0JqBJWm3lZBKY
O9ElR0FmBX5Zi4tAuhovuGmrmZOSh6nvizgpxuPd8MNoDnXbvKZhVnbeHBBzpkxO
mYUxzpo9CSdJbaagw446h1rfL4X03tVPNruaCIDjRavGLJCe3fv95C3lWx5VTl7R
L1pcxNBBjh5qo1MUruEk04qU6c0+a1KWgu9cGmnj8pNfuVrDInmTs2VkOwM+eDyN
Eovd91aQa7mSr0Gkf3FClh7SGp/OHqYka2SZCvC1JaMo1OMeS93q3s/VbaWTxtnn
Sr7K3dT5XjlNHWPg6fHlMydZvgfaRsy6bnzcIzRGJDm8cXQp9i59kOhtnejHxx2X
5gbh84hdysaU5JjAjJiPsxwejpgMMqpn/xXD0RNk0ELZr2MC+PNqLjEBz/E5eLqH
5cYf+NBI705UyKilpxlfvrdQ5o1lxWUjOYMxmliqkw8UmOesUVpBCCfbqOQvYQJi
EtsYzVrCVDDPZHP+Fh37857kO1+TCLTmJ48kOCDrZJNxsAsxB98X150aZ5bQrpBf
x/9d6q2IVep9G7XebaBpaEnlqjadnE87ceIGRMU0oAT8KVkhknq1dJa137Tj6fYo
LVhR2DYE1erm2mpSPoxu6aEHgsD+XwVWWtrNXKPAIschfoEuvF1yrwrvV/dcygTn
dMeK3zuZvEwMvKLRT3maqN46XlQ0ly2GcaSBXH0lLEzTuMnbocTYwkwMoaTtnMhR
603ZTPY0CyTiYxhHSQKp9Rl2+Dqxe4cL/8pt/PGhT4veAB3wZaEo+LUylqd6TM/L
XORjPt0593leWOuujJcefi5iXoiRSi7wY2K+VqWnzdRHnzJGnA+FUjoQITRSAITy
abMC32yckcMLu799Clb7MC7mLE5JAofngA71uVbBfbFcAgItM5xjvR8PxnR3PvLB
dmZioGWxu+1Tqm/P5C3TTaAEjklNP/8I+aJ6sYDU52TIVvjqIh9hVDyliR1817d7
xOrUm0wUmlhaDXMFe6sWn+nfOnxr0x3EcJ2klw+3gRPxzkMP72OknEz//uTBW/vS
VdvrXbyceOZOfQC0vXND/g==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0GNS8ERjeYwOiqLlOp1BR5PY2TOuUzRhw4q/+lqnofTNOr4oioKvhLozEt7HLAd
FKx9ixDponE5f5nmI8Ey5oyDB0MbXClGzVG8dDWfRkng0ujkT3aYDtU2SH2yh1Pe
ccUuRerLQq2E4B4WmUHRZowML3zGTxW+OAapcwtKxxflypYYiuirL4o3qUQWeU4M
se4lSBDgnbEQbIDszEvksvf+FXIqDl42iQCpZxv/15TmMtRWT4yR/c85MpRpZzRs
RUosTUWQXBeVHCCZ0amNPgVF33WdCkDN9zKdEahfGJerapHg873kiXmU8ZXrymaw
UiTG2ELmUkHHsjLWVXVMT9/0oBIuzwxpY31u6zWfjg9w0CoJVADve0U1BpQQYNwq
WtcpzTwlmxpPsOnEhMhk62ZvZJRn8SUV8U+ny2PoRH3vOJo8ddNzlzRfAudi0HYO
GL47dScGLsUnFwiWdjLZDAJ98mmQoKjBD8ncc8SXBR2GSTvAY2sKezvHs2NgKB59
/1Ds/SdoATklghYhNXHF4ZmAVgUOIQu/sPBvxUU8jfrZX6ycUvy5RCGFkYJjX0tt
dKFaNT9vVUwlXEFr8kaeMgTZYIgl62cJuad88k2ik+tGroXs69jkeo0NCT8Yu5t9
ommAcemA/kDj3SCT/hmFVdKgcRozv42yLWLhbIvq31EN1gSBtsaYJWt3L9wqPaCe
5TIwHFVuSwNGYs904lrGMf7x4+TAq9S0nMWJ0J+VASNhtgPJR3SDEwed8D/Te6C0
W5Z8ZdUaH1I0/f9pjGwmueE1Fj30KPGreanSJYMwkGwNr/jzIYrpP3qplJ2nwKZi
XjFDnPq6AMRxgSo1A13Yh9w0sJ+4tKynwEuLChsxBk3wZm4dpX0SKH/9wlGlEQE4
LsFtHivLdgjDxQ2shCK0qLrdUp716jBqfdAyAzJ2J/WpBhRC81Zzzd2fy74hactX
nFBpZMd9wNhXIrXLFQ4/qT9cJbk3nqjOszQcfk41lJaYnVfaxEzEshwNjDC8efD0
b+p6Vke5t7AAESGYIoJpAu5k8h4RDSXt1rcWhwutZkfMkEmbD2bdhdo/jKQxAI8y
9uU7TGLD9F/ZevSi0iBCBDruqKF4uRrJgDghY19xEpjp/d1nx9SOGA+/31LDiY/Z
/bq2UIjfLDRCmRmlVo2TmERxbDvKxStDcwD0FnJxX5jUGNOdI0FlYhH6aQtJjFTK
MVlPtjvtk6eI8HeyczBKV3sqdXixsfX7I9dZR4/S1LKfgaZ3G3Jmzn5NaurVwEiM
/JmpVZDQRzvrgYUHP6Jld4wbIWDxPjufBmVjJFHRXCIplllbFpyuRJ0bHywTPbeb
6buJt1h1WroeJFPNVn/5auy2Rds6P9lr9m4UPbrV9ApQtXb5g+MKqkGW6e3rqQ8u
m0Mc4eUCN2qfHVjEXvCaBZ0xJKCkfWHKQr3IPQD0dyqdd4xvMmQ5NllIlQecYAKX
HwtUqFyoPUP1N46MUjbWww79Vs3W2+NpIJOkbKrjHgLB1kQBgpOx73oeELRyLUDs
Z5dgXsXmfucCruP0lG40WXQPvlra1Def9A42qomqM06zFZWQT4ZGc1BdK/0qA1q/
cqB+a5OP5oglIsei8d/iERaTE+7lZgvAKCRM1CdButXfUhiFC03jnw6zVSJDyBO8
pAhEwtPZGs3PdVTdB6eT9SEB3mRIGGeshKPTMFICLX3zCNHjAEBLG4clA+ngjm6W
rpuJRSmjqObkFMBnjXtKYpfB28mJ8RUJpyxXJcYGbJtbLgdzpMVlMau+Qk3WYEGF
s0K86vTTNztplqgQ4wZIhY6sBU/bCufS+cAEC5/j5BZqTyMC1gojY60rEew/k3/5
GV5vI/6dhRumsMN2l30nTsO/C42TseiKAdvnDpKal1FaY+N8dRxoL5GQl3ULTyqn
VJJ7pL0h5mBKtJVTNq5EFdoJ2zao2Bi1HAvDfd9dzk3LTpr8cd2duV8zZ1a3Kn0e
CS0hBuGlsTmvgkgoAmXUvOhcO6/d/zE9y5fPUDjEDEQ7kXsKyXNo6WEl8Syc18Ob
L+WMBhQtyrV6toItubN4gUSooNYoRgJa0z/ofJwMBEfxGvmT40asiqnIa7keRfzD
Nxr5+68b5pYAPvfUseZ3LYRUhZ+Sm9sUryggU4JsiFbnLzDnOai0iK7UqJ/rARya
ZWEYt476ueiCP+Vqz2OLRVwavN+00SXyCgJWB8BxVR7PHesfYqikwrzIH79ZuGWs
EGF5EzTc0GS2t3Eh1/hxHiwphIn+6wPp3xxxNa3ISh/rl2+2hB3aHtV1f/T6+Qja
CZ/ZvaOK4tquuhzbmjPa1gQxxyArqdmBdznspsI5ZUJb7eCPS6Tdnv/+R0dmDZZ1
qTwi6t+s5hC5RRlq93iKlYw9rzzxylQQJBUqih48m9pwo6DdQWv3llRkfaR3ecF3
mJK4BnNXsjbPIAQIerUSwbFo7/44WHIOoQENjj5UPBzhi4wBc4TWZ05tF6Fgi/cf
/nIEz7PIW3/LbzkkWyO8ZAJiy3hk3SjaWNJjwOukSnhd++9plh5KdhiyuXI8hC+M
6EbMRverZ4bUEzzxn+tP3EwZygHOvq+3Ur1U2U4+OM7XA3i4k7POvmF/C0gBC4G4
miqMfZFpPKSlNQX++/AUng==
`protect END_PROTECTED

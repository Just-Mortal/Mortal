`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZilBxBjz8F/zFl6+DkfDuUaQGbzXe9vbVxQ3NlCApxuhx/SomVlnOAEiZHE4xPU
kkNh2oSWe9RW9buCgeMOxGTs3/AUNZ74M5pT6UpqVVjbH1FuNVbMt9HM41j01PbG
XctCUKhYSK8Zd0GKGEC3UCZuLAfJNFGvmCytVAFI5MDDM5e9ubC6VHFusMfPi1mZ
/zjrnwGEdIz17hVqYoFz6kKbxi/eO7JBXq2B8nCpUfRXgIqbAw0R2+vZbiSK6lhU
ChkY6S7f+NagLlQYCPHQ4BHBHguEzX1dPwIOgFNaxMj8hMG0AdiVMacjFXB0oNe8
hWElpCIXS0l/GwczgSXRCBwSfEM3bRbMLheFPeuhu43KM6ngYrt3T+dowwaPFjjz
tPByfewC4eA31ISdA1UTStjclEv21rcNDTbinvkg06HiQJkUO5gjOYOo3Q9hAcI4
Ct5Z4rQ2pjZAt/+x69orz/ltOYhgopPTbYp4AcCiY2+VweQ4oVvLbday63hyA+if
QxbWPlCwKqjtk3fwgFtDLenfNYz9mqN33I0+jYhqm9v/1NyvCzri2fOw3CEbKyPA
g0VLdxBdkP/1UkJi8Zh3GCozAfXF8DyTP9ehFcBT1KlubbdTQ7y/iaivfUrY603O
NgYYvPOnD3AzZDiDYMcHZ40mPETfMNai10RODQRC9DAabaXo1qsIJO5rAjyfm5O4
P8hwiZbfNI2map3+Ok4zoQk5o3W9sr+uMBG04PwxKSPzQlJvDPbzMq4yTEDkogds
u7qxbj/gbZoZdp6L8epflJEm9M9Fk+BGVbpU/UX7TmHKeyqLnwflPDLw6j/Dg7Nu
ihu3wSULNfNMH0u8kNKcvalLgpKNMeFIHisalU4PE908C03OJOZexaLwjNC6pRp3
C3DoElb6wI1TF8HcOdCYjAsqqM0ymltmKF+kiLSsMNjssOupKbSbvir8pd1isXkC
bmxIbXNoeVsTJBl6dH2d4MjkqTmFI3kznLy0L5OYWeKYCyGfkBYEhqnpcKDgZnep
4LUIT9nKNXvwX1hjqj2lQOK6FCX7+GaHNi0gLP2z0KehWUj6A3xeYB8/YgjGMS1U
knO060B7mqkU4cMPtMtF0mxxsyKw7Lvg5KXOA5PyQQNXl9pHQPBC68gUDv1YciY4
F1OIx8Si+IWcr4IqB9Vzj2jr2jcc+Wbp8vsx/WS1cIwP8G/SQz4uVhwmWsNbLpjp
yj144w/9Q/W7fiG4hBNXii3HEYGobTb0UxoPXdK9DifB/3q2YhqH/KTDOuSvWceW
d3Rr5UIfseSaPEchpgXH3EVCkWzrG7Sy9gAFWHwmFJSP4U/PAnoXqv8qt36MGst9
tidk2pfMrAn2mh4NRlzEnSxSVhCbiyP9Og/LREFJwKAgRyI3641Bc7s2rRRBUsjd
Y5ryWcrHWHI6e/K58KMsUfUwJHjpHdmPnv6Z97qCfNwoyziKYiHJ6QVSMpjHCG3K
yl0c4B2QxfJCLytOJCFAfUSgMhJRiW4Z6+zx4M2CbcXC0d88XVZV/KfzjVCgj+hI
8V0Q5/aziYnP55Jjom/99iraoWArQHLPd6FsWn6p0o0yygS6ww12LsENNrxOVwvZ
Zek6zFsrKg+FUieSmsRl6KDXqBva3Qg0wRJ6bEGjEenF1M3/anFmHEmPvw0brJaT
9/1a+7pBQjI95fIsnlmS/scUIBExEZSdAGrqD5HSe+jXcLTHOir4/1fc+RmP1b8B
INkT0QtuGbLE9FBJvj1hhhYlctGCTtcj9kPEDS2O5++nJlKKcP5uZV+OrT2JM5h6
n1UflQxHE8ftMnpHSfejTkYtStYeVLkegeHunQz1L7uVHDvu/35YVOScWIzefNOY
KEEJ3lSlTO7vNUww4Svs+J4AI79ttnmhkzhlJ7HmPtrZt/4TPb1vsSSaN9MblLj3
q3q6YL8s/2qDBpsg6onmY12bha3osaMMK1PZ6OSBgomID+iD043BTG4SxfDJU1iT
0uUHkCw9pcXJDytpiy2+Ed4sF24B4/LbGnarKNr+EOOJJh5Q14w2Do9hWldCdTbI
aBeXL+CUkpdXFUIKrlm51EjOdH6FBtqZSAZR2jOiUMwI3dp6v3h+rs/n37lH2ZBM
t4fH5253YEArwkmPCAG617tp662KlVwA09dZE6R5wgTlJ8w2rbzQqWmGGouivHip
TJIKFroAXRTI1Ol5N5PaNFGOd+sEf4r69HOPc7EX0lud9G6V8myBZ7a0ihFUonLH
q3ZZqvTHT+UhfJKp0DAMFgeT/+nkWJPTW5BCsr+SGnbXoSSEpd26fGOUz78zEWgZ
nzYCoRlziSfFMQdtpXVP88stcW36Wi2OwqWztzpETr6nSPuWBIvQQlg3/EM5Wtjr
nSvCUqc8QJcYA6sOwG7r4cSL7C67jxhRTyKFWcPtus6IHJDZVENjoyZFKf56C9JK
`protect END_PROTECTED

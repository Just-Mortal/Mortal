`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mQKz4yOtJM1GivWVBTusiBJHp4VfuZG9Aif9PNsk3o8cUw2DGaf6eLLTaDOC35i
ZJbqdL2bNr14jxFL5qY0n2T25u6vh0Lzo7kIAVVLudVrIZ3hebUwsuQokZwDggPu
bAtmB1XPwVLTsPBH1BEH7gy6kjHmJ0Ynp7Nm20Xpp5Ub0w9DW+BrySlXeyaQo6q3
zUJGZQba/61ZvXEChTg3z9PiAIO1N1Fb51kjYLGGj98GUOn3UhSSWkZzgbBIC7Yk
XOAqY531BO5WKQYPw9/yajmV4QBxgSMKjRS60i3Bcuvfyka+ChxFlz3IqUEVdD44
oZfJHrGGQ3pEod6GJYHbaynKNm8hpAhV3SxCN7APFVzUq9WMzH9AW38lkk7sc5Nt
1fMw1wNIyzhUFUZQWLXSOIrpq50ej+jJA8rU5XIy1gaj7jZE96HyA1iqO1LSZRtD
apbUKPuwZwXl/O1uXt5tyhKa9Eb9WoWth3z6hBvb0L2UngE53qA7aldBETehz1aN
3XukAv+zmxzMOUI9Oz/SQ8iHQtnTcn69qsSyf46vAXZxPGc4yg7yAw0rSR3UaDHF
097ybyymIadAy1gdbTClJ7kacfrFNPizZO1r+QZGz9ZqWW6+zGi4kCm4oEtd8AgC
T6XUFMgqJpwrJ8NyTnCXN2m8QdLgc7sjRn0Qa1ZfNLkDsrNJu9fJvL5AIVVRX3C+
zdidNWO0fdN0WHx0dNyQmYk3ea4usnzRqATsCot5gkyxs2sYEDmbEVVeH+9SPyGX
TlT33NQvYEPKKRSGo4iJJ5ITxWTH7divBgR2PdjoGQy5x4h1v0MNeqxF+qBR8VxK
w79ouB6p+0nd8ZaMA1S3rRqBQCqvMHxw9TFLyIBv5Bb0vDjdgnAWICR7a6aks634
lx1FoiWqXI2aPNBReC5fJQCv/bpV/XoIs/8GBYj11tA=
`protect END_PROTECTED

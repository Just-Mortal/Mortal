`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LMkTgpx7E4ZrRbFC3Z/8O7kFlUKkTCF/funf2DUC+NoZUt2x5y1yVXnpfOTmg+/b
1MjrVBOpg/NBX38FWk70X1GIq0RefuVGJ7lpPW2FS2QuAnwOKTzOZ6Bnra34C/cW
a+hmSL/bWih7e/SVY86jxSySNKGZO4KZl8IKovu6gBxY7Ke+FgPfrLs7KyCCCCB3
Di/wMQsJ92Wp9plAFlgcbXcCvAThRpFalKAwHWfddZGq/qrfKt5CdmYKt9xy91sJ
SHOW4M8e1aRAJ0qRN4IdCiY9sDjw0AWz3rY2lpL1I9cOvYyi+UmaqR3631HFA5bc
sn1WcuaC4WiRnvstga1HWxFiQ9ywb+gFgAYYyA0eXR9+rPFlwb4FOXtnHsOoI6EN
ZyyeZ4J1/q4m7662YHOB8KOc2i7F7hm9CYyT5nqZYaeoVn7eXLiMswDWJQ/KORK+
xbpcvwoeRdkE//2taEWaqVsZM+XeQvUBGi/L70NOycWWBt6rX7k+hx/Tmv7sFJq+
UkWsMAAc8A4i1SmQU49sjmRn11eTzBAhheyfej3YXWjURK2LiR9xoh2/mMsKbHfW
niZLB7OkvuczAaw0wNwCudQqaulRVnGz0ipghGvSbO8+cHSfS5bVL5a6374V53Pi
2MGiYGhQYBFUowjRI6xuPL0KkbBy0GzHIQBgsuA04iPyowLS12AK0Pb1uLlRh/4t
9pUDy28AQTnzW/lOy+pO6tcC+lsEZHfbdnCjUJ4Avws5lQwSm0z/2Hs25hn+7hSB
RHTP8LDHbWcguz4Kie6j8jvMWvKrn5oLY6xuNBSsfXeR+CnBtKMWlSxrEzV0Z/+5
DxH/tAiJwAOZRT/DHd4hYmbN3HMuzaG9HbIIG2FfJ/cemAmI/OukKjfqEUCMzMkt
drAbs1k+VIzBM8EDlMb8DtX06UVqclCL6TYEAl/ICR65EgoF2L4fMJf1ofb91lU6
yoBtXvpQxvzWwCoFAjYbvO1rSJr4AZEAmBUxTkHTZGFMjRUzEgIK5/I3wK2vvcxs
hkcwE7Bhe6ATgxcQ4x7A9vKUp6yTfc4lGFFtvbCBRu6Gi9qjC88LhvNKyJIRne9V
hLtjyDyocUYN9T/L0YQ7Hb+Qs0qAXepbb12WTcQvlXDDArVmnA4RZhWkMU9aBXHB
svG1e8azcxt45t27Y4VLe7nOD7ja/6Ee06pfJjpRP5HVwzFMxUo0TLUlo0mzUmCP
0GpxT3Qcm6kKMi22zcjyB4pacuBGe63513YSVbsFBOlweKwfLUAGGv/9xGlrdifc
PiKLSnshW21bIoQnwFYrZmo7Vdhu60s+XPXa6NDj8VgB/Ehv55V5nzLn1T4P9LFY
z+g0ZwtcnbeAgInqOg0lYc+o7aFgsG9CkVBXI7wTqKgG8OdHJiSwJRWByQsvFQZj
WtXEHaH63/rtzT7yL0O3jgTVfMbNZtOr511CCEF9kwkoNHb3ofl/4e50T4kTEZkv
CXij8Z/98zaTgCzJkoZ/mPGkR5rquahjIiC8CkFk7gfSJDSJLJTmtbp2bqG30oMk
`protect END_PROTECTED

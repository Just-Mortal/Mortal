`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjMdlv1CRmTonci6zR76SpUZURTN99+68xdVaEqNv2gGi34lAP9bbTNbGebEDcQk
TfsQtWUbr852+51bEEhtSIMp/vOBWDGYSYHVr6k1q6ovLVbTJV+1HFY7rLSoGXp3
inwI4uJ6EwEovgXjWojDsDp1rZCBGAE2M26sdVBqd9ttt6nKa/VT+GJ5fV028AOf
IIc9gjrHYN8A5mBY+9y3fHmo2tW/hpmARdfcNlxyMU9HeC9J0cLWc/gbMEi4HEP/
i9b1JZNDU1wAcZJBnX71HP71LP6QBKtLFqQAJ4fvgROaHCp+fdHdLI2hYb16o2Rc
21yZXwgt/JnYUdl4H73XhUkV8Jz/DUhZ0WkwzaLOkrWDqjGBfSuaWS0MJz9vpWjT
/co7wazzcoTXgVu1jlD0jvi3X+7uOJxjdB3ZQz0nsHDdC8uMOo3HxdlKOW6a8M0t
LouhftKazuKVG+eD8wf5GwOKXngoBHiX3enuv+cLFXmnjSt2rBuX7rtfSvm1iDuT
RCuzm6EK4ZwgX2QEXPAV5NMtOEF59G2gq22EYfvf/3Xfzxpuyy74Kqgiex/StRuK
tbbL8szLUkFw+JAVlPezYGs9aPI34l5zK2LjkvQIfjIbqB8FOb/f+JKzIJ1PlR1E
tJ+UjLKjKvsHcY+8YKAVrcQ6qbyyhsj+8sk/rQ9xwfbhWS0soX1KQlrqLalZ18Ss
MYRQHgOrAuqWcq08MEDveN3i+g1/okRmitAXSyyuXjln1w7FU/ZAZcomoBvuKrQi
N4nI6rPQX5/T3UwRl4BWHLFE1swkEY3rgtZWAZwOeqm164bJ9vouvdHMLu9yss/1
QUT80fl7SEHDw3gCA9rOQ+D9BBeganepJ11aZNnA8bw9Ow1GX4t1/nPf04j2rEK8
DC5lE/cr3XADVLRqGk0CI+mrJbImw1hRUcmHHKPYaCrZldPbEg3+iiLCiPORKOPP
kf8uxM2uyYxPH3mO+5/SqloEoUCuI7J3/EVfYndywPrib8uT6O5Ub4FfQHmnNTBz
cUCfg+qP/7CiBFs7peU9k4LgOWg9+YJHPIXDjssXZlTucsjZq6AbG+dYdk6H/yL1
BoEAFanRzRDti1bNa81BYt/Y/EbZbARXCce7XLBdSQ4yu9Ess91oI1jl8Lo0aPn/
1aetltHKCz2sl6ocsrCuV5Wag7m6jchVt41b0VlVs1dqYQX4j0VZD1GaVfr56Bps
3g6i7E1VEmiqS2EwQ7fUFKEk92t4Sqpn9kBEYhfnhFkyO4FErLK1hB3qkeHRFkeU
Oww1igGX9YZlGxSeDltrW0CwLDJpsFU2O/OWq4j/yrBsOUwD1s9lvRDzu7Huudaj
cOkBD/o+CcfDqwzcTzoxXYj2jIoehcowgfBSSdp2dubzizjMwOVf567mgX6n84aP
yEnFjNWpZw0qXl8ddOV1DwMx7j0euLkZ0XkL+amuMs+xERSWDr6BAL/0hECmVzbS
FoOYe9Oi4UXOu3kaaUVA++1FocFYxFa/GLxxWsb6U1cfAxpkIWgR7n9sJnE1DtYT
ih6rboZ88mrBLizUBIdrdt2srGN9Si6hbzZwVI81iXkE9lIqRhgRdfttw+d+Denf
5Ebcp6zwhxUJuOpGEfQNanxYFSCVrLP0B4xT1JpRB86AjGukMWvrAkZ3I1QGDDHg
3kWflXh7Tgoue2CnxNUmh1HWPtpbB1Gh+BU01fF19FNBORKPJMOpmrBY3gsv6FLR
j6hY6eD0O8iqGtCPqpJ6hGci/Be5s90LRz31wD88p9JsMx69y1MBL+3fzFvGQn2/
1N1e1vDfYL3oq78fNhR8E95l2u6Fap6nSsRLwUUFMFdlt66wds/1uzkN+FsIFIuT
v9hkmB+p3im31MowzEJyYjnCDQaTC66JYFbhlKipkvxte2IieNuiPDcDIA52srK8
ele1bFAWj3rMnqXgWKxexrN7v/VwZqsjMmIdl+m7USRuKSWE+Ucc/tZTV6gnEow+
lDZa2T+zWz3AS8FRPkvr0UZODzayit9aDQx8u8K2UwJKccn0ScPeC2HhsWI8lOHD
r+2e/wtmyF8a38ckUHYXwIFJDLzo9g8S4bpwipLzDYgcLKSG3MM+oFdeQmH0/SLZ
910PQpSSaFmFUOqRoSJ8s0lNM9ClYBTUa7u7N9CZiWVw9gVdUp1fwjsigAf1JFHy
41Ok4jdU4CwuNyK7ZREkY1NjT8U0xWtEqstKU4jD+8jV7Xjnye5jjfa2aRoYZ1ka
Arm7oRHYam3gY/bsMRnFRdWcBlED/WtpWCqDQilpovvZKPCAtSOW0NcH1h8WOSyY
onwyOKh1bq+60baMGD0l17pdRMS7+DHPZlUSki7uhFOAcUbZGC9GM9fPStruojkS
oks6KVyY7TwwjVRU+7w8ecx0ZRoZjvkrwIPhz3FlxTDpNWKvIb2FiId/IEsIOA1g
n4vCcyPKnxumLG5xzOXUwObTJTR/tws+8YLyhe7D+3xFC7WZqwz1mHnF13yXV/oV
CiTUsWi55Fylbb3iSGn41SoCmjdz+wUkrLiWjCxxGKGivuzbymEJx17ZirEqNoF1
r6yt0L98G2X7rE7RLuBtFaPOlkmItp4k6g5WRqgcc8UMnNlZS4+oj4a5oEzyOTlR
mLA6AmvenhJieIY+aN5EK2j09OCZWwivWxfAlBOdmFZYQj1388utItJHz/tqSpEX
3INER7pE2duQnv6P5s2F1gj8uKuBB0uU60LUpMNIXE5Tps6eLvWS1LWpLWxzqUc8
GQajVUUoGIb8JIP4odiQdIMz1f9iA1dI51tuQSwq7fG884+Cfr+xAiSY8M28jssr
MEpIo6mjJ4YR6wgaagNwJSeT8wSSByj/d1s5lwZ4jvDflO3ls2+mZHjJZ+nLuof0
bu3hOiQjGWJxOIrwrBrcGKLVitYklDvxuZALI+v5VBayZ1T7urJB1qhfDVl785Ec
MgiwnJDBoCZGxi48nN+eKgp4N4wj3FH9BGM+0LLHbEPGq6HNhGazVdTgXhrHp2Ik
/g5+cP+g6zk0p+t0ipGhak5JwElQuah6CmXjpBps9i9QUv5nHZLbRBLJCee0Jots
gdAHYjt26wUSZ/pSqq4E2zIRsmvk4aJGab3UN9wtBMHfFVIW5mkydBReg1rce+Ti
NYmIrTqItdfO748kpE3MRS0tVL5FXwkTNHkkrH5n97kGTDvdqAk+iOGlBVTs13uc
kOMBw9gkQGFowc7/hi7GLmxFzNuhVu9CBrUcg9Sc0uEeQcT8DPPERb4lopCXKy9V
8nei5Y28iRW8aDcJADEajzALja3wwV3WReeaN9Mg8f++gdhdCOYv57jkzAs3+2si
P7tHJvvdlX4Wqf9NvL7gN2ln21oFmKavPV54xrNSJgMNcHYGOM6xBmi5ZILKFLaI
iYt1l0AkKGMVujSrH42gPlnkwum/rgnW25UkFbJItq0VoYXFCETpEMCKwRO9NzKv
0aODteLCbg7w1dEOhSUMnJU1EXUEMrluGcF/SrRel/nzq2HM0CL5V9lhVdxaoNX+
5CmdyDWuQIvPgrOfPY6L50svJicfEawa22yfKbwmxSEx0SObDifJZtIfxIqr5we+
LjNEsh4MnISj0UBKNUnogT7+LIG8qL/T7yzniah7ATWt2unFbAYOhTgjeHUZlT9R
8HOh3AtssnKIWLQT2xGzOSvgVZ0YLBka18YBNE+5t+W+A0urLGjF5f/S0zOjie39
b+f0M7/DZ1/x1XYkaIkFvVtnsCR5z/y+7OTlQREhXV4GcTH75Frbzps64mr9QEuQ
ZstIEWuwnU7MCcVCwJFcUFmp8bZJICcK5H20zL8LClH4FhwVJo2INJl98Dzq+Hc8
I5EFnZv/XEEIge2/LPylks5NvkCmrJ6S5+lbmLANLRqSEPnky6sOxJaCKoy5Jt1g
HBKEBXV3xLYYrvukIpBrrEFyaOf8Jm2WNDqzXoNtEzlQ7NkkhmmLMVPWYQScTr6U
zb1RmQUJ9TBKrNtG3rIsSEEhcSSEzHkNWajPtFgUIF4cvnDlUnhLm5qyfUo7EySY
GWjkch2Bt879SO82W95I+Dv7aOlhCXEgzcmhAUWo312m1FWtRL3UFXO0JP61SaAG
NC6vgB2P81DDVpSybUoV6kXKtjGIZZg+z1vwFPaYCKbR7KaTg/PXeEgVTGRO6TUO
xZm24Ti9CfUvByVZw5ilya7mu7GcBNtaZHPibsGhUN842AScm8OEzSRI69B7y1t7
ruYQ9BxT/3/zhq6O3vhMMleyVKIufiuS7LCSnG6x2/Q8sWy4FhMctQybgmABSK32
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZPotwHkbRPre8NTI015C/u8gzd7rrI1fdLTyHgzAGndgBc5yY5EciARso7+v+R+
Bd37eeLNm93jfn0cjQfwLTf0/XDUeAEWQbHN8ezEwPqDOkvRye65gaqNVrvQ7P3P
8Mvte2obWwRDeBcITlPL7L0sXwWNGmqY3gZLluPAj/32PVprmhalRf9y9I2YP5Dy
VK1AogFQuO9vD3jNtYvcQGNCfanNhptPe2SPcB11F2Kdf4LKUtpCGjtO3GP0xwg0
cIn/FZLCCrt8XUBQsBl6C3mXtrx00waioCW15lucvBvfAGsUYp+BDeGDnwFsXtJR
wyZ0J7QxwP7PFNpDsF3neRkp/BmyVZET2Mb6iRwiZlvyZQH/hNOSQM6um26CdNdm
X532xqJLoNttp1eYQ1Y/ZpNvGHu617LQI9akgFXFApM/KygPTGdlW1J63JnhM0Fe
xZWquDwaK7aO4XKpKl9RvlL60GTGMPFeIXc0bSpTWz8YdWFKhQbh8TftVrE4WboG
PvEsTfv8hVCSwXiQzAPmsCu7JkSrK9hEgOFT/w4rTavzzf8RXeoPMRodqsrmqQV0
C/ggESoVN5gfXqW/ZEeo8YTYaXVHxCIWx8YA1PDc1nIbqw4dQk85n5j4M15p7mt5
Z/auTEF5a1hb3bUHieowBgQOImCoBmg9AIzEAnamSBIAZbzbNOs7AlghOvsbwYrf
5SyOP+NIF0bVimL0As9aF9zC1tDCG8vm6MFBibpzlLpGUi5NFeVA158KI7xI57zw
hQ+qzCoeYbQUJsesJAJeGOGD1CEt7t7JNqTDbBtHsWWyI5rV9mjT6aAKrTxal7+o
anfnuzzqsMyxdAgPeV5eJr4g2FsggtcWEjD5V/28Nb0YV4z5tM37qDlRFK9C0HO7
3qgnAmLuNsepWy3efIK9RoTp/xrp+JWAQsjCqpdXa+vY/eLg6b/hBwhuS+TIYLdE
MbCwqZPwgiq26W3+2mCznIjgII3oWSx+Ca9u/7xT/P+dWYzFUCPlPa7ftfnZ81jg
TBnmwiPRSwiHds1ddzcDMrMQ6gvzJSmygJXFX8f1bq5yZ2L+XOLM+Tpfz1CBtbXe
4w1lwmrG0xisSLacN4NQ59mVFtVZZInV7DTh6ys5V/Y=
`protect END_PROTECTED

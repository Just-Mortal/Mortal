`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmTyk6raRulC3bfhDcIoiBB7j9ypP/rPKcyh12FvLLRMrVeFKUREoCMfaORtkL4P
C2SuZgqCv58JkfgK+AjLHUVNt7Zti95MJYfPNZAE+mo8185nT22wRYORkR37/Hyh
Fv+IlHIYTtvaS89sVIDXbG01Zt1bLG5UmOAsppOYErwM4w7d4yuFOdM62Oqr2vDz
hTNEforW/aGVT0MXP1P9C4ogwexQOIgQq5QB7XFu8dlH3Eap3RWJRzEu80Vqah5r
ZXM6UG9MrX95aI1aI4y5Eo+j8khJaCjhCxuHcZjNcACtxdqL+Jnsyc2MedkKtm30
parN3gTlNXsJwZtNZkmHLgCyQe6OPn+dMP/gj6QGwOY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9BsRxJxX0gyyRHN+8rGiMQGCt1RyN6HiybbUfUHjMeqCt76RjkMIE1BIOy5HQslr
IzlbdjE0mSWZqZ5sm2PZGcdztAF7frDSknELT0avtv1uHnD8mi/pNcFWoxlBgQUq
gudxdhNTLy7Juhi+6GDbdx0JShmGt/zqmw4Uh1iyGvB0FtDNh3gH0wVPhpkJgoSR
Apv8yywZaVB3ZXByR9t1cgB2D+aipV96D7bqhMMbsAaHFFsWC77TSCGgyQs8tyrM
6WDBVjH9pMSqhCExRmnTil+HebNyfh7RnPEXdCk13q2tjYDMqAGqghRtsKBnnYBz
If17z6sTETn7G5RRutdmB5A2QwUeb8IWObcNumA2d4Rjg/4ZRC9x2b4frE+2VEC3
0kYjp3nL9VGtyZAwTH2qVI21KgyoehDhPGaZCK1DqLQuqppCiDiOsRB2Q/b/CVHL
4ogxDcen6o6FVTXOgfQ0pf1jiRGT6fH4bX9smalETh7AqlKBocPLezd8Rr1YaDWL
d2dACuzmpT8Ej1VCoDBqWk/FySlafN+FydEQlp/x25u2G07KG+5XHlgM3o8RG+8W
JSV0T+KTruuy8ijrGQIJib2ohgcqMOrPvIi0igyocpHt97nf+cVEVsQk+1srDz0e
8IEXquOp5joi34zoo9wE/IR++0bztEahbhN/GNmTeD0FZcbWR1Qoko/4bBKIjf8O
GkYtby10BxsG0dgXHT8u0LC+wEZpyITSspinJaC6RfGGNZONLUnfOX8SdxNNXmoc
/XwpgWLJyb8l9Vglpr5lHzGmppB4j8eb70qKbYYMxk8=
`protect END_PROTECTED

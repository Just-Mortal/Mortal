`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1cMKk8YUm6Vr12ZHwuDu4aXoc5vKPj8UmgrGTuQk0gfs9fx8Ep31p9yCPrnGzuYt
8ORc3e8eydDSn4rzXcvt24xwUKHcgXOAIwZg58cibVsCKOZbtwyzPXKK8k4gG49w
Xa/+KfjCsH258Qimjou/VzbozaYXkAhTjCFo7dWAqKQnZNxNMVv0Z7yn6Ole4Hk7
qZlej87EdZg3uJ6yAItCzs5AY1uD0SV4FHt1NW8uK+8gG2V2ane1Dj/z73oDPIPj
NrYQa2ludh5FOQzlMY6hSMn/NivNMpVl3F6J5wfDQ4FlF7gI3rZSX3ZN4FiZJURj
pLzPgocv3yLpj+1pmlyVlPj3W5n2qFKUTR+hsX+4lS8giB933+tk4knecKCUjGwP
yE2VE9IqQraf1DALkR+qRySXON800DP+3LQnYDxlDzpuDu9Lw1JEGBKXaC+OlKpw
p1g2iAy0Oy72JlIAh8dF3cIPHRRL62w+X56sg+OartTPM7QC2x80WAfM4wMZ8xQV
5rZUiGUpGw47nfMib07JjxyY/Z4KUQW+8Xbp/43H0bB0XIifGlZ2xkkHnoMYr9/S
MUNNOuyC3mChqllo/4pyN0DrlXzllPS8GMVYjyOVNVYfUbOM+I0UGY4yCsDCoMhU
VThOBMVCg6tcgnvaRwCAuivpzVNT6IUJ9au2abFdbhfsv7N5t7JaDnORzb9DWn72
IkJqYkL01bsd7EpCmklcvJNQM+vxs5wyH4brZfr/LaPPmnOAZdpfm4N3ZFQDGuFs
iGyDwtQCsZTcan/LDJf8Jq+gUKtA2LvKAkh+MdBPnsgPisg7dhk6v2SgTM3285SL
6G8PXuP9Q2SsRgxMe1Crl2nzAUTJRZFL/qQZHWfhAJ6pH9IO+MWW+c8ood9p18Zi
GkpIlsQk0589SR7Qa/PGDX/MzZzxz0VLulweG+GKYSmNc6F4swPbGnJZ3F0prpgL
iTy0OuONVeao93y5sAKN/yfWerCy69tMo3mPpG+ayKbn1ev0050PsoGhxQIohE+G
UqoI45pe4YwS7EZEw4NxSbFDztn7tx3BLWZ6eaJRnNLXfT1Rq05FLgtc5WqFXCCk
RU/4vOwoWVskxl5AoFG5zn1fxvK9S7Mb3vEO5eCtjpecYydLSHUAk2OlBigpx0NL
8yneOHhQ1xMzvcrsMnPguh9Jg9scZ0TsOsaln015e4iiNAMpk3wweNbtqgJ1k0c+
tZSe+WGRKPofv4zM5C8/Nw==
`protect END_PROTECTED

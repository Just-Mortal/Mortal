`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bFDD4Vj67UwVeRsmBN5++8XWBIGYnWPhRtp6A2U01wRizKz6YbcXwcSJWtu0hU2
SmXprDALq2VBgBfiA/Uz9d6gBQyItskZxSvI7TpPi3BqhHl3waGwIC4sJadxsxDc
778+6kA5EJxUsFrA+I2WHuXYPfl/rQcGI8f71PBIjVYd5v7qjsWPrzgf2DfjVkDG
C9NGapoKE0GOIAioSlYF8XZRkslqaU6DEwL8+OJkouOIkZWpaIFQRzJDacgP65C4
RhtF+b9ixkd2dOeBcior/SpLXr5tAM8bbD5owWxRZj91QmHaMZSeHjkj67QYYhtZ
Y9Q6rFnZXkWoVYdgtuVFAdlF/kYr5nMYTgJ47/TEleCG5laBpnIgnwpn0B+EE/yt
mcWW+mLKbz+jA1yUzw6qZN1LfIXRY2dS/Sko8LR6bs8dFb29ztVhPWU6rZXjIP/c
H+JiZo13Vk2aLwEkbUOXESGyneJir+zHCxuuCVe3IDWPgEFxuLEEw3KGJTzkXOSp
8+1IV2gaYr2u3nkWmUm6AaNBeS6tGKr3NNTI/rxy1ELlyh4mppw38ycdxFslbeRa
NahMunPjSO+T1waGzxlZKSfsDCU+OXIr/GCzYXPH+NHbZQT0UOl5UbWGRwwouuwn
ggY4hs782NHIUnxfi/4liQ9v6EulmYpO79ZSlwFooU1IA2TPkMzizN3SwvNyNueW
iIp5x50KvvhibSx/OzVRtxsftA9AvSY0v7eWpC7p/rg0uBxgT6vOwHgRpY8qL4fH
OcY4Hm2AhUvXN79us8e3Cu8KgA0F+T9b9Fw4qWXOIRjb5VPNzdysiK4OEdZCjuqs
CDU5rr5Q3lK3Gy900mPfXJ3CwR11is4h0bbfl9rhPq7PAZWKW7VZ3FQFAo6tu8XM
38A1OTmWpoCj3tL+T5pk3V58jiNSrE5UdMQzgK4Jr6mAXzDWl20Mjg8qOnXq3DOS
uuy62SWmW7uh8Ka7/1cDVUw0+OytlS9c+ajeyL0t7HEVv2nWgAGWtcsuZSh0gHZe
HAA9Ek9qCbuuHy7b3dgATR/OB0vXCH0Tuwdahp1/eEYVt0onyTRSZHPgyvl2w+3G
mA1B+xyqukR1FxKYT+MsPwvPSWlC9Two3BS2xWarS8QBiFgW279yaHHSy629fqU9
BHwn6Gedfa927VhrT/zywpScaZ6a6nL+lIvTkzZr6fhwgELIT9LiL910TVc2cVCx
QzNM5CJAbs9jsX4RhIBBn4DfiFbMZpMZ5Kl9lKM89VMEbXwIJUnBxCs0NqSojlOc
gQQH95YzslznH7fBvB1xkAwLXKnJ43GYJ13iybFcx9GgRCp3+sjyWCp/+89yY7X6
nxinGYoCm2GvUhEo5UF+huj/F+DWCx9OMT6BhCZ4i6UPrECL20Kwlf+bQjrWjunO
StLXL6YUx+ud90CnPrVygnyuUoo6ewg71V6aYIVnEZoM+KAEjH/e3qECv/lw6mUn
tjDiGF/jTqqiZZzbUHmFaY6ZLYVAHi+92IaQuA4j+dH0hAgDRXDyde2/pq4iwMrx
UA9CDtk2FCAP8iek4V3lG0U/shmgNuoldp4htAw09EQ+dWLfoEeh8w8o8Dbm0PHp
hoWG033fZJgi7DsQ8fLtrLWGp/X8Z2iYHLBsUqbrTzZIH2A+dAh86FiNglSg4YA5
xnwyznrN7Qba7BOQ/zgUNJ8pQ3vpCpdyKnNdcf/6HgsSt77Z64x4Sg5TH368oaVW
ruVeTrFEvRq2ibPDYhPspehraAjFb5DWa+fhBcT/yQBEaIK+HTwbTciUTi7LrtOE
uD0jDm9czuP03S2bRDx52rzj64EIW6rCfJUknwInhy+HzZlu/ryWJe9n5d1J1pQz
AZGJtUIeOhN5XwZsnjxuXr6hpquJCfFf1BmH+cnUl5Y3hDOrv27Th0Ep/v6NHJ0J
3BBeeyJBZwB4V5sSnD4YJdZL5DAFKN+uzuDu909b8w2eETvFmHL5A/8xxtO2oaVE
aPTbvql4NtMPAgah0zeLem4Cxo464O+bQzGL3qhvo8o=
`protect END_PROTECTED

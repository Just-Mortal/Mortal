`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qes5T+Y7X5qTieFbiSg5sWhgqerSIqmdql1gpBImFHSdu+SbAAyCnbFz/r2KfuS1
YqjjtXSgqw5XlYzYKPAvFT3R1ars+tExZ5kG0SF4ns73CaT5ajTX4c+gyHCoAdod
voaGTLaNPNwGwEsrNRXEphWQS+EjAId5Y9u9K+jOLMA/7KADJ8QqiD20MDCBZy2L
o8JERUA8Gn/ckRMpyzGdffZy+PbwhzXvn6uitfFSQVrODpp+H0oZuARDIRVfU8e0
oy2U+DaAv2fTf4vx/wspk1hVd+NFfzKdpr1rSM0gdbxYUB01SPQsyv6XuuEksNYu
OFxuqRImeABAvuZUVKCrVI9ldgO2HyBENqewXqQ6JZ+YdBMbaMDQp1OlcxXDIv66
+XhAJXvkL3iwJjOUZn+umgDTchJbU56EDoZ0LyxGCkF9LS/O4y+sCRkyOReD17qk
WowT7RfgbIRjOM/qTBaQMmp03ak0lq5ogchZna3LlSNvP1wiHb8wRk9B/RGtw3lg
3rQ1tJO73AZmnLgyd9WGtKRrGMYYgmwcbUKpyCtUt0yOX9526ixjUZPTlK1DFEjg
8eIisCBzrMTb1LkJinXsC8SUIRMDRexD6KVpC/5idb92/CQwkcMPx2cHPSxP4GIw
HtBunM6H7nuWhCxPoD/Q3/5JIWv+ihM2/P+YwpFVuVFR6tDlNeKgAj5A7M9/o93C
El41ZSFsf7S0ipOfczAvkMECeNR7old0+Dw+A6ZlXLKjCk3ZxPG2BCHTFsOkVkty
ytQdohaKHPNOs+AY4iTBcml1MRtqgzj1S5hw3FyJE8EUmq+cqKg9NvWGuZdiZrkM
qbE+oNVuwsB1gm6m++NYLzVZpi/umda6NfPp/4ZmYc3Vt4DVMlk+bixLVY+pq0bL
/2gAvuD3EqjzUyKNjVYF+Le6qENzLOoR6sPCNMCIe1jL8BZU/remqOwejb261O/r
i9iaDfiVEVU1N2OB3t+s1LlRg9kbyDsqzCY1JVCiF58wNuoDIdB7bRFgqxztOSeB
Qa/ZKzV/nhmkxiym3g7vyx0T60BtMn8TPsUGpaZreBRZ4O9CybHrY41ykYo0DBsa
K4fYONpk+Wy8QCWRr/zVTGbVebyF60SWVxmZo5S+UYwaEFZC4IyIQdH6c00tc7Fz
fVx0kdGczOOUGBPYPwQihrqThNSwhKpz/9iSxJ8CoPdPD5UJm2JmlinbcTnk502f
FgfKPJo+Q3xN5pFHBYT9WSKMiwGI/CpFGM8ktJqfFYFR9QO98gA+bJwI8SLGN4tE
+vnHT8mzX0WgG17h83pgIAI/fpQB57VI5uHPjSdckBTgSEeRzvf01nMCBxxd/bMg
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbN7bA9VEq3cDW/mwK1Y1edWZI/Btvb7e6AJOgj+q1c2zL06nrkdmADJ9dkp3FLP
VvhiaSjC2Lb9RJT/FHRxHchZHqQWicE6ZVV9BLVW7/Eho+ogEXPRKVigS5kNpl4B
Prt5kmdOEkINOSBk/pHkVkYN+MiCXf4nf/jwy1AFvQom/0VbyQ32QQsa30fLSSGj
kPr6Z24uOKX5/MRLDBvjRCp1ezZRqbW31+mzIkKVbxnA+Ybl777fYreLkAR4ep2E
WWJIeSpfwzoBOhTb1rz2mFMdfKstzV+YfqgX01rgCYYQc35X38JT6LqyPNhiE74B
2to7SQs5PHzNNXME/OeObcMjvCTZ7LcTxDNXhEH0xJVNqu6EEI8PNXgBSQ/cmtho
SsnT6dXEzqbI9jti6wwONU/tH1pcxYo4egWuIwt5gB6qD20NeBJfWXJo3jTFQH4F
SXh8F9Vf6zzf1usSjoyzpjXkf8EWYDjiNwXg33tLgRjhzr8bdQE0/NDDHhGbJQo7
E6YkCh/V3ox+vbR9KTpD9wgbnZOytXqQhYpzRN9jTa8JGKSANrjC9C3HVAZeHH6w
eOIGeEaht1P3x8mD+kK71oY1Zi5uo+l45rAZyjD1hft003mm+M4Y41tCZohizFm5
MnuEafrNGCgYKyoSluXNSh26LDuFBJ43yRqaxO5n7I5Qxx1QkzHGBA6+bNQvMHOz
HiZhMpLU3kqUCTUJgR6G4GRDtdDhyVJznUXy3R/44V53YNNw8j9Wjdkd44ehjlaA
CFu6BPzcE1ouYZp+PlNZwKwnXlQ9SAt317C0xor8bjyoRz8/45DRZr6xtAoIN6Nt
N8pnEx09jir6P6WsNIHZbH3gvOFhdMGUj+yDXcKhZ1V1ZK6hohbtZ2/qmQTLawhB
FYHqzP+BgEVYmu4/trx8xZho6x7Y/l6PylCoFcAcsR02BEXEEP3fCg+hVJJiJPX7
OfIcqZJ7+oGEBFqi9TzAHL5ZOmqJkVLuGKZM3TzSy3tqGaQwgqdBZvQO6lMK9rd7
RIjl3bKklL1Kf/QrktRlzaP0dtAGbhq6lDWlWDGJ6S+t3RNWshXpCAiqAOGuIM9L
FHk++VrNQg5KTLsObXDNc1WRH/N/syu5G8MMg19KPBpoDTKmlI3uM+S03h3pWcmL
QbFvpG25oSt5UZPd7m3yqCd8WgCv1CEXGtnPQmeVzqF0iYAxTvv8n0KgdoFi8EML
WITi9Vx5K4GO/PQO4yK991oDEXduTFqrx9aBbS8Kj+CP92LpFmRVmTJp6FlpNDht
3V6WRoGPf4I8VA+lQZii+o5kZELiwO+NyuJuTTXI9twwz5B0pL5Z9hIXbW3aWxmC
x7tzbBVEhMuMLUlYw2d1yfVvTLxYiNMG98H8dqDkokU3scjG4FN84gnyf6c/lA8m
NHsTP5cWWmrLfmSg8RA84Wl1/Ca4Kgfx2GLxCnA8TS53tWacRzgHV2JNiTwc4RuG
AqqRcG7bpdBnrvIu2INx8WWeDoOik2WK95xa+LTLDehCwsQ9y+2mukSkEFHH8wbB
7jV04LHtccFMvVul+RmE7ma97NMc9XnZjemjFKZB5kyQVxL3zJjlwMqiw8ZrLV+M
9MGU5DUCqm7+niTqQ4irubOLQHjF8aJTfr+ifwyP3A/L8OHE/r+TPjL+d97UAYiR
yC6h4SyRQxZ1VQHusLSr3tEJOtT91Bgcrxo3lbfZPAU=
`protect END_PROTECTED

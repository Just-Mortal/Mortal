`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b199T7B6GY7FYnSagrpv0EnUu8zwmCkupkZTFuI+SEWrVifvs0RL29SqsNiwlLnh
/kKK1H5MkY43ysdG01q8opKD8MEcMLVXmLRhZRQmuI1d1mttMWss5YRxjEq6bZXY
QakgQ9SyxZ1cFc5SuBD9wVsVqIoP2loGeTGXT8O5FRmAlHIitzYH993AscNJuo0y
IIVPv8heYgIbVHzk5eM9O8VkvtbkqR2tuk/oCe6E7r4I1oaCRO9q6zSnI3+soUep
iXCHkrMfxTa1E84cG4+UOb3lLfPB/n63M9RmiChZ5ggh25P+YzDUv1dtUF0nfUuH
lbVHE1f+I4B1bUodM1GcsR1vWET/GFji866Cac01G5MjtAM2TdZ7RaNrLwDLe6Xj
qcaiRgevfR8KJVBSEWIA8VnKuIHMALpmuaw0q9gfush9NPgcGTJBb5B3gcuO4Az2
X/LmNuBj184ARr1mGGujkUy4tkzySsPInRU0PRmfbDox9wN1Yw+bGuSERhAUXi/3
327/d7gMUOoap0vRwdeTsRCcvf8b51iCsvaApoonhZnI6P+iPH7Gz1OzhOUplVnc
5yduXWSOJkc7/RBVn2dZ1YaMskEE10XXA9nBnFthAY2Ws0HJgXkFUTXn2W5OLLls
859jf0mO2WBu+gqYZ33G9hcG1FR0OywQj8kJI6r07qG0eebQdY0NyZrmYG5NxEHZ
6ynBGWJJDfCsuGfZR+QzDuF9Br0gbQKlnk5ysWPwSDmc7CYpzGErF/WkHw2A5bGw
GItTKRSneI9DJy/grBPvtnpKgDhvcj9Mo+YNgt+nXHbCFyyWM9h0P0UUhB1SZl3N
WA25VafaoeCs9nAwcl+mgVrxq6cBJBxbyt7YcJZ/rPdmaR7PVcvQ6d72WQJ3K8gm
tna6fI80XW77YFtD/hRXAhl6oImvxZQ+FZLqhBirDfL+8jCsjMm7VU/NSC4wsBsv
kiGijEXGKt6l8r+LL0xR7JLRX3eWd2YfXbP1c7zTFvEjgHAILJkYvIGQg3RS9IJt
jiluk+tso0AxKHt7dGT/AoTtNqrEI0leasFK11wFoMnClNAJTRMTv8OXMXhal7PT
fL7AX8qYemCiR/HyAFUTrD4/zAcK43B6dHaEnJ2x+H2Ytjp8PgMHwW9EVnUa2jSG
wYxIXdXUsbG5dqY/iQ+dudJxFp3ZKd5IimVJBlyelS8vhlvT2npIx7EKzED9802n
vfd87u0gslf5lPKQFf+n2m9wwlfjwXO3vlgo42Ho4CeCtsinhAJosR7Ydu1HghQ+
k/R0b/WniZFLhrI/ZgjJmTiCUJL6zdQdGMCgamil1isPvNkLZLPv3eFJACb1icoC
/QY4C4WQvXVMHFlmFQpf8/+SEiR8hb4RyhYbVhhWFgbbOA73SAv3QnGfUEJDq8Vz
5pPm+e3acZkKDcwWYgg/+P/1nvoXF7ySosRHTB0kPQkMZYt3mmnIO+oLsFavnZfi
AWMPb1v36iduQI6Xp2ajRyqSUiAceKrpFJAJvtBfWOV8m+HucZaT5R6McxOKHZkX
LOnBQiMwCkuGOrLtsIOlANk9yRketqLzAZ0U/eBmaEDny4EsUND/O3Z92dLeUU0g
bi2958+BL0R9Zz5UIhRuXxbJzOuXLEeGkP1QTPQtchpLamalxYX6va8x37zYFBam
A8PwE/kIsVboXAC4ICS0t524vnbujjnnzVjgYmpYhoq5KK/DG/lF65H4dcAVlfCN
gE3pN6pRBAKW1lnl/mMURgwidd5a7NnDxGc1jAurAEgiPPzI4zRE8iGEUUvAt4s3
78VbKLjNJbsxG/YgmMSlqKx/Hnj4mpCKPYgRIM4ffc6HYPfcKAUs7WOBaFYajtaK
spcfV0fLr/Vn/vL6aaih68AZhvy5gWvDluE+cuRBWQ3vccOr+Dd5hUoHVbCX4Ccu
wP4HRb/GZfQ6ZSq+HExQHUkZEHfDkAe2SyOCScQos0Rq5Aj5ZzsBAYHHXPess4oQ
UFPXTLxPh7e+CEfXXxtyel+1Osjv+YdETpz2LW5+kAyCXg18tEFIk8BkvP7vo0nG
5I3kkQMJ55l8t1NiF6Rsv9zGKCdJJPaWC8vFxPAJAxEPst022XGFcBJ4tj3ixudn
bCq5hNjU0znHSVjQXGaqLGi58sVU17pMHTP7QMv8X78=
`protect END_PROTECTED

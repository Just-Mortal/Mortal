`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iTN+SFjPw6dbBNXysoIAIHVPQhRbCF2Y+R981A2H5cKujrVRMk+qgVWWbQj6pR/B
B1YvgU+ZVrHNovsjDuxMb/jIwSvHcwfMWYcxjjSr6tzox2JMyKKYIlKI68hOe9mO
eiHvTW1q+XPxZvSeGc9NshidEPfkqo8vkTHXYhswaqS+8FvhZLaWVVqHF5n7ramd
9ZszBpZMKXqTxhDOBx87LkALjzMjbf3jslJjnsaJjtuGqsS9GXg603wJAlmg+MH8
daVKRFcYHWrB76VUJszNtZBFxyVy0JgHprPKsDoQvkRW0ccVyIkrC7UPoEtlg5DY
lNrAIkdCmybNTkmppkiP9vvxxLbJuy3TXsH4S/toViX3SgEXEWGCUiIxt0d173In
aiuNu3F+aME8iSFxk5twA20jsbII8B4SGnNBP7akPgurCuBYkHWJjN6Y0yoonZDB
78AwRG4hcU0oO/7Z2+tGK9QT+no58TQeiP9VlGUOyZNe91qp8p/VoTo6Z7ExLoAW
ecXi8ZTbn+rplOAyjPbVV6uLbrC8WWdpKwhO/glA7N9v/shYaxUQh2R8C9w0zZmj
u0/bOcCb88/SpTaeoj05eP4qIs89ALpFHghBHLBFe/E8aGGLFjo1R6Dp4z05opXR
ctm9G6qI4uuaGKRdFuEFyNCxC3WYiGrlUjd9lCTKrgH6uk+mnOvRNDNJpQk+WGaY
lAmmdRtOiN+FnL7jWhTo499pQkaxm71LP3WITOxsyYc4GdnmobM9gqSjeDMgrA2a
MkUN9QdntSY0SLEX9JtcUSciUunUM5ZerX8R6wyB39EymFrzK7g7dSLajM5fkmML
jBUuCYGqJTlQg28e2A1W7dTJnjpZt9wO1bohdQu78vjBOLUrP3SYixmE1y3D4Exd
us4FS4hoti/aW6FMEyFIVw5HZFhdJzD8cET1FfjeMzpnRlvuAI6Iw/dkbiy0BkbU
9meKblnp2V5Rz8NcsPoZ9eonpnpUQo9whBdv8+rJkbpFmzBTdR4EiqYl7TgfUJ+e
5rsPrwqfn/ZGV0sNd89PHQVJbIuJslcENhNZM5oWYi7RoHh67TuaH5ihkg89opVW
rqNY6njAWNGk3VTBmDfZesxc63xK4ziRrvQ0mCfsB6aqdgxlAYiLcTKYNteDfRJ4
EXPmiA/rrssxHlEg0ezg7RuDxClJbYxISyGQl6nGUSQCxq0q46/23O9PxPlt0u3X
pLQjhuFnWpMMQMbFzJzVr3Qw6Oll/FANnnsiStomwSQ=
`protect END_PROTECTED

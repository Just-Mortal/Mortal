`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCDCHUa5ywpV+dPzw4nVmAFC3JPMA/aTXpZAMgcXdEQamCBpnbhohHY6pLZOcyt5
ZxLAceBCQ78nebSXFhAslRJLrALIV9Q0DOCKg8Y91l+inNaa2/0WBkEPCEeVnoJ7
C8Ez8skmND2LsJD8HNbAkQj5JvNazQ887Rqin133SVpSi1zSd4JuWTIHbq0FH6bm
hencz913lkLf1Vgczc64XvuxBLvCqLw3UzxoamAQK2vDe3vsU8PKFTypxLdix4Ol
gVmIGUwFWUIx3Qa+k/cbLftgSgPuMheS1KQH7HKWHeW/+ETl71qJj3cuLRYivz70
bjOdGRjrnBL3nAlJdX3MrYuS7p2ahit/GfI7Y3l0e7zVLmftgS2vt20PK4eTrfH/
7kO6BJ0o7061HW3Gw5o9o0fqJhBNC8gmpSiir0p8QvlZ0hZtfSw2RHD5nSgygpRF
4Y0w8GPvS0dvpwILFwDQtskAkvh/0n1+MLeiIB8U3xFMJ78bSanHxi0lmWtSPuBf
tiijASH2ZXOnslaEe6c9+4dpvwv5lBegqnA5CtGM7IhJXdiOM+SI1KdhKWQ0eC7z
nd+lmEDF2rZp1FSfPJScGI3fQGfsLT/qMSpeccoKhFSO6e1wUTY5JRidttKK/K4u
WeKMp3jIduRVyT9mf2jk9tXnA9js7sTOCF/AogQuoiRwp5hbJY+LfyKM8YbHOULL
kxzfy/JypKYg8kNvfSGwM8jGFwKaNsv8zV6jPTfKKliQKoMZXUJzY93+0ts3jj/H
sphvwMuYf86Dxgjsg0Z946G8wx1sMyDJmHIaFOGxDO1yfNgCoyJye4hw2JyECiu3
x8YOaOi7sH+qmdcYbNbvZOmCZVHsmJwRNPNmgn0bHaynhinQo1vSWLSjcUv0v6Wn
tSGezX9BjWLoIir6FYz/ayxGI7get1Q3sJI3vOQ9G6EFx4f6Wosu2WZ5sD6KZC6W
ZNiwi1w+M8AeFpOMbOhm7cEIOQUq5ifulI4JpafiBSlxd1N1eUSFLl1OaI8IZtZg
GCRMY+/3GfMv4cMRYWoo1dOyF4Kt0eaYQEMdsK4Y//h/oNBHc5eYZsHoWJR4ONdu
oo5/ePyktGxAmaDylVB2TZEgU2fqQUQRj9rI0TwFvw8VrA/Pv3nyRTIJnvV+1TJV
5Ai+eSRdzF49IpHQnaWglZx7FyRuHerFfek84ubyGpC+Rb/gVKwwXe8nnf+EeoGR
MYa/3gr/PB1OxSBZXlEkP4vkmGx1mhrQr+2tarB6cA00sdrypkhy9Rz9qAhnSOk1
skpcx/6RaMatqt7jsDmAPN20tcbcZd9Sgqmr2fjr0KwD9wkmx92LXZ8vjyx975my
9ROAyH4k+Dt5bwWoT3PPpivl+yAP7licpVjCJZROdFLQ1XDOcPOzxmrvyCGzRKr+
rHSub8JH9216j3e5r8IkcqjXTdR+uPqk5zSSLzmm5/k6yUONmvrZDAzCnpmzKmqh
0JHM8Rc9bCBejnbVUhKO80sNU5fyPeCL4Hf/M+Jrw9VXReXyatwY9y2K/ctrvrKG
BqBJaeYWRcnDMKKR/Hz5wFAJVgqU1BGhmE4gGWWYgEYitciLoa8lv5fpGwdFTapw
mEF85HKseRNaE5qXHylIqgys4Kz/n6ap/h73oISXBr4Okmr0f2TMaaocvB8rDUUe
tfzQ9CKDykhaiRTwy+bohCEYeow052xDIGEgYMrEXt3XnE9SBSqwf2K5aHAZg7gb
LjHjYVTiH6AX5/KcCMJ7RKQTQz3c0IFQMr28d/HuaBQ1zNVHXx99tA9ptzH53TOc
Vhw7Ml7XhuvglJclms1N4IoDyo9Re8JFmXScZ6xs5EtODkbtzv2meYB56chASih2
rA3pkbJWUQJBrd2iRrkRnAnaP5ZCUUXYi1vmepqw5HaumXcFUC5081y+p9K5M4G6
F7fBqQbBEVW1oCd7YkG1xWNtpxi7QrtDkspOxeP/XQ7iwxo7dqAbC3zqUujfqAsA
H8ChTiPjV2fgdgUji9ObiQdQVrOm3x+lBQ4be8pHBx6ahxKjkmU4vm9Go4sMLFGC
kaFd9xHSFzzvBHNg0eM9EG/Nxp0k9TLsCE73LESxEfQWZUfwxWU70Pd/AfYHzC1+
XU+4lWVMKAgXojkrV7Vy59mWBblUmzHYsAfF36KUQjk8tPaEcPyYtCpOzeIY0EEf
Tb3LWRmt+iuHjK3+7bkG54VkRfdjYncXRqeZsixGyr3sy2zh38Ni6ysSrN1ZzN46
EBq+S9X7emIR4rOAoR/lFvfN46bTpCJcCFWS/ak3sPlkvaYwBokDtyjP86MkV2uS
pw6ZWOvJfrztC36kjIfXGcglWwDSHp1iLzU3UzWy2Q40U2RzBObNMRZba0CxduSj
KCuv0FP/h6+ozIvwmgagk2wOgdTdY69vEPFCd6UfTOFNRBOwsHKpcsPdIGfNqHiD
5/Mc+YMlkJlTCP7yl3dBKLkC26BiMHjn52+L8+bdveaBKUAjCl8xPjwTK2/aapSC
g5yQsBLH341FZTCZsprZFNoPicGoUgUYzVedSrjMICXN9hvpRbKXFDB4dCRnYrt5
JQnAo/JsJ2nzQPOQxNfCWuu2vaTfnbmHKiOd46vGfFywyFQ8XVpU/wmF0BRKekaP
c+Y2RRAQ7LxLFPEP9oMdgGm6xZv8j/HrZaYrQORj/hDNmdYMFlRl5U9syTGjIMXM
ropZ4TR/rhRsJ1WFv3SzWa0r8+9/UYhFHAF1T6S4tdd8XGvOrsljl+coZJYVDfl7
tq1ZaVDQfyqeBSNWNE90gVRjuPjzezAWhgmCmJ9G6JB+UPoq+FQ/o1M7/bMUZ3Ta
QCATVI3So8xa+ZLbQRTFHcQSZpHrmrfn83rALUNtpT4tdGLupd/3FdgGQsyoLQox
QAALEq8bmqPtyTDl3HaIERpjzutRDFPvOqbFL1/P6ErkH2xZLPSoeCmrtnmToDdw
QB6iPv7Ds9bqU+O+zVRu0PYQiHG7cMkV2UOAYN+aQdGVu+VfjkOOtDYAB9TMr6Bi
IoBxu7RXxAK3U8bytTZF5W9q6+TQjuDGzOy+DbViHTw7ObWC27JpKL5PKK1BGsnL
xiOILF6WhH/EgXRQm+4sQqpLgBFaHjt8/M91FrVVqnPpc978tUbnChYPbP3QeTen
Q8VFvbArgusXGakATM6Gr3G38Yq3KrA5h5AABbqfjTAo/RwzX6nyprTVr9mz1F7K
LHnNt87oVRSVWjOP2qhCsgco19v6EjVZ/94mqArv3HWojK3UIStLXKO0J7245Ya9
lb0+mqfaeNoGJ+EdrAyKAzEAu3aUzocQqO+twOTUjQhuQCyvBqAbirXZdn4xm199
Psqy3Dc6mmabg+30UvZnCJYUwfumO1Nm8zZpKoI7ptUNqstcKQXFgtkzQl29aSl4
MdgZFgwkvyfOTsg9nAj/avBryR8Hwm6f4qinIeEVC2dmfAYNZ9jUWRn+rQJ6iS+m
m3gi9txbTg5JSOAVyGWDXNfm8DS6LDHjCv9YvjuZVED2/Aq8Nbt0DDCRnRvT2mmu
XQ9AJKAysWB6VJnUigJyQBGjbJtqZKwhzXw6HTDKC25riphq4wCGPaIr4+0eH1bi
uNsoFQL+r5a8U1OGQbvJln7r5P3KCHhEV4GX9s1rf5F/6zelTF5DlPAs5iFnxeZT
4afOPDryXa3gpZkdLHheHcvMnfGcI0YUacRYAHFpojmfnOmIj2BtYrXCxR82AT4s
6XWOTKex4igmZcFdm7Pl+wGBtWpn+414CTrM/Hytd3ba+dqYpR0JIbZwaTsvha5a
fx2W/dEq7meotUZRihpP23Y8QQ7z3dg+E+Xzw2S36NWuDYE+ud95pMb9qknnh4p7
Ze2Q0wW6oG/08oDI8SDAoof1wbAFBxdhmFYpw7364nyhVgCskKkqE7/w3N4Tpveh
iHVcbat6gxFal4uRzZp0ZGzWBpTsu0XNnbN32VDvE/f9DOco+mtb6CI4hVedAju5
P0agLcXWefePPtVq/i94lLO4C/wIp1kuV5sspl2F1qfeiW0unalOfVTr+tWGZmkL
LZ8y3zBPTAec7LfYHL6y4AwgGarJuZol32aVNQiCsIwlY1MlGXRmOHHsYfYu0ZXe
yjIRdH0DQuD3chS46lPwoDJSl/aY91DWY1icmHSvRcMbC2H8OUvGK710DJiLaa+e
jC0Pxhz+WMJj58DSeaGEM3oyvIaJ7YGH+sq1Enk44SmRFVqAXCLb21dzil8CkkTm
F38cJCNLhS8tXXpjrIz6LrC1MFxJ+JyNBeWpzNaUxDhVHkY6TrB8NckcG6x416tD
PU3pC6LOAfgAup2Hr3QDwCy8ijNGSuHO89oSG+NrNCa1nqXVpVW+iAfVwFb7wxC3
BhTN3FYXpGz1jRp1VBAAQ279GuSSdyLTMr8EKNUQy1jitREurPyZ+R1B7MjBARub
tX+NjyBqTQ1pl9t271BPIEOEsnW6QSlLd698JJlqjLcSyew2ZPAm9YrkMzZ4Jxcf
5S2Nhk/l0tavh2/MGC4pk5pzmVKGJgPFhlmax9fS2XnVNodydFQHIxUEjaOQMqwf
ItOEIjZPai0HHvmDl1HLZ1gnB99S+YuIi9JN19M9Cm8mZK7F6Ys8BJt1TixN480k
Bm3RLWrq4QbM+3PPsBAMKycdSC38q84ezpUBhWvh6Pjbqme6qcyzUdP4hBASxzjp
mPBzcClUuGzVf0lxCgOCy4HvBlRUusa+XNCCGYtqU+peDuDbYLEybmoIs0QdWtzd
g4NB1i7MxyDmRgxF8jkX/zu4GIiXI6xhRZa0U3LwXtyQ4ZsAhB9/vBfATiBhLeaV
gqPVbH+qSIm22VqK7IUt3ihayvl9KZec2zhuF2yzwZ7x/T4FNOISwY2tpSMou2UE
rPa6CSZkItoMIlgG/8PyVCG49h7oJ/cDya3djfshm/1G7s8Ng0tD7b1PhakefJ5z
m6ssegcwp/4EzZyj6kI18f73M1D4nzGjGCTvMc8Sx/iZ3Zr2nFNngOpg0bdEkHsY
gQs8t83vYCqE1JFgotItx1PPbXL9HcLxeviFIDyYE5VzjFYUgamp6W2jh9FG/1hS
0Ns1/6vnJzcvogryLan/Wr5/B7lBurAbzoOEaLspj1MbHqPoc5Djc6Z/VhUbpy6W
7EWGb/+ZN68EnkAs8j0RhHmAqutqzhDyVPEM7HvJsCUp5/uB4o+P4LEM75dbpt+F
Lw6+QtibRL3VxLQKrLoSEMj7mzaVdCeoKG6uDHZ1VNStwwCelYTTDdpThY2GxbHl
UmUlLePNxKR/SRLzIWbxO3YYvkhuhGnsCMIMVa+ZsLR/iqctayP8oTJd+jxZ+qe5
EugQ8jG19ESMthcSgtaipqNCcImGQTvQbNvuDM2hUk+uLQ+2XSTIhQJmRRUok3/y
WkJqBeqJSt3YRpvYe77lXr8Gv2Q8xP5MkBmz3zpyOjXDx/CNr8et49eQ+Bju9FYf
4hs7OukRyltZtRug4of0MbAvd7T4oH4eFwiW4gnqL19bdlPjNZQmwF1FUZ7v/1R+
/BV/72OFwDFNf36tksqyRtc3DLDBJYbuWMxHtoTNxdZ0S/uyw2UUt6zJl8rKPJ+F
hFcR9kb2VKOY6MiuQSDAU/hMqRn3SR4pPolyZSi2SLnz8CCUjfLYRaXbaCwWiOcl
zl/Le8GHM7+Lfr+UPQgULMSbB2XegXX2DpQaUEzGmHWcJLHxDnedan81/Gvd410U
VxKHW1AF3or8Pl1RHwwetQ96GcN6wO8kFvkLaFfJPbT5OKE6f8n6fSQAqTc9NzPW
/3yUDinJGROj2zxHq9cQctkQCK+k+v52lvjkQOVg2UHSPf2zv7dW4ag6C9bs2ACy
URQlVwQAuvIDtym+Ry6Jz82OZ6b4yIdDZ43tDLQYzJdQ7r0HCEOgjVy9GA6xANcc
D7JJxP6amUFif7Miwp38v5R9ggvMlEn2N3cxF/+VtWCWaWUNd3Mc+DJO+y7qGhKP
I6KR14+Ab0ibPqax79Yys+TQY9JX3gb8zRDjUg0ttFxDex3qtQIvjkc573oUgXJs
0/k+3GdpfLYCBBRz3g9MUgk5eBTYmKsmBn9w4EB1sTMLIdB+al/2GmaUUamOa7rm
hYhZ1q8iWPovWPdDPSflYu6DsLCUiqTPIOZwXnGxuXc5fU891RDetMllEBidALYj
p9FykAENtThqXIUhVwzMfYjwXuGu9iDR7B/5t6tsGCggdrifwokLXW/KQRblhqXr
Mj2/96mb8yhO/NydJKdfHVWMQEtZeIRBSinu1ynBzWAtOpixn+/VUxKpVOjtVDaS
DSTBHAyxCKSh5c4iIvTdZjHOW1Y05e5e1lvUGTQLYOWXzQ1x4cm3uCLYBUrNooeB
NohkZmTmi1UC6KQ5cw0EgGY1CQio/mfv0MBTO12+HyH/BRarszNITiZ71eoUfZa8
H+gpF5rTcgPS3AagVdlLhyoVrCgbNc0K3BcEWFZj+JDdC75DIt3zYlQlnAz8kTvQ
88NopRQERpV9DpGxhZKM2bxoRSmfESw30yKY2kBAWb4HRBTONa0w7SDX18KbC+Z6
ip0RidpavPjB6othqxpLBF3GAW0yA38oek2XFyGti3KJlp3R6pnbSW6fZEWOL3TD
Ej0+XO+v2lMpOrDwCgzviGpLGXL8o9XXmjqnvxalDe6p0OOB9vrkCNDX45YyaCW9
h0dzun1pzXSP5yOOTzq7vDaecakT+I3L9ZhqlFnsKTgn/61uYadCaLEdOfLX9Ryx
UMaABndUQ9de2edNaODdniSOcbVsVTFf8SKkJeE0m85BsFrAF9yjMVlFpy6pfcOo
dohjmQelyQqxcum0YpM+rIGpZVyo942147H41p1Erisca43kJ+dDG8aNBYfYw1df
CGyGkSHFSERrTsl1+Wyxz0Fyi+cP9zsgNXlN7pQMX/GlfOSO1ZYfVTgRUr+ACpWJ
ZUdBlvBw9QSgFKZA8hVPwBQp4WpnUO7sdDnlMyf+dw9g2uaLSdqFtsBu/3ZKznjf
z3vMyjZ83q6Sn5mXEVDTICIFzPLJE3ikh91avekH6d95rp6IC+s7fv6VmE/EhwV5
QnQpBVwMSpAeNvnyl4LfK7EJPFRCpu5VA1zxwh3JAa3Rlcadv7psnHqqBiTU/CCg
DYHphMH1PaPVzLNgxxQQ7kyYRPBMI+4/9DKfAI1gl9Lnpatm94l1eSDVOJhKGl8v
ytEk1WV8uEcp83wB1H1JQ2SxQLBbJfmab5+EWKinbHxuLKU1inVu1CPDPykmGcXZ
uw6DNzFQI4onNg/wuwC3cXR8js5WEH7JGYdiiIOqJygO3IS3yiw9tU9dMqGztGfj
05YZem0lA3ryt3K8gh7v5wnnz6uSWtS0flYeYkxH6GIR2w/Gd7E+zkqieyCAh5kx
L+hT/wjVekVbfiCoZPOE18cCatDUmOKoIaNTCzEUg9GBjG8tXPNcl4idcXx3JG3c
knUXW8jbmVfAM4wbZBGZyHZP+TLJwDLsCP7g5ZiZHgLVvuWJVjuwySZP/mxg/wGr
DRHfcniBWzODIMa+/hEf438Cl5EQ7SpvJ8gcJCXt3heAA5Whj3O/ifi8WUVmt1PR
5VgTwHfuvp2s9xxY9M8OnZO3v46dteXFXSKnQbamHTBvWr7e0sRl/QO/hn8GRh/G
rfXSj0yFmQFYhwlfWYx4Y0h9MoKTp1dLUVsTU1lUxSFvMQ2JngAm5d/nSEhPbQAx
kevIeTaXaS8F4pdi04M9SIL3ze82faudniNVpzbPmKAH6XLnWFy5nk9lrGZisjxV
uh35jQlz5RP+D+geaKQwEWbugvRl1XiYY7dbeJKSPxwvv4DkatMACIRS7sJSIntv
SisgStfTWQ7w9x7lLTriGH1iz4FBlH23IJSv6SI0nhdm/5yrzVq/6u71RTQ3QXG4
oYjJzNyu4gJRoPtXCO1I9ymKAByQ6DRM+/8LdHaRy7Tuj6MXZdWo7zVfo6Kz8mGn
KJSeAvI0Zw8bx68k2Lu+bLELGoZKftAutQdSXRpoMK23GPulXYM7sBtULdyeaB27
bCz0cjGYjvROSGc+dnP1KX+MgF0qh1zaNHRwfbGm/JYSOPycOkLZlncCYZsdwd8O
jc3W+0mSJA/IcBN/9BXmyALEEZLSE9lqJmnX4byzAxf0HMPOmr0eehufJH1Zi7bt
v4shF0SFhF09iK0E5y/zvTQc7mQarSMybKtbIYB+RDh6q6AdcofeEZllNFrTVUzg
LHTsuJq08A98OGrdodZbzZIkk2BVxxbgYPbdUrZmBBTctyELcjPHHyRU9Z1K7FUR
hRJL9S7DRnH0s4lMDyLpxmfLTVcvhLarxlnd3XRfAS7VaQtrv/OtKmdACJjNPGdD
MaplcCCrFEeq9TOzcAWHHRU5ZmPEhnbZTlaK76DUdMWoosMXCWbutPBeDzNYdo7n
bem+/qxE9+QWnHu6ZxJV3kJ9ElgPFhE5sCIuUlrWiHOnZKfM6vzP9sRyc0ie2zSk
y8aRUaJMrP6E1ORtsxzCFaN+nQ+j+kq0lJLCebzFzPDOOmCumg4ZAzt8Qp4pZ1UN
akGD+RgTNtK3IcAQe7IAecRmeiddVVe6oJJLu560W3SclD8hcpIzL85fQWnNrVpZ
mywqSMVjZAaVXTlcnMKVxX68kQWal3W7XVvOrTnxsOmoZyRgIGNXeRbYAObYpDwT
UegAFgvbZKblkGjq0B97IdVCjkrc+II3sr6Syg7lobVEV4uzoLF9hFVoWd8WVGNS
aPK8MUbD6ngcKHtW6jHHlCAJAgg2+hRvyfGs6r4Zj04aOMlYHdqWG/dGvR8ObcYO
QWjnBuj4eO4KPg1B9MVYZV+6dkC1Hu35PKyoNGYE/G1Z7dL69JA6DXk5fjpkLzt7
7ADLe6vQLD9t+Pf4MbDcBqgi36Y3tHuxSxVZ6q11mOreQ8aOnglNJ0ZmVvltMNZX
Hs20os6EJJ1qahdeoQOFNe6I40lPrcSN92Jes2Bdaf4mwBwQKKU0vlZP4aUu9Oxo
vBaVLId9dPk1GiU9w9MP0v5Qhw1+q22+tZS3jdVaM7ii2FZVfOYD0dX5ccWQBpJ/
FUCrJbswOaFKmJBdrlLfJEXezMJbHTEvy1v+nH6jlhPfwih8cVvc+EKm/jyQTIcM
DzNodRM2hF6ndQjO/Gc/A5kur9Msz/HVxdVgCwnF1qySwGLPLdGmuVhcIJPh5Jy3
EFgKHN0K+/KrGdON8jmNp/sTLFIMsLs6BxNylsxMbyY6jK+asxpAEvkHiK/S1f6L
sTix7WV7r6dbFDkMt6zB1FKbZKsEbhBosn0hj/OU3Tb0LbDSaktt43V3SCpgv5fb
gFFaErKeKsYbJqPHhi8sBNLPrshMBFAhQkm+h1xIWS+cnlqgV/Iq6FQifaHu0oUF
VL363tqv4pplqelcmFGsf5PESKxGV6BaSw/T5sesGi++vwHwS7Quu6HnCgW0hyDG
laD7rj1ty4qBFNSMS8+7f5DXNNMlnPWkkRj30AGCvip9Fzla4T1+KZRyP87LHuJn
AfJLBRkSE5BPod7oSZ5z3bHQ5qwK6ldryqv6XA6nF8TsgKpNBKNAr96ubSnQRzZB
30/SraxwfiqHjrNfcjNLaN1W07XtaMpPqj9+TtGw8auRzqnMleAGtaYPEyLXFURz
Aj0zqSSQI+lupZE5/TpfzBEw9tx3anDtPWXmBfCsKqRryNCu7+wSJNRWCLaw4Vrq
pr6U5Dpnz0L+0d7SQtvmhWGtyh6JfDVvU0MGKk7dy2EZCY1c/GOCbsOlWnrPoZwN
pNkS01p5mIvLmURoimwNVqOugXdrUlZFqLZIHfH27nj07T8gBL47NJhlfWqXJlYP
Mu06CqBtdPoySGyLLIpMz62l+ljNDLR0hcUt7qWNO5OWT+00Z1BGpNfJd2lShbxO
R6N5nC7c4ziS36qVswUumccTaoTMl4QQ8+bcaxcNgrHbpECPZLEayH+rSuDbN9zb
8DlIr9gHNB/YF5ofpiqSa7r+z6UfO0v9CPgJkzl2YpRi2OwurBe+8+cVO8iEzTDK
s3JUdDJgyReHluXi3nZLnqsw8dQpG2qqnkRsifZAR5lo48RhOzskGXczQkHMUQjh
2C0NqSAeIKeC7GHfHC3MY0BGsNyr5JvOpOrBmYu+U6528CUiaqOcggq4xREqLeMx
GlalNpRi7oFFSkyicJAOeWDPVkwJqaVtynDH1Xoj/0/XV4b2r8p2yuQIZP2IpKf9
poU3EaEzjH/LJ+/yW2xWsRMUw2lnZTB42Hs5AFqCdapTZI/TFq3aRqMZSrNkzG8s
BDWrXJTbMiA0ik0a99/LtCU3PcxITCbb0Jtqe4grfx+ycIf7/ogOBbLH2/0rVFX/
mbfBzVC6lfYz5TMsr0Jno1yGEqNF1cqA7g5kzn/qEVwzwwLr6FvLqgfUl21aTJz3
9gJGe/AFcY/uS+6sXHEuYMMnQxjTO7eO5SLRJAXEcPxs34UZ6RdLLTmBpQXc8wnz
mtsshZenkshq2/bRIn9SSEpFHOgh7lCoKKGEi0l1DQ2/P+xkTaMyCcnISgU1bfgi
6XSj6p/j5KbAIEy3djoA57Mz+V9VnN3y2iSern0O31R3IpsMYXAhdTiI/iXsb/al
9wv0MAAPXg/GZM5oecXwp3pvTn12dzDFcZJ/xMpDjehIB1TyGrdXm/eeOlLp/eTJ
hrBV50uSkKXSxJ5WoabjQ1jCHgAfVhF2m9qiJIfbOlkDrXbySApN9YNbhzqQ4HTW
cdxgGWxynQg6Ptr5cjWlACBqCRCbleWVLZxK/6pE30Dwdr8H0ktXMmvRuY/TsK7q
XdbK2VCc8z26V0r/Wlcycbo+SQmYNP7zE8Jnwsv99vQpdIo0o3WfTPybF/T4pbAu
mSyvTOTS7ynM/x1DZjnLB/6auG5ZJLT0XrWsnCryokDKOH0mo9H/tQy0jrTku/hV
XtnBw8dCxA0bkP3yZcGNpxHkeVp1av5WgS2L/ZEuMVlwm3NwaJYKAen7PAS0WrSt
KNaF9ULBmEQ7KVpQoCCRDnxrV+uGnXwSszli8r10X7dmiYM+jvyt5VpXjpB0B3sB
UlCqsUg7UglGORLBdCLoXAugpd/Lk2lKZXuY8yXxf9YvG5+0VnsGrrTWz0PpOrfX
72kXxbknMNmVv3aHom1jScj1AklAIyOxC1udH4pGEgmiHdjNkQm/1A+pB7CrZibK
Rv+oGpf9GomNSZllcYATBxq+HoPk1fxWBTI3+qHRsHoLjYfS8VN2laIoZU8mVSob
qxiFCXAU69uAGfC8GJ6hA6Kaf0f6uadcoXLQUxRMYcbObQlCluV2I7gjt8yw7QhU
1AjyXUFI+pdITPrAa8nPbxLyOSVP7GzsBjEe72XlR51YxmzC4g8XM5EZAQFD/mXw
mi1/ztT1f0mJPszfDhXO7Oxu4qwCxjA1Ql1e/m5IAeXMk2dP7pgghzG4eKCtqhv9
cX0Tk+sTGLeK3LLoz+WrQhRukXAnog3aGC1LsjBDIErDbKs6tWtiWlurajbLcWnq
zewuacovcyWT3zmGgDczx62c0EtFNk5yZnvJ6fI+HD80YQhefgUuYpt7EdA14BwY
Y6Q+IFq70scKxR/Cv9hMAufPy07ZBAoFEcy55522imZ0SCJg1/GDoTWD87qRzMS2
lWzwTg09jKwttbxlkGYSRvPzp3CcfCHJtClRHv3O/4uctvdGiBbabTytyliknkip
Crh2YY+U4GeU+s/kitlNp/C7c0diAMBJ9m3JrDEW/BdQseQQ6RnhHCjfc4x9HoIK
7eAr3/zwh6/C7LQg+kgAd3eVvadeUZCymUTo5zI4bSDBUlGuM5D1HBK/RsSSGSfX
MowbyNG4BjnnuEspVCTq3pIVPxEZEzr+9gm29GYdJ4X5+GcSTa2EFiI885Qivom1
ImQDaI3VSWGTAOb3zH9xh2IOkHKOAv/7+Az8YJezT4cP+iFpFyaW4uclg2PboE+5
RRKNR6Iua8tG3GlFCK2UVStTwh9gJIQR5U8dKZaxwODTcBW5xxcmwn9J2zcB8Rip
D4jixb03oY+GOa2OGjdIUWjSHAX25yVyRMGQqmvn7zXEY/bWW7TOOFETEF9eo+nm
TWa40421SLYzy6Wj1shT9gLakwoq+aVwnhs6NzOB265OTD3RO0A7I2AAGl86elnR
01PmohyOlOVK61ILUeaQKs2mv30fzIRGkiLs8nADWibpzejzOC44jkgXXIKy5unR
Qm2V8GeCRPB59CCwQBtQIm61RCy5EX56CeJIrzGrSvDAJoByxkSNlhjN2WBcqUG4
d1gKhV8LpQD4DIoMNZqfwboiukMC71MHgT9DwKseL4tVU1ihYRc7azpD6Pj/Pd92
lqs05S5IM7VWxkmiO2ClKRhEB8orjyo+R6SwwKrDcQheKQJAymw0k/Lu+S8s9cfn
JUgaWBLLU7leiLJxrvXhenFEtfOL7/kHyqxPbGf9xGCmI4xA2ggbP2U1yodDCduR
3rQ9HuXa8UeT2yt0z7twKwltidfG2J2bj9+Ou2ooQ0S2nw+cQKmYQ1lMIKrU+/jY
gXFcTZg6EJ6f/CSl0aFVQQ1dITWBOOLIiyunUe0AlD2J7/kL8nQon69M9ZBdGiyx
tIRx8+GOzzDy9DpjSNWqO+PQBIKqXZHITrnH0isqd1HQ0N57YxpjoLEx0RN+vcJO
9fPvJ0d77mr8XC8bRJOSHoEW+hVZsDdIndfRnH5/qegBrCQMndGiFIGKlc5234Oa
9gRg2Xsnyar3F3m+F26NmpJvSaOzHvjlfwe214WzCpqS2fO3l4gLONf/FLMNtMWb
0WPdAjy66XBECvmHhuC45+XPb68TC5gv4tAuPO3eQtmCLvsdfZgI8KN2LuCEslsO
YbyJGU4WgKnTqITE8WTciDQvZIaZtejsXNbEXNKNSslYok9IpTVk8dH2wg0GRbgW
HddWAxJyMG4nhwNGxR72elfAn4pL5bk7KLcBuVEMsqlOEw75OGq5iliqsqPvZsev
abZnENWoAP4RkH5BZNXy0+OCV7lF649uewPyXc99wuqbOAaCB0g6hrqyMxSAu8wm
S2BJoXvLAnX7VSZQ8II89kX6wi1H6HlkPVMcPAP2pN51OYye3m+tIGncQC8v+IbV
6LWul7XYfUPq6wRAcK/6HcYSXn/W9NlBXuy9iKlA5hS52R4e6xP+/4JHGvvn7e4U
6NCcj/a7nvfB6Rf0eXa34fvDxgUAYz00t6Id0ILW6ZSvM/sGlOTVNY3yRuviTNo0
/K1MrHYHsX0uhUJvn0A5t14Zptqu+Yek47W68kJT/ZY=
`protect END_PROTECTED

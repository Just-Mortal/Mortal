`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8Z7VyQaIfQgMPdjRzxfNGGK2lM8eAaF70FGIZDJzkdVp0tKwpsVXsbqPeq/GdBe
GqvHPMBwpb8DHbt9W1lo7irQWsv+jkaqWSJBu9il+auJYUHQFNgnE/Xs+D+/SQ85
5LAvNNiVGSSSxV2ypoU6VaCEe8qDv5PpQExKut2wybFUh85xX3VtOVHCOTJ9nCB5
L96jiv+aAa1nXR5SEVYx/mYdGsXkwV4RfJh1geKzM8GMgtRmfqu53TPBakApGwg/
710YabjKyUr2UzqfQQyCeprguUhv2bH118hcyVG+7l+iSdvZcpcFf96+158+aB20
K7ARB1WrH+wjXQ/AsH1IoGNKomZBPPtjDWVgNWPkomcLRk9JUBkNzxvVXLN86e/z
Bg+0bLlJoHCb7NYdTsfHNlUMYBwCj//HfmSk99lt3G0G4GobfnpMvJqBcfor1q8w
uKTMfDZXsrURUxIQoRgZfDQN8M7nLvlPcg91FeLWbn6hdX0RUFepGE9uMAlUqfZj
0/VIfv+Gby29Lb+ENdCxxhMOTPYXY3umTDPEMZYMyjc5gXRHewz22O8vaPCG6F1E
rdXM0qIG4GtA8Rxge3UNuLO4tgd7OK+ncJiIjBVA5boAHASmmbEjNzIWqdltVh14
XKJ8SPNb66MkCaEPxgiB9xoVnZEYf7qIeJElxhRxylUfg5Z5eN39DKaFqdMrh5dn
gl8YRPXHlqcpIIJDCnr2drYdFI2W1jN9bJv4Zqp/ckHUbvdIwsHzWZui3ASLXcHt
4o0N07PMtw+t0mlw9BEWUuHPX55MVzwLmAMEw5fxx0qIw3QBVXqZRSMq/xUJsmbc
0aD1JQmUjNjf6S26y8cLftEMrN6C8DeUlgQKR4E+WTvljrg6KEQOy+pJSoY1NvWk
AYyGUaGS2mCYihZQsj9fVroSFqx5ujURq4qpK+WEpWlBUh5gfCo97TTFlNLue/uN
jHm7qkKmtmIteDRa3iK123OIdWrfMLkXYp8tBh05BCdyonZJ5rjv+4iCANb46w6O
2G6QQAQ6xm3NBwS3ilg8J2Wdb8dRGxx88bMmGPGLCiuyrfz2kTjk7wcVw4ilb5Hi
xxiFAs3ir3RXG6KTFJLeHfiq4o2PoDKrH8xvhc18L0iQzya68WMAw7iH5yuSSaT0
zdxZka65UUyKGiKUMTZMeaJ19Kh623ueQVZW9KYEFSA9tWrKZMo9CeZF9p9fKpeC
rhCi63Fw6ayOodio7CjJ7hEgVBqJH8vnD/ZLqV8eEj3fhW9L+HoKxKnbWJc8jUHA
f6VwWPHHyLnqcnynlOShIiZoQcAZQ0osakOJrmm5bX2wCV5ZtbpMu90usAbgf16d
lnugcLisvGVWlrZ5mtBnWhqWOJuwCRfXVN27SITRZ/dXfFRKx2qo1MejLWrIFvIH
yeRYNHnusxg+NiYD7NEbuwLBjqm1afGJ6VK7B8X5m6VmE3AVSbClHrRoVQ5Sk906
os9MxDNBsNzXkknGaxC/6pBsHUvR/cr8np9HSSpuShunKpoxrR5cPFreIofxrK1h
RCLGNzRPzO3gfDWpw+XQpaAmFVJFDRKjNhFEyh9q3cOQArV9+/AvRCdzehgD7mqs
lhd7V3Ki8w/mt5d9XY23q4Yukae4d+y0jX8GEfbvzKWKjivsdPeQw2HtL0+/VAVy
uemoJgd5J7mx3Kv2Hk/TNbY/Xsbt0ccfqVLnhp8RGPcs+LKYedlrC09sBAjLmBId
r6/Z86jJ8Gde4Q1LQqzC/9Mx93F2Pt2j3WDO5p5SkA68NXgsIQKliWXYOPp+1znh
FnooNX/lVshdd/JGqq1qQjYlzKY/KVRqkj5ksRO0crVybToCPktsunV9ln22AWH2
rQBsg0IAQ9pLW7dcEZUESfi8Lh1Z1MURg49IDw0XKlyH55uWelZ+0GxTnqAipO1D
qHb3fAAAdSH/HAZirjVycDGbP4VSrBm3khIYf0vl/WWrX76GodRDaVvAatAuQchJ
2DidVFEeuS9xDNX9n5uWfWYMCFsxcNd2CGLh6V3n8BnmxYl3fWx5OKjGvD7ICahN
WPrkMgANmgLjheUgK7sGhXlK/3ghdyjXwCbuDyGs8hH9Pd2sI/6nq2ikNsQpdPPB
wui6G2Be5eYRg509fVX80xLB42k6dGTtyGEVEa/vTyl8mJ3wilOYuWQ/F0gA8y13
xcf+mKPXT851w8MKnAM2ZrCTuXKBmZt8zMMfpNCwjum2jouJghL6TI/+UzV2LzZl
HLTOMzzqH0fN0Aswb4y6jyTStSJpOdNHZGBnTbDoVSk=
`protect END_PROTECTED

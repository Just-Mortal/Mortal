`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
75nS+jsYlp9lu44CjVbmZHwG9DWO4YcZDL/NvTXiw0B/zQWyr8aOgJRKoF3QwKFP
/L8SsuQ4xK7JobNiL1sy6x4+66vy7YEMPyKvwIDQj/KaQBJAz45uHtzgndb/q/2w
t0KvNfg++oHJ49B+Pg+Kd38s9HSBb31uyQuG1K+JKj1HYfUZ29H8R7Fe5uobxTai
BOU8sWEtK8yDzk0WIHKCZ+QuLevr2172//D8kKP6BoWFd2FY2zDemr117G01Zbe1
gWuHJiHm9EJyKyELOA925YrmCJ1Lr1CTcd1evGe2hNM+cZLeiJrvmLdXq3d+wcQy
nYJXgylVatQk1VdfthJ9vLKvp9gP9dMX7IbLnAwvsu6/QrVrGkaR8EAOiDK/TQrm
1eoOChTRtXziyunJLOdUBoFWmGjSY2QBbeSFwzpF+Wolcazfwbklpv5Ll+xvBgaV
LZ1FZizJxyFMufx/CEFGuyy7LnP/xHjH/6JjRdW4a8MbDoDuLpjxOkr0LqnDWgIr
DmE5SPeBqmgql2XgoLTBqgeWYxbGiqbaKL+uQleiyxsgvZ6LrU2ZnaBSmlrmVQsA
b0lCZuJzD8JOkkKQ2C4ftBV6m3raFsvaEAxaKFZnBwsmFYCmlXtFRUT0tqPOQauk
NIQqmR9qkCSqP9eEyAF8yATm3CPzFjSmgAf2rgKXBUoYTWvQZLh+RsRtteacl6Q6
r2PseQeaCDAadLRPev1XcjEhCLvuUZhcK9jFvmUXcX9idUEcEK5YJvALdT7P76Al
j1HDee2RquLaujD0L4qeRhOPtN3Ee/0UixRAK7adUFud5uHLZdVTTZI15mtD7H1J
FHIt+UAhfxBcHFuENs+RQ3GWhmxHHH3f3Kz7HBPbsEvG2UidqX5mbeNHV6PJchep
3JLfvn6VegfyZOxlK1cJ54MuZF3ECeiWmoX305uFrO8j3HFyVnEwMoV0OL36S1pK
zg1F7b06BJYUvbxbouimPIyfzYu8oyb+3N/fte/R8cY7aY6YYM55EQI9WoSiMQnp
yz7q4dbfk3YbQZkUr2IwMAv5Xtk9tlhBx8A60zAv7Oq/Vdjw89pRrCI1bvg7stGS
3FQZk6jeOu60zyLlJwBC96tJYG54MjJsAOqAbreLVlmTRwevJUCZpWt5cspeMqh1
xRfAtgnM485ww5URluJDcj10Rm04T9aldaWm2on/SxJaANCQeSTcwJQrD7vf93lX
+2U8cCrScU/L8kW0uruzw5KoHa+T5pzLnmvFOUqsk07Wmu8KNTfnm4XYQ0+qUqj+
0Zl7nQtsmC1LDB0CSrFbUWdiZ1i964oGrXtQj4NIy8pzTazMEDmgGoxgb0/uH+Dh
bFB/DtnBDlz/75hhRFRqKaKrGKgOxdwjhEVAJggBbuKVKye2kNhO9OZBNMZNJ9S/
o9fgFtGUN1RwiRn+GkjkRv5ObOemWXduCOHlmtky6J2kammZEN2Zo+gP+aKqI0gf
CH1wpofsY4yTtWLKnbuPR6egFy9Hd54iqHuGWm/VsWH90d7WcQUFdZzIoT/JbTFY
b5js12uvqLY68CMMumc72lZGPlmK4v50BJSEoKhgS4xTA6AAei2g6fjNiGv3nIAV
6CHr8CQhLrkuzDzqKAAXyuJQhrICOwINj6gDFA7Qoqz/3uiy10mVMaQwTjAwi9hA
5oiaJghKtW4U74s/+c88LPD+WDwC95/XQKta7fsAW2MmfsCJ4qL3rlzy9StqgfxF
KUxDInpwMl3zcMbn+ZmizNkgbaJ18OT3LZm67rROsPeIxnz0D/CJtJlgCZ5HJfdi
kLWtPk4E3mmRBF81oEJUU+ZfcCIkqbYXYHkVZETtsOiusC4oyZ1l3vg1lx5xUPt4
oLyhxcQB1E76EoHgwr9eYN+ff2cY9BHQBxwRai0BK+FK/ifXusBN73QDTcIOt6Tn
B3HTBCW64k+9YUVgCY7QUDukbyoerpORtli8jN35HufkKGpcgiC3nuELb4QKDd9R
uYEltj6ff5u7q7+MgvW9ck06BmD5IVCbE4sb8AE3lnHPXzH2qfxPNVT/3xfWbkUQ
trs7djtnLkeKYaYTgRWYOQmzdwgy7QaAW6uCzWChA+uY3fGyQ9Rji73wLV2TQKz3
IZE/1/pvPo/ZY7mJNs0jbzSHsnqdkV6lkzdZ4R6D0xs8FvofFKjW8HOjq0AWdIAL
1pgNS4ksztvAPaphd+GMoq0zCDmsELyKGVBfU3axuXHWmr8NEYlEHI9PW0PhBnoP
2aO38SaECW0JblGHsuo7KWVMHTBWhKmx2rte+AShgBljWpHldabTVDcDN/ljEYxq
fFNuXmiX6lgZRU2XwtUVhFvSKf6StsuTjABI8dZk0phlt877T/3Cxn9oUv7EN2Ki
/s4a1rhqJy1+w2I+KzLepa4Q/2Bg+mABr4kruQIomsno+bZ3xvqLbOHO2yeujxms
AFG/KtRPw8xgRGs0zN8tNaROysRvHt4woAmcRRfA98I/u3Gzv4f0nbH71Mg5yY6I
TdUQFj1U8gxTHIzCT9d4XrhXzNSJnyD3Sj2/pg+Jyi1/aAUgU+GeauG9Skyn6gWd
ELQHs0xavHBAqBYw9RI6gCaxxF5qL/d+xs6pDMMWlfZvwbJYIvA9/ibLV4Xy3iNd
5nrJYagvb+fjJORIYTOhpGRERkCnI5EnEB2OxkWTjKYzaO8/sZhqlx+/TY2ix93T
sgEvjBMoktKTShjdLQkomkjwN8weWcQEopkKkYpNsIT2DYjnovOSt9LZVyrL+kUl
ekD6WCf1bg+POAoI4D9L58Ba9PQmunA+F6UdQEfsrERFomMaZntK6ZeETeAUTkKk
12aIZf+FguYrmA7pMs+Xhs3Km4IgyZQLW/NpoQO1DL9oOQpLjqN1GE9kOzFUe5rr
g9XgZRIJ1SshhL6N/8FAUWEj8lTX5mbjfi//fpT9RWS4AbNDdyFhkYfTfHUjw3ji
eXa0xm+H0aIXd2K156kK0BI60RmmmiEvG6yCCpGdt+ds8IrgBzP6xzUk7KxFXak9
ZrIWRbjIlF7w5ciD66UJ9t7REB42AflEjzy0BmKJmUZnjJjcvmry+LO8GgtaeViO
Tnz42jlrj627PPe/NYw0SJb9XBwPKQPvABsuM5462WNFCW/MVtd1EvrEP9J57UCY
ZYArjkzsVI3TUH7c95rE3Ct0v9pkqc9LRzHBq3Puo8mfhNX17a6fhJMTxaaWvN07
ruWJhiPEzJebZ9atlUWugmnCDAYrI5NigjLmNCDZQrdr2OU+I4Pry/AA+cfs1U3T
BjqJFq0/+gozZj3btQQdNqVqwA4HIiySc4LBRnFpVMsWdcVUffKGLm+Yqiql7M3y
HMQYHkz3YGVrN6HBRz3NOCHE/fJnVwJLM9DXb9uuGPRzR3vWOfAqg7r7HFcGOIE5
bAvScXyHaFO5Fs3/EDW7MkZODfnX8jBh82LN8OfvPnsgWyQ/9CwX/8vWoZUITzWJ
n+ShyynqychBPMwpTd51H/6l2j65xOn9AcHT0UwDgpk+uDAyhxzSHUEcoLEqn5hR
n3TpKjEdqP8jKTKVt1AApomraDLrDwZtl8v9ewdlwvA+BIs5hUrFufj5F0UMB7Qs
qOQ+AEPNOocFxOxFW0GHH22HxvyzRc8KLBfkRGz1t+mzRm8oI/Iftz7R7/wyutQD
mk+QYrd9z1twiIQA2qU04wprM2CePY6qOJS3YSMK6d2fO1et89W7xY5T0y64Wskc
d+UM7aBVQbQDdzsPyeC4ls/n/i+d2UhAR7bK6Wo5rzXBvtlHRYDNk4WhiBc1brN2
ytSWdBdQOAjJstQKEEcljHrlt5GvMiZCB40RhzydiQWcW4Xg1RGQa9qRX2F9xJN+
1zQfbpdw4Fjfqyc6VCEERy5fZ/dpxbCS0WhzooTdGRzCZs7ioWy8/GYKEuQGRUAB
4KdwQ59ZXzPskB6rYEK2P5A4qTek3Wlbwti3mha3GljTYZZubMV9ulzKgRyVY22q
HeGtMlAPHp3oQ7Q9CF6McUaphDXgjAu3MY7QcCUVDLZCyMl+k5Hb5Mlsh5G21WZj
my32IQuNhf2FHfVkkTd6fRk643rrc0rKaEGg5jYItZe7QU/l0D0+XkV4kEnaZs+8
XOpUJTlSVqRGjqJyNzVveeR2fqHa9vXSYi+8ga/QdQvf0PZeibXGVNPCW/bTlVpd
WDh/09zdxhwPtq/Ho7vSZV2c9bAuHdMAcVDvQPTbxu9OuFT827EYSaeanbhztHhz
ui1iRW1pPuTSBY52MTXgTlHm1bE57kPE+fk5h9eoefNdodQhDhKbCBLVTCI4ggK7
rLmy7Y7hejp/rsEdQDWE0HVZa8ZV1DGB3B9yHK/TxaOrOYX/xS4gdtfJI+uIKKqe
UjnP8U+ZvtuCVWqs6aiq8b+YYwBrkkC/IjNp1tWpJ3tUR0SYxUtbYbCfTzFDbDYb
tgd00Dyt1pk/qLdHpVbGAAC4DB40LuCmJW8togedawC8UtG72o1fwMS6W9au+pjy
9262pEY5VMGx5lWEaYWkqZXIGW76ZLKxnZH1AEPZdwp6Ah0aubHWcXt+HlzS9+L6
HL5akxyJC50eGFSzNRamnWHOK3yVQVQIhUbfDF4k9HazDOb0bUHhjNN/d2SyQp1w
7R9Zh9N1maUn4OB7Toqb8NmvHjt8X+9f+at+oERiVLkrzrMwqav91rvPxkXAQ4CN
0XmBXYctTVcOi7dHBEfk1HxXbkuxHyRHYk/uN8n+NbGcPwhUIjLEa1IZrZuwgtZ3
ePUWLBqTta63Gg2BQY0GBdKfnD/t2LTeU+XU25v8hQxODn2yR8z1IE3fQvjDmob7
GW33Yw6T5ZmT1M7Rld9daiJFkimzCYH11sZ10/q0ZBD569wtd8Zw3w2QDySRcvpy
IY70Nvlmhh7j5XshKgjJGGGarnkEn/kwgv1ZjFcL0O0DWagyQRzdDdTHiz4258BS
FthG31+OpFSV1hqzU6RGbizBUNAU4mf9NiOwnussjxSmiwjMQx3893msnUMLMwdY
tXqErItitPBQtSKXbD0Ch5ptlIG7xX+OHZd7HPR0fL8d0ElpmjHRPlmUMSJy9v4i
oM8Ra1xvJLMXdybhYUHKeiewUP5WAOAbMo0QwpQ6yU0k2St1uK+E2xZvmmCWDiU0
bMvyczUBVeG6EWlhSmlpKdHkEG69Kt21iP/vMR9Arh29xzObLu1u3yXgqGxtcnQK
LKUSiIUDGLTcSJpIxiHmFHSbNv5ZB3EaVoPgFzVydrOW8oc3ZTYrbCDMiYNKUCBc
4ML7OqAUbltly3G8Es4I3dxU4RujuEsvUg+qq538Mi52XK/T7yCqNsldCPdDre/A
RgZOxn+a4mzggM0UdtOrw7huB46W/ecL6fpwTENnguBQ2zf4cNEPWkP4D6kAxGpa
C4fJ/dkP62Lzm1ENJz/Mbn+Pui7Aja8eN6+p72A8DoqdLl4N/hoCLKaQkqku2kFw
ynzwDE1zKogzUEYUa1BT6LPhL4p/0txL2OfqlcRPdrJFSLdyWBahmbslSegwPINu
RZQKXPVnh1pP73bQq1Sjdr+EkIotbOXcHWVqzpeW9S9BvQLH6lSO4GATRhCXwjpm
V4lOvINm4A50G2bI9GV4EeG+6lL7k7fwP4T/2bxsvNR5awHsn/RVsMccrfTxB6Ij
vjp4qzYGZJgcsz30yqWxHzB0SOXdXfkD4ZZbca4WsI6Z3NWAbMpcVHtquGlDcqPL
ZIyH/1VPn1ejSLKH1idXtanNX+4tkGlNQ9Q77/M+vWtJYzgaOWntyMwx/sQp9t0P
cVqCqqFtMfRyIAkPpWE7gavZ7uFqcgW59Oq49Rt9HDyJuZ9UgF6pRGxrpvKIIRR3
weztUtbo/iMRYd+c7uKgZPV54oqkt79ceJCihknhFyM1mjkZ0jxiCC5Xe7PYWPnp
id4LCpb8jBoNTYHZomKSKQEArjYJOluTp3p6db14H4S6BnzyWJLFzeQoEKAScDO9
8Zj0DYqLJYCZP6dOk+LI2F0NsWHABrZkXGcUHmF0JvKr0PlDJ4+RyopObGp+bQQZ
zUE+JgyX7/ENx/2tTdrzFc42dE7e6hOhYEn7XtVnqn7S5oKxQeMsIW6Y0EGEyTCB
n26uq37ozSshuE+L8g2MQy4gXA62TMf1JxNU3aAgk2aMUqGzjbnctbK8O+cYPv7f
HsnXHqX4mnRknWjqttbugNuEgv2Pm3DGKkBHxbiLqV4ZNDlr6b5TkDvxyeMOfnUT
X3f2joXskZGir4fwPB+BA4sjwTl0VoH7MlH/q9YnfLdwjJBVQeJjQdjhFTM9tPMm
Xu1peWy8bK0DB1PRRHqeruScWpv5swukS6jpD5LMzSs7txeMBWs6acBt85OUSpc4
FuX9IzsxGOVtEqfunrdJ5yvqXGYYTwNiU+yCGlLUf4YlZYL3QbR1ax0CAs+WDs9O
npx6gl83gTFgg2JZo3w7HjdhXGDuN4AR04OhisgfgK6+QgCsjBjeFlZjszP/xgGB
0fg8E4MQak+yJ624p/RtBVARpvZvKP9tr0PWdy/vihiLY3JbEC/mqR651VgrfHBX
UeuDIhPt6MVJp0iFkv4exrCGejM5zE6KmeATRU/utdUvijixCj+DrOq4U+WlXShR
gLOODCPPVqLr1sOuos7E8n7Nxmb+GjtLwcJRHxAJp0eLRQZExsqQuXSkb1Ej7e3c
O0+g7TO1ieybv4JrnzOOjp/9V+DPh8sEdYp2zE1p6SfwRj+B8lGvrf5dXiKyLYbS
rRnfDrbMi4bKYwAz1NtiKGrovzMeu4//Gm0GD5xi0Vk76uHkptlnRKCfhaL4h31A
0L6NQAeVqREHKTS7qiYKr5wiA3ye9IgOt3/MEKU1JcSs0eRn7P2gUX7fJh09X1Hd
MGbMqlzZHt3PeMxO8UgYdNuMHpRKIneOmzEA5V1+zLyP3gnu4AVEv/vcsUME9rqA
dvkSbG1CmNQpm44QuPYWHK/NJ/BmRYVfLrNqCbHJc+PNjPWWQS96u2NR3LR7al83
VDFJ32ODFl9UomgLic9phs43H2xNZVRA5GKkJgX4EDpXq+6YFJaZxQmetZ7ISDBo
e/HwqLkJHuhkJrjo4NginRbtIBOQcABDcOchzsJkbhTls00dkg10BP8qawhZBrWg
/jhbjMrYStJNgbSp0sx1QeUgD1K6bNOCdSEf8Edp/gt6U+1lLPY2O0Ig/Egp+BT3
R1FBIC30ahQediSCTNLmuLPAr9OCUo2R76yEA86fooZGwYr0JSC84Uu0QtXjRNIp
L6GkuTk8V6CgzrOZfmjrTi39nxAtN29KwDuU81a0WkOSwBk0K1+do14WT54g7Zd8
cDTPXvlZgz9/QgW6PO3UL5DqjH0KJhNRY4+UYWq3UrEolDRrDp63SAPaiebdeQr5
3ZTKotka//gQsm5WybxKwU85xX7wc/rwxT9NZPkRbO6j4xhlzk9l6XG5vvxxRSOw
XNd9DD795luZOKghmkd0OgRQQQaE1EqdsmmqWOVksu0zdJjT5orLkSk1l96W3vsM
0tg93aaRASPxxKyWmQWefkskGrwPtEl2yYZ4J5sM/TinptE9O8B4bGwX1ZesYoFj
sYjnGaXTVtRuXHaWxWz9hG764yELTAP9/a1K5zbr05YtAQryuFR72+C96vX7pbt9
Xx75AibRX3GQMmfxFvZSIpAeEusefONaLxxb3UoD7mfLtY/gMqO1B0owaglrWhcB
Qqc4CMIKtKoM5ypBuU7EVsjZdi/s9VVkTlwb7TyjyyTc2NVhPY2svIn7ZseoCL4b
CYqoDrBiUvzdkkdh4R4rLBc75CBZ1kJEohy7znZ6uVIbWKDjfeN+4xiC2lypiYmM
/pQahT0n2SMXg5yxl24XtmiDqn8ZtIPCwwxE6PiHAPV6OPcpT8+Si6PKIkbwIrH/
IW8uM3FcqJmGJ7IMpYZ5r4c5e8T3JC/rj5aCpHUmqzcFpWETQvkV0ls4JyY1rnaH
qGZSW/ptZdMTfIaEEz8Sfy6E/grAy0cNvKfIi+xXIMxbQEb//8tXcmOzfhfebVTj
fIeq4lGEQRU6qWwtwfmFnwMM0ZfZkex5jbEljd5kMbVoseXY3NeCfc1BjtsuwSFy
10vnWC/LA8VO0ZMgX+OhoH0z98rNfjpoX4sszHnoyEcSSZbMP1gnrVsRw3RkwPve
HnhxIZLo1PVFUDEY1auoWSXIc1TLIjr8bIn8nzBk5d0q8LSI9jb6IAYJ58Fwik5U
e3aVJMdAgyLRT43b6mOvhwqEXonUGwerU61ceFYUQhdNSKnAT1k+kj3Nb7bx9c1Y
zvgFh+v0aGvYt88vBakLzxx3c+AhKOn5HAyefSiPA/8I6dorDaCZeM7wkspbjvyR
OrJYvyZg/WC0bDstk3pMV0H6rd9v8JX2xowRWI8n6LMgyYk5tWXSyQ1XG8kbBjjQ
6tG3bEAHBJwUk49KatJTjvLjfU9/U1og4420X3MAsa6gto4j2m3l2uPhac5B5qJJ
TDE0MxGfyFLbmOtBSE8hz2l6b7aCEkCMBAD9y+bhBuXS7rdwvUUJ6ac9tK58wcmx
am6ILohDwKUyKxbd/JnnW7eJgYS5XeyY5HACTWaVuPcw4tCBrVirHmaisO4/CU3m
JmXw2KFY+GqjZLFO1BzZeLN0IaTsNxkVBrr5pPpSS3RBParZ32QVk6CvwapX526q
z8vzCLikM5aQd7wYsD8OW2XIXo1Q7wO6plHMZ35bsoyZBRZD4f+o9YoFZjtbZ6oE
9+lKMWj5jBFz+dGnkTzf2c2leHfv5O6YEqONxWWMhIGTgQEg5iZjPGtCBk3bBvVi
gURVP3UdP4NTUg1/mAxUHXj2VbEIbPyfjpyxqjOQzf78DD4uWh97KIBqUwCzhFJS
NTetE/kfClQY6I3wXDQUCrgM0XpQYFLI/mEcjdggNoLRD8TnmN2kDfWbQsptLLy1
yhfcPceW2u7HGZrBEdljRKp3tGWdcRK1XsOm92zqjMxQJkgfWRfbefXJI/yBdgWm
BTLt3Xh3bwcBOJOjuM+ZHetSpaWPf5Qrx9ei0onkOby5s4Baxg4m2TT2sHOO/NXA
NTwe6VCT7HJDtC1u4ObBojpWAIUPSnjQjDC1WlQyn6fZcC1Dzr2cU5KEiWeLqOXu
K7oeWoUMqmVWgLnvz1DQUhoRPUh9HKV+sxNViRAwXiZibRVMqIrxPhKjubwN4ouQ
lC/LvoBjS6RLdemO7NOya1zzFXlDy/7E7Z87yynINUpZBgYERpc2IjqfEWp/jXO0
Ba4GpdxryVsMz1x7n5F7ro5QtVe2u1nYe//OmdRNFfFoIIHBynj/nKU48usseA2q
aRNRq7tdScbzIBNNinBCNFmuAAt+zVB+WXeOXmDyNRLgvfzys0D/f7WGCjoZBagQ
B9qD7Hk7AklPWCdZJh3JtmCD0KhJmw5cugvI+LbSGHw9yY9BgV0wb/VMto+mSXnK
DME0p+JrpZ6mgrlzDNe2OhVFgaXj58EzS4np/jY70b3pXSmDDXeRluOaYFQTWaKd
Q1sGh+jLfZU4ygOiWOCVIgH0b+YZs0Ks90aZfPyorWmbXpYDZHekx05tNQKCJXIR
/i/mWXbFdwIi+t4ig6vuRn5k+pbdIbSmKXeg1igAxzufgGvjX+wxRMZgIpT8g0M2
oCYf+6b8g9U//KBmitCR4vCLgDuuEBgmwausFg7EWoExXt+FUbxRQJ/GqIXFnMep
QSUSJFfjMKBlcCTCIMO2nYcBuSrqvElG1AuVyqastPjk5EkcnZQEiMPoelK97nU7
uu5fTfFm2k2K53gL8lXX/dkMtS8+uUjPoDWse1TUQg9tmrpWTgG+vwlpvOxtIL2D
UAR2S139fhSO7zECn+Q39/tf/+6nOu09wRRrDy5hyd7MOIJw0Egk4nUbqbbQC++w
CjK/w1T3RJsxuUOd0ank0gcbu2B9vrqMUu6d/mPt0vBdwKZqD+dUfgjlZrsHMNcy
hM2CGPoKzgJkTG2S9cq4wVk7HqY5qwC1L/O+iLNV23d0b/S2KvxUjqgKsEVdo9Vv
iAzl2wfoAyGnl8nQoyu+CVV3YevQvspMelTOdmBrv0kKfWA8SyMEva/RUc7203ad
sjRr1NCJCcmdApuuID0CCBtjXQbQQEeVH3+MCwC7/6NLIIEnHylnFPbvCAFLJKM/
hZgI1d3XNFZuFds0VENtxcxZ5+N3tyzG+GkAfwCgfhgTQAhp1G+GSe6GeHnEMqhL
Qpe+Lp3Plzo1og/gA6Fsxwumdj+ck4gyORLIRG0mhfeKJeUSyp5nJmCvNIeXzS0F
t0ZwRG1r8ud/YJ5qVVd3xsBq2yemIwc6IttAV+PD0VGgW9zJbLbW+MEXsxP7UoG/
F6ScWmq2eElGPZuxv1YUbinLBFRqmTvugBJ3VyjJXoVmmnw4GTarP7Cs3iSzOkNI
ShPuL7ERniJyR5uS3aYhdrMRK1VqwwdpSv3cVhaRmHKy2jRB2CJn9rRNCtnaM8ip
meKwDjKXmz7635wkyUvhCmc4i2x9J+ixICl2lysSOVBtB5L+LpJ2VA8NAvOTtuh8
oMoP7XUkDfVC5EyVipRy4m2fCHyJzBWvoiEWnGvwDNQQGS170a50w69BqKqXNe3F
U+kMHIq392gx4FrrXK2IocaNzwDM3m8uP+6xBAaP5jdE7kXRw7sdZSPIWmIA9FCN
nGeW0PrN64iTuA+ecKM0SEEf5KUIbZs8AmX6pasACbpzOSlC2DgT6SYkYawPW0hV
2ZyO33vfn0l6wje4ngRl6jrTzCwFsw8wOW1XcjqVbq5E4Hb29RPV++Kbze5h/dpV
s8sdhBE2gR0rxr0OUWSzbRdscVrFsds0l/T4ClFCJeSJcguUT8OlJUzH6ApnQVSm
WQ8oA4C0o9NvUioOFpEgqIcyWJ6282vpMWNN1gAOu7ibSyJ7aRkgNBpn9k6l7cK0
O0nH3u1MbLTKrq2Ervgc15s4IwCkYSyKp78DaVSIgl6lAqMKdvWyiXJvpisdUiJ5
DiEqBRpW5lg4vAdkxKAwqdz2RbM1MZBXE0FAG0GE5DlqwiijhWhcW7Cw9o1DricU
tvnzRDiRExv0SNElatOVeGuiQDpJk24BXUiFFbeOcXBohrkZ7tVkspkYixL686+/
hrJHxXdgN3Dk9i/9zdpJbGyZjtYr8vU1hXhBOFLbnLm7M1MOWQmgBA6pol6Kk4Ko
Q4JlEPeaOTALPmhgCR/+2PfLWfVYVA3uq8F91coCy0q0H2zoyfU5NhYIV1/ZpIgq
jbxPePbaigtDpBRRvzCFeRzfAxA7GwtefZfJHfopYt/AtyayqHM1Um9VUKHlgJjb
NvY+qiBemcgq704d6RmEXYgMiuoQWpS8nfEgX8TWHSXuwjVQstxSn6OdNxQlMLNK
VUlivzkiYdLTZqnWy9ujnkXV8UrFbORpNLZYTmRZBSGTJRE4QsQNkqQVQBDQzPOg
A3+ImOLdV3W454rL6r5k8QUQXAmu5Y+exQ/sx2MY/536/IsdAzFMo6QXzCzf3Crh
0miGhlcGLRUwyfIya8elj/CWof9MtRALO6XjjIPdPT2NYcnyG+YJ0lMDVnnwMYKx
VF+6UR5OH57CXm9c5SC3t8HaGGWEnZ7XLts9E9/g1GqPHfYF2eTfD748pwFfQbi6
w9J0nTP8exe76TE+R41v2vOIvWMYUQYDeVWvgq5dksaFuGiSrHjIx7WBN7uQqb/5
6NWanslUarX34t+jVpcgRghEOO9stq+mFIJJuqrdDWogx0nZ4u4zVZAuLd5AKUvo
vgcWbp2o0XScMCkpH8c9/ZablTy52Y0fC03OvzOo9EsdKv2+ebFg9ww8kfgpmLQF
fSQuDcQozVkKmG00x/D7shwxNL9CZlJAUcKCLOTt4O7zwjVYJKs8Rr/8XVaZcT+F
ov+15OZFTSgEJFmHHBckRgG5QlcmUp1p4PwlfcnV9rrZOLPAcVLuj3si+8+6cyYg
5PHrfzGpi1b5SKYIz1CBGGZ7HQltVDxRRriFDyZ2i9PlNkej/RnB+kjlQ2L22848
eUZMif7VkeIkzrRT0l4rdkGAQrvuIENJhpSYjHlqKMSLWnTfeymyM+7HvGxZmtiY
MUpdueOLhYiCHavfradQ3ldvF8Nf6613Zz1HMyfPPjhkO5GCpgOCCkC68II8d9sg
sgcpGgKPlAzELpKO+SZrjCLSXxEAE1NvpPq0m7zXgDCFajHi8c22/Wkmv7qmZelo
PTMc5m4w8BT/fj3Jg/oESPrnOzTJ0uXhr6ioOlYgHsUvrHcztIG8PlnB8fZLpw2v
ranXUN1mz2LMu9ZTNqVhx8+Nl5ZK3e17xGZcpIVjvn1DspEP8uAUXS1dcdiNh3YO
hjqByecXEiIsqO6FV27CnN+X+2mBc0D+LPjeMC0fT6lofg1nuwM7ANAuFaE/V0Mv
270mfNcuSERbfnGtaJfvNFLlRa/Abb7ZIAIvHzUMZ13B8NDmmwthCDYpL//dUP2+
nszEQmzMAcEWxW6ss7CNgkAwBwISu1R/sd+nWJLjv+E+2MvtqeWdm1hxpK1yx8JB
YGAheYZZ0LOcDvCPIurgLv+ana++oYtikkZDYcRaTEkUdpFgUhMdkxJS6Wfp8dKf
VoP36d5rsjhtRpVENl6FCD/fciamvPAZXBWjMIweeo8/8Zdvag/mtB9ZvBNPSMM7
BUnWRPBg7NDV+DBQc/63mlKwZi43C/8HgCDYQiO7dwF6fDEjKqZFC5qw52YlO4rQ
6jAPzc60Ei4EmC+ZVetbZRJDqsl5Z9+EsRSOgwnF5r0PTfDg7qfuuUyO0vFfA6wm
KgEL/2pBqAXf+3EGjZq669Opnd0pfNfm3jHR+inx6tS0Ynm0YC7CQjQYAtIIWkWj
y0yVaEtfKp4WdpzMdW3V0iI+FC8VBb9CSZFM8MLSfJHLYqcE0vjk3XGcsDznv3wl
Ig8dYlJzW/vEbVoCTy/NHLXC3bhXLejnMoCdqLL/mG7K08Sr8S1qPMZIpk4U7qbu
zrb9Wp4tg9s/0RcuaLXkZetkrBoV1XcDmTr+TSbXcR/ymShIikqm/seVW2mRRTTi
9gqEc527GAhDiWOcqPAgDuMJoOGBHZpbOzP7prgMdeQqAhrDSxo4vdkY8y0LwcOK
/3sWcYcgxVmNQMY/vgA+0+I4d9WklbAX62NMsB5/oWSU0n0I6pXyUMY/cu3EJQtV
6cetsepi29i68ED4lcrOy4IxUTU0c0YVpDRJuIcVe1LyqP4t40rQm3fclJK2JVES
kP5x4xltGo27zJPjQ8n9L4HoGvWzgtZ1O1AT5H+TAM7Cvd/pALX0vVCrtLlwKUZu
H1vGOLnMiTOp2H0ZHkWc9ofUsjg3Qd/FyKIWxcilUQJbc6rGb7m62BwpUjDL7FHT
r1slWpU+S3EnEOOuZSkF/TvTnx3TY9nrfS/VZpup+24i6sH7VXuns0FWFLjoZQJs
CcVZVOcp5TWHS1Nl61lHdA0WThGZbcSZcceUlFjbTlbTKB9KVhZKieVvDqT/JYXv
JpB01fLvC9scRbrKENZTe+Byv6qGMqyMst6pNwUJ4IkidmbL8jQgAZgx33DJjn9S
rBhwS4zJhsv9dvZoSLmRlcvmJ6iCo90CwScwv4Rz2ROsOb//9qAs2fKlz97OQj/o
BhEH3TsV5aeWDpTAlQnvKJmP0RQlOikKhLaK6jiG47eZuvG9nSzSwZlQeJ63/ptR
sdNEvLLMUHG3L/m3OpPg6NKa7N1SA5dD+Oy6WzgLdLPxHpsOQecxTXo6oaECVkBu
Ahs83AN4XO5caGVrNSuAmtd58b4cSbOFqm+7TT7IUBYISu9jK78BdOmoZQXI4mTp
lnzhrmR+oexwUDs2mI748pDn0Sw47gM0IWYMwdhX4yzRRj9gfLTCuMlrkqPjk6wf
o8lSTXIEri3Y5KY09SgOLxSo3XZlVjOWrYUH5VrK1puqU/ra9xnPwbK60M1cOOPf
Sj3cpJaQM5BkvX9wU6Dgg1cLSRXPbycA/dtjhePGFds3NNjTDpzOfroClN2413Me
wNAU/Jkq6ifjIZSdclh47jT2R/C4rBf/CsfnLkCA/pe4HXGhtlxXmTGKyxA6rgT8
qFomOxRM3EC6RAM+eSp1gW72QxqVd6qTfgInO5X9cpxx03MHthYj3r6b2t/9YBBP
itHGI+lUfLn/PB2IdTuzEs5ttmWeKroUGVSXFLH+FrfaNB/U1FkhVzYQpbK4sstK
gL3FzSgVnqBr/HWTAJvWefDWNoSC/qxTdN2BA5882H41tAn8z9As6G9PJHZeu0ie
RorcwBaCiVMmpLpPm2261oXJ9wX6D6tJ5G405Xkdl3L6WEcBiq3CvVZo8U8qc4Rd
QeUINcl1rre4K6NZtUGgC3ZBYbDFTWbw8pvsvpql7yIXENujEgBj12N3/aLYbLkV
L5njpIZCaV5M3FoU7G4jw6ryqakoWcdTsq07OJLd7LrOK8ExRv2BDP1bi9APDNih
UX71TkXK4MnjsTCwbb+A7U4HSaP66SLOemCWQzzyo+m8wfxkG2cC+HjzinIlwjSX
2si4JX5btWzIa437YQ/aw8PgWk1BTvCWIAFOfc5V8O2P/TsPj6nKmZPJcCnRihdM
p4P480qz8mTAnYtfgmiVTSlo3B8BoGs5NrWK4Ver4nrI9pb8/eJ4Kjo1smuQJpQw
X/2hcOMhcmbkdCRvoFr9VuYwV/yIpImTRM4CRYt62T2KJvPrxPE7qvoT5ZwjqcIT
EunE7VtDE6c+ebac8vVvpz4gPvwkB9AwwQlRLebPitoye7Cnr0a0Vz8JxxBF5QYJ
+9I/b2ne+Ju/N96UBIXcJIkbAqo4M5KWqdQdhWqxrbo/SAhmRlz7ceMQjWW2kdt0
d3OsjgBHR/gfB0NPlIRoZAwcFm2GTslaBOgCZ1sFZZzvtXPZmA7KdPZcHyjGufZo
XVtzUcdqyl3YblDSPOTrmrJ84tN35+XEyG9BP53LCK9oog3s1d8T5yDqTQN8gP+M
hD4WmsR1aKi9ehPsGIKREyK3MhXXpUlQ89vaAPHMR/Nf7nTqH7NzLfhD2IfiIvtz
jqW3W3p5w8xVwgN3iLOeQY1M0mNrdm/foOVkBRlfm2lpa5e5x5sCkDvck4dOlEKn
lcqGsHBMSyQ1vj/EYAJCeU+lULPGKNqjEDVhKCXYheNG1XFKMzFeOysAwgCpspKr
3fCSvEWONeA/xE/vVhNhChEotT3YQDI9UAEcwYPID+AowjDUGXwwnj/JNbLa00C+
Hf7vF6V/kruTbq3E3WMqI+Gm5GRbYoP2dENvJdvoK6zj7iDxjgOE45WI1FcQvgqf
OXzrNbBa/OhrxI1j2hBZQ+YhAqYWsXDzI98jPUfZUr4lQIJuzdJDQZlQBNyOAe39
/rMIS3mFGBh2gSimL4xZNxQhByvqHaF8hUDv0NAvzPw14CbcKmxvGvMmoXsQMEkn
1bbzr25RS2/Dte0OmYCfxP1ypuOTsZ/EIndfumJT/uBXwy8xZdlbBfyaXb3rXkAa
6yaz48l6I0JREL+tz2/tcFmZlRFddy27IijqLP5lYS0x8kJn6dEgEqmGifntn8Tx
qpniYGz4gijVBEincxqjZYsLKzq8pANP11nZ9pEAWRJj/V0ex3GD4nBX96ASIH0Y
kcJeFvuKewHUBwmtC7Lz0T++zwi4zVNJCrOsvWavhdNELs1up0lH5+0Sbo0OKosn
tfFMo+LSd3ZToUNS/NDwlmGhjZX2jCi3WXiav/llZD3XdCjA9QryzhzhI/yl67xR
GcfzPJ9SY+/Z+P7WrgmcPkT9yMYvjMM4TRsjrvtbNOHYPUdpHT2TSpHq7He8uOu2
EW/0do+ACEBPrLIZqqHnqV3scqZQ/WxT2+DD1EhKeOJWne0qNv2vu0mM3LLfdeYJ
q7dhTeWwufqCZLTR0CopxCZuqdUcdmBkx6WviyMFOobjTLSXNTMlnW65z4dwW4HR
P4bdQ84PFwkHgM0fHU59TEI3YhjYjwZc41Pog74Ljlrk2ekEZgs/sLstdiE3iJkw
liJWzeW1nlVYEaN4SeUDI63zEZffgCpJjSxDYQ6JCdACU1LLBq9mReg6faU2wofh
3zx+3lDQGinc6ewxat0azzg3cvnM5Jv7SDzOR9awPsJDib3Z0dTKKd7ohL8A2uW7
7rd5FM6NVCctkpyF1pcou+DUOdKzKD3Eu54hY+s5RXC+iU7bVs2Ch71baz3LRJgn
JJ73D+L4pvsY9SjsJQ8L6y40kegk0Hc8yn/Yei4lZFRnauZTx9TPIPHH5KlPfiZV
Z4/7f+fSD5n9qgRnxw79jhq26Av69su3NQSQ7Qzc6pTD43JVuXfrTWBrjzbIyUjq
a4ZIR6dZuGY/Cw5GqL90HjtMoK8bVErTf+wQ2DjVjGdBk7CSfQqHLOJlYzQAeerj
6YQgPJVsmEWDzKePLGymylZcrXY/ZUctZULUl4aYErZr3m+17Ptgg85y5ZnXZigX
U0aGRZT4sB1cXlRhx5QpOCVmDZvZO39w3soVHm97m5xapgWswnJXgbqd5y4MZUlR
cO3ZBf3RguuxugWnDUD9zMnzaJHQ+bAgL8tE0UGunXmqaXRTiDq6SShkqFxG2ugc
WuqAUnXy5qbOo+zrYlKaTlE2xRWfaFhrMwYu5ekPJTBEqVyKdv9I7D4ggx3dbEGa
EyAR7k4W5mMAJQunTot/JsW+L8cRrt144gqwesSiusW9q5fvpNOgRtE5iwfoRJqE
xEPAGQUTONogHXX1vtHuSe+CnoLbGgaoA1tplFwOGWWW2uNBCptzL7o2AL6qM9J/
o7C5Km8ZjncoN3/iVNOftjE60AJFAZVvaekStalz6Sqx3McThXwejWhBfWmLjFqN
q/+i4Xa3DXpEYoYUNrKp0rTO3i0oQpyOVRwxF2wQZyfMhjo+SI6BQ5+cYr7uB41p
KNiG7iK6UPmpr1HVinytK1MDOe0vWW5zgMbWtxSglTzGDGiOcJqfcCd9LiKzG4oi
YN0ylg/sJTnKYm1rQGtGAM6E7BDQ1MjIUVfIeu4gguh8sUiM47epQMYjjdLML86l
ImK9mV9BN2zsPOzy6zQ2uur7N9q7nvzAeGvgcU9KYJIorhIWMiETguP2RfBEv9gr
HbCDks/+N11cCNGYRn7iRBdryuPh0hV6hBfEUReAliBw44Kj3oPRxeWwIaWiPFsP
vkKDCjHo0qivYAvUgeSvA9UlyUkB2S2xAkmkm+GJdIrXEn/j28ZaSaGaHgsR1S2F
FGKNJ90FDudmh13BunXeU//XGxkkRWQn0CbBMkyOoIjxc6K5kfcl9Wxu3lrTJv3H
iDlg3AaTccy7xWSX51XkClXKinLh0HQq2Cni2Atkb4EWckAGipmFY9XDXpRY79aO
SbCDVSLuYiBo0WjBYCOqVWUNheca+l1xFLjWmz0+rcOKsMI0EWIGOO47wYaxCQeV
Uz+AvqX/F3eU7JaR131JMXM+XwNO0Uj2cokn/hDVxJF2Si7JRxrv60q18qq3xkNk
d8lsoxNxxqA+kw2qHSGP71asZZ5hHhzZOj6jRzlKZQVaobc6aYIrpkmeZhQOy2XT
rCQmboqKjQVVwDe7Fa9u0jIXukkKbHD/HTi79O8T9Az7Icr21ppxW+SKMSoWlOi1
P32e1NSG+R1IY0Np+U0a5/U8UqrgfSCWXp3qPVomjpwtOPjIPkq+SMhH//wgka23
n07qHGq5IEgOn6XS+EKOc9W5auc5oFcpXU5XjbLxMbCB7AvI7QO68guuTeSsk0lg
tRM9oKCGlaT7kJzQR01PYSzxSlDtAyxDvMt+du99m4vGZjgrvRekm3QJR/1sj5gb
2CaNWJflo9aoy/c/t9mIKOBRkDK5aAyEc26V/qMWa20PQ9ZBe+SrqoSugDztHS3y
LepMxS1tpBzJzr2Uc4EfX8VfgsZGyWmLZM2O9xIJ+PZz7avMZmCtSX493tTz+5mL
JqiDU9Hvfb/rpMMJ4xLp+nI0CPPlVxzTcFHENXRXsLlMjs6novdTXdB67Av4oPX8
jfAWCZXrA4XhEVnanJ5WHh/l24JqXpTUutdU5bznGI0aJjmY58+KvTSDHNZLqTiz
G19qvY6EIYMj3wsGtNv93+/i/obiI64FQg1F6MHpXyFv7v97lCuI1g2qxrUhYF9m
KRYx3+ABamcOM/f7XVKkaSosjvIbsdSvKRAQJJz9WqoTem0YyedzQ089nIQXCJ1c
VYpz/7rAreXQN/Vw8rfnzUTeNF49tuJzhMnDlcqn36fR6vTG5fyFEyxLBrAktVyP
s34pPXBG62WSUe7xc0PT++FpxuV7U0GmA2tnhA8OLZIdLGAdwb7SaM06oEv0Dhm0
NkCB//1d7sdV6RwLd55iixDucBlVjeajyy2auEwIudvkFfJYwWbW31peYdGWCOF6
iLSyNUMY2EZJwdsUbMi86dwYfmdHcm/0L6dtFknFfApH9S83jAFL3pgeyh+s0myq
d78+lrnYRi4oF6WXppd1IvhzUmaCiJdvcKbyP4hxxutFcrjCTc7cOh+UxTyTqs+k
VeGpJA+kUmqCYsjvwD19TbcxhAaGeSy92OfG8Egaa0hEO1XUNzTFytpvZYMtnPnT
epyBDIURcf7sJBWbgc+cPb61n2lGw+1TDkmCciFYStT7BZ8aZQBFJJhbAqVFaMYf
NFJ/AmDCzQKb75bhAGBWnZ+34Nj8n4dWnXLdMv8B2Fp6FEeHT9nsKx+fYH+rWO8/
pU8NSxKFC9SruMw/9eYSV1CGILXvg+OXwAdWrMzb5W92BglvHFEx5+peVmjKiINA
8dp7hMPGUVzotrlb5LR0X97hxREJQUbdS06xi46mnI1gHSasmtIxRO+XoirEhgAl
AB1lWEdZ0LLaYC7Wukt1g0Qcl5CweyJggU5x71jgwfCq+mPxHsauytRuGh3oeEO6
XfRb5ji2eoUZ5UFC7kxnBSDwcusXzD7AiCK2SFfZp4SMjX13OLDVY2M7//OqP4XL
yapKSKsU3QdeA0CbeithHXZTPk8WAeq7tQForA+KXyczNF+BC5NlG5+xJIUdk7yV
YpbfgJqc7zVPg7CtcwrHte/CC3ig5jUC1OylLe+/y1WmrmorTHt5eMsBal5bWXsx
7/7poou1QlTHp2rr80Id4urbHP2g+yGxsqPQHhtpqyo0nVScovcuPhumc6vGiUIf
tRbawr90qUFYQxgdXcT4ofG9+NOdMyWwMHhCb/PTfPaiWm6ypWpsYiq0lDUlGJpA
MqVYRXvrlTdb5s+89NWl3CxTkZMaaVvVUEDeNuQAG3cLEMvJXUBAPTEw9jEFxQY8
TeXGXCTnEM1mywYV6tismyjrdaHbKFuW4b+EYXBagEwFg1UFiXs8OD1D+U9OEMHp
sScIGz92XpQuGVq4j1fhwS+LHivoldtqEGudw6HsnddocVtwFizz22U0E4vMNLdz
J6jb4QB/UPcJezAs6wFSq5bIPdeIclFXsvNDvkhMsfEEKfPB2nfelZYtf/seDj2i
uWaGSc1jEjx4MogYIaRWRya1CqdQ7O4SiIZMGkkC2B21IEUkexQRFU+iS0PLUjT2
H1MaCsE7gLcdvOwFlgGCa36TZfbIoKBDxzoQDG2dtOEljl085rP7otsCrp3+zJiJ
YTq2wRqAFbEHF7VBTrJ/B9Zan6Vu3oog03uh8NsLI1CkzitxWBvicI4UUaOJrqmp
XH9o5DK/bPrHxed6kMWoKqFOjBgzqcOdiWYZb/a+J2GlpD/NAgUeEnY2NHzLcUOv
8AXbRfdoRJLqr4r2MRsyMEVycj9xj1StZiY74OMMKMg+y4q0NC5XsR/7HnbEa1lp
vKlFIo+Ql1Ti5yhCbu+29qFNP/XO/HDhFTb6m3p86M/Co8SIIbeWhwo6+J4TySpY
lr4wV8jM+dtg7H0BFdUrSbtOw8N+dFM/SF/9QRDQ8TlgFcs60HyERyU3yvYEbBwZ
XbU/3nonGOeCrkecfXRTHEOHN7nXBNRlpTUUXV+qIIbslmcN/dgRQRwQzJ0mcMAy
PD4xOGOmogMqld1/czeEx5To02PG8ELTK5xJn3V1Z0TSzAOkFWoqYD9RyzVEMXMR
ecFxebThQbCc6AC/R799I5nCaJb/Fq/DW0RKcklWI356gX/ZUIH0YaPym/BIWh4J
yNNvIsKijYFl/9VTzANgdNfVPP7jNaGe2Pc6GEw70IojrBdY54hu1cKHx9zsIaPY
KdLlEyOhaZiHyiNyQheoWqv/IaUsIiCldSEChZZnQQHclDeyKWMqWSlGn+9Qw7ck
RPGzVswUC7M+4QP45qi/2/0Sbq3nxrvAq7CjhKTljKJkdby05rUghxcFm+uZZD55
bcWKSTn3xeXQMzDejxufDi10/swQftqBByUIQxb+gy1BIxC0OOuR6YPeRB7EYq3s
5JXmoyulmzG8YEHCjXTes1ivqM/lS0kZpeAOB6H3V64V58asVMjaNQx4f016zzMg
3VsHsbQAOFewTPP8u21c2dArsQrQuuH9DSQRcPAb/7+wJQJ2sllrVPXPRHnd0zh6
kpMxi/O3vodj+3jlDDAgf81F8nyMiNhoV/9KmW2dC4ALGj1tt9b+vT21YxujckMH
Itsjmaka7zvt6OUE3791oDfm1KsAZmClKyHmiOIR4v2C9fpNwfu1VpoBW+uEOahS
w7/RSLX44TAdkDsHgei6GyEQK0S+AgdrKo6jE5UTodxp+nYr78wK3DbMdaW3l9B3
BDHnpwmZg/4dYpkbmu5r0yGYyWCzQwpe5YeP9xvCSBefikhZ76BK9N75KsPcedbC
9BWbCk2Tuqq71tJ7+htONV3dkxQUGb9+prO9JjlJiREHWy3MoKcrDN4f2u0VKttN
o95tg+IHqoi4yhTLOokesyD2kfB44Tj55tvV3thgokrSTgzvRlmOtuI2aJQHS8iX
Fkupj6xLyRl6U+tnbAjb+CiiQ1e79YmLCk+GLzI8jjE2R6k6Idp7YjmbhdVoyFEt
FlnxrZ5ykiopAQxiDSo0gvLXFAeiwSQhOTK2OZyQTwBZEVPCRfKgAkL+BscjbjKk
r5DPTEkOP3fgtobvnjNgXl/MHC7YwO08uhhmbg5WVg0nyXNvqXkIyy22qm2qXieO
8wMRd18HwGBOUT93ib1knV6qaztzvW3V1vsdLEzGFandZ8fuICfKDm/+XDmapCv/
Rf2KY8pco4oc/W64NBhbhWWMzJOS9zw9frneOkIatAjvCALQspQbnx7coTlJD3xL
aCYKQ7S3eYoI2RVH4MUNX5bO+I0tI1wdh0W2WOnJSwitXjIqN11G36P7EVQRZe2w
EPtGNkTwIPHvKR/XVBOU1GPBdU7gf4TBotYhBlaOOpSaiGLLiRP1PhtuoCsEXTix
o3j+Ra6pHI6hYmQbivHW03H4UyaqBb9EvUncRyt/ZJ4K55iBaFlLOnQqFpPy95Rc
TixUObNfMX8pZb3YwmEfVgZGYVp0CBts4shZ9N9/tXIViHJya+qzT6D5jitF4VmV
EbztAb4XnastcrlTpCG2qU+j7MzdKx4yyLW/o2Gh8A/RmaM9JPRlelwt4225U6qU
jqlsZiMhGwpLaWkn7EL2cWHDcRDIDyjXFvYZDdxDcCIPSVUW/8eWcNLDvMSC9nLo
ID03SkHigQJQFEf4q9B1T9ds94M0tFe0xHEqzL+qBbztlPUbM4swjgxZEnjoyG7u
`protect END_PROTECTED

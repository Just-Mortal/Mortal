`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ksvtY+UuY7PJe9er/DSzN5yk8Uo+CbQh4wdAosIFktxrvj+RfgokJ6T9XDt3qzZE
SJeeizpqfYBn7AhxEcOdaVM0IF9DhcP6v2CrRuZKhSBF4Ts94jhUpG0Fs4HuT2eM
rLc6Ntz8RY64MzKM3u0PcLZNb2UjN/+mvpFsfSvaNdCXkoMtFHAmENMN2Fn4PwUa
1o35fDzejcmvKsSRTWhwwU9xI1Deb+DRwO4lSHMzaR3Nu6mHKDzeVT+bMp8/lCw0
Uo9ngrFSKwhfvalJ+XtU3dqjBKECWVXqa2h9MMN4aeFp8We7BAMEf9aqVdIZ8umU
G7PHsnNhfZhX94u5K8qAtN2fZmult11ugkyzI8m0Fv1O6vGvNBeW1hZ67iEbMTUs
8szx1tvqRyZSovVQb0BaBLQVmirfkH/p8UAKw11Xs+BDnOCJsKzwwmrP/Z4t2268
lITKf8OnAEKs9yssPOUNy/wK4//oo9QmrEUGs6a6hvKFQ3Uoxq8PscdfN1R7qEp+
eEV8lPFnLN3fMjGIclg8/Db4s8ilwaUTC4Q5g18TwI1ytejRYX3twWQ1oV2ZJjI8
kvfFPqIeaxNKaBOHd2yOtAkJp7F+MWs83xjTmA2X4tyNsVuvRaJfobyTe4dFDXfU
mChzMXpNki96w5LyFePBOj37IFeVdKQGj+bjQf5Q9x5LK0f+NAJgkek7lS6mOtj8
ORedEf13gbkFiSeT7Y37ijfbkmLD6nYwu44Ct8+jT3XGfwEq6xwE5UDNxAoFDmkw
IfX/6JIGL0Zy2kF26G4WZJ7/Hy1/yAlhCQaqX7L8V2ZRkzgml5Jc6tKyRZS55Uun
wWK9r7s3LO9WsQbsnJi6RuqQgVPaQFnRMk+YsHpkyyaEIDH/9ivLWWMmJAZGau4e
Tow9HOrdihfcHW0usoCpmUYzH9MXDjqGq9GEEX0DF0yR8R1VLs9n9Y1Wezi02KiQ
t2XsQBGOKCfkYlffh0TRkBKaGCclUIJY+FPxeI/0elRUeSN5288hjE6IN759/MMp
HPit50bSJtEM2D5P3Rmavx1S16BTWuBukitKzwL/QAf4XCo9JyR8ZNljuV6jpK7a
RRleORaN59hV9IrWIXOlo9xbMM7dvZM18CHX2lA5Pspnt1tPW2/wVPOj2gFExrjz
Kx5FBNnQcWxVXd9KBug3n1vNO2VaL9WGr82x+bmzD7uuh08zFORKeGV9hjmGw3Qf
2U41HVwK/uU/MDtukN3A1bQR2dckotc+1C50XLZf7f/LtI/wiSj+bN4P8qjJzu+r
yQj/3gbrljAzCd66SvmqjEtpAL8ZElzIlqnGvbAg2tOVduZTtOck4Qwmv3+v4M+A
eGgjWtZeLiO5S0WICSLFV1zleSZR58udhvm5plfn8EfcIvypKE9YZvXmyD/YdzyL
apSrLdS0ZTEQGxw6gFVJppNHT4V7VF08ii8VSKxVfseu6ZCusiQI8ufooFi9k58l
LhVYzxVowxRIryFAy2R2iQYyYmvvXi4HYu1rEesgYalg0SoMXlTENfDDj+620xLj
QnZCvk1W540byBpfOt6UzULIgJrHXT2M2MUU3HstfmBCqJ2ebe1WrLmyaMIw++5o
70FlCLKpIpcnLMj34RNkeJ/39FifCRHfVwE2vwjFBV9qkxFdcEnXas64azuXoEv7
3dSWGepk+XyGi2sQzFPe7NrZZ/8tduJrRMeIqcqvLSj9OGwF7/0JkNJcw9IhWd3j
Y/QtaRl0TYqQRUmY4iGZ+F4ljKW8p5Lm1uguPrc7XHkORx3e8I0sXOpydBLAv8XC
ng11YN4WwHx91+A5iGM9Ubba73DpKg2fOhHarjc7RtFKPdpi9tUq5LIQ48LqFBdS
tLEHySINHOwACw6Izo3PHuXG70/q0mJzuoqD1wT07ASDQ+3u2Yo+Lh4w5xSPNVxA
UWHZgOAATBVS9y2pCoVPz8F4DeCtB197dKdX24QZ0NmGXwXFzTzmJUJTHjYJlomy
61w/9hQUkITBtPLBQe9ClV7XEtoxW0O4K6tokV49IwywoBai8nsU8IkUPGFcpLaE
NF24tTcCXW55jlyGeO/JW3y44dRjqVCHNKGB1x19e4SZ8+A7U4BRhIaSW4F3F6YM
TYSsifZ+iQOaCjaYWEAj3WvaYck5ubrkAhqxOmu9pcppurrpOH5ceBaMBH8D/sVi
gjCDImHvMDOlut+QppKm/aLWbAkphqyPsjUNAD+0Doob70BAIZwq60lkz/vEYGJp
ysKjKjPmmaff3CBSNBq0K2ud51MmuWSYqX1AWG6HdU50wn6zscVOY4ByzJvDv24t
8zN5YRoLg2vDfkAYVR2dQcI9tTGqA/3+GadgFLAInejifDTabUFtRVO6uHHorZPs
NlSYPunKMirqR/UzdYY7OscLXnEA3P1qZQ1TpbLQbmRo9EA9tl9arBRgSPWwxvOv
eJYDAAXEpwNx6853Q//Dyu1P8yk7RvWkJEcl+wqiSz7UzpfAtrL4+GZhUlpCzWyX
XMrJHpa2nyxn7N9VZIU13W0xoLfYT3asGh+Ecn6uAqSPSS/8p3YILPEEZ4D0Gwb6
Hvgn5KjJVoTizdDOTgp10SX4gaGnoKgZByfr8NFyBEkJuJj9PwimxVQEcV1M80vv
SQgXb5J7Xzh8w8a3OuqzgVETC74NIW6Qq9KRPO+d4d9UnlCMoazKjEJtoE5+i2TB
r1Ae1ACzoxCt8utQWnrgaq5PfizljBHILucNPu6kDMfR9x8jvWgJMh0syyay19Js
LIp20iaOdEwz6BE2gX4geICXBKq1zDoaj9kWDsF5qIS2kFtqqeSUcprx34KwA273
qPd3GYvaE2tee8boO0cmwKssA27rDvPXUGbClmuxZ2Qjbn/UxJKMMdHvXk93pUMM
F2QaQfdKgR0wxF7+xxOaaWctR9LdVYISgzRK95GtbZQ2L6GLKu+ADFM1DJMZmjZl
VcCRfTlg3x73c2oCWlCY+fFi12+HYBILgMw3lSyQtR6jq+ceyL9j+5jtyogKq88T
nxXBeC+kUbnhTrxw2jhE3s3hXGv2d1pZyFeFwzqJDycIon1cZpwB0ZzfqsiFUb1y
7RAkGOyvnLCgjJSq+wlT6Ws3hGGXbKeQ+w6DWyogOaDWnT9bJeBaCQiU5EOBrrqU
RJ3ds3T0wwbc5VPrkCHmLXjuTEGABFiuZG1fSxJnsmkqM5Cdlp9Vuy5iiBfJWeLe
ObOjnP5BoIW+Py0JiKxhzw==
`protect END_PROTECTED

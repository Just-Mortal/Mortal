`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hMVyoUCx4J9koZOEGa6SmkcSNRgtNY931kGjScoGU3vSrgyghKVHKw5Jrs5WgAD6
YVAyKeRPdi0apSoYAVcTj3RRF2QRD2WvW76dfCCaF3mbv9Z1h/uv6EoYsejI+RKK
DyJdaXj13ofW5+8dGfpicXJmgQps6MIJgevKkm+mbwY1/kFTyFdRJGE1L/MuVZgK
ikzAWd9fm+Dkmi5CcKZ6L9Km3SJVB8XETuPTKR8mFVqfsmPt9I6gt6D0LcJUWo5c
Vc2obgI4i662E8zQf/flUmbemNycVobzUka2RR6GCFD6tfsTKk3a9QJ0aJJPO0ux
eUy647ndVkfrOUCA6LIvl9mekPLZqOtrwDVZiVePRKb9jhYDJsHGITUV8sABfQkO
Gx16VR9cx/h4eeeCdKHww+znGlE3aO3aXoAAwkhSREj2MUpzE+aeSnPGuHSJYYTD
dR1E+xHrvmQU5N4BQb3wJMA6ykmkLavQXdpaaQYokB9mMG/xaWz54EOv0l+ntf54
Fl9qOC2r+3WIDM3RzVZgPDYSSWBJ+5FlktjeQHfK/RSvqBfNk8vKjXKsZKRaMCuC
xafVWyFzndCsUk7bgPpLhEkBS5V2ytj/Vbe0IlsU5wTI+38B3tAjk4g8fi98KJvq
OUjjXQ6fOvfsHtLDA+VSzK6C6fVF2NBdNSP45lUXdGoUtJYJ1tsyS8aWzGXWKG/C
qlmAEloDxCXWAnxBYYYQMzoYTfopiybueCfvFXr+6G6ZS1spva+i97Y1Km34bVUI
7A1uRZRKw9KRlUP3HE5N428pRf8MiJyyOjqAhQGiupXtw2Y89LumrzMzH2fAkJw7
/Hwag+llBgvVaehZehWJrCi26mQ2Nc/RIC+Xx+v7zQ7OTKSqfhEQTJFmyBt9uqeH
NW1v27qJ4ELRNfaq/Xw1A4W7n2IgPoFGcWtcXXhMcSZDVnqsqhMvnFSpjnQL8KtP
qsQBvl0yFxTeSZtSptAkG9lv4K8gP4Dr4a3iN9f0b1/aBemiNmJsLwzLz4zdoKFG
ye3C0rZ8XvA241ujde6ROX15X9VRXeUBKfBbkvUGLl2QytKPGSWtInn3WmZyek7l
spr18UbVghozQp8P1N2pXJIvUyNLiAYt+LrXn/B7o+qkWAPZyQBVZjQZgikQEkx6
h1+xrmv7lvpXJepMnqskfi3UEr1uCyrIeEA4wEjDg9zMboktgqsZ433+4zlFT8F2
p0HASfU1f2hvYp0S8pCLQqzxTU2IaLZ6K9kTyvsDRjih+slNdytosp0C+dfXwJ+c
DU8IdHCbjTzfKCB1tj6zbzlgC5jjt3PLax0CoI1LWG2hEF0Mc3lax1gFoYH2TTxa
OrE+6WxbrXyKh8fYbvXfHzrjKRBHdUvt6Nrn5T6zLQBsm4KRwBw+bUayPWc33NV2
v/qYz89Ts4K4E5bnxh4StuJN1xAoWC9PRR1rQhH/8nmXskFxbnHVuMFw4T0y9/PY
QJN/P7Sf/nSw2HEGh4q2rikkGOI5B3nd3nOC9+zHY7ELE7rmUPUS8Yvxd8t7pCBS
zv8ayCQWnmk3XKMLvwlnGj6tHQQk5qoQxL+boH53oJxNsx+dr82cuD6GVkRePiIu
YUbp2Tv3fXOVyE4CGgOhccIKIQOvv6BlBz5z0wELldGkrNfTBfJhvI+wEtNrIbTz
nn0XabSnNQwQ9qfRPGGrohTi3eAZdRM01VQRyZIa/P37EGbjnkbctdbg1AoyM7mM
snocBqW3pHjIlHlohz7f9z8u9uOabq9Rsj+1h1kkb3kbPE7K2naD3coxL7XcfMdo
1Lkt0cCQwdbNGvjf1kv9UA1hRv+su/nnAKqGoqhpGb8ZBNdYaCVbKMqWDfDy82SN
5xXLHfHEgK4rJpD3w92wYl0fgCyxlk3+Pyfyyk2sCVm0GKJuymBXSZVIYomdihY+
W3d9Y/UgXceHPkq6gMYZN/8AoZiD7YVpN/zZ4VYRACgsF8pP0aVgR0d953pm3VXF
O3xSd5TH1OxK/VK1Uset466oqsj1kP/hYivQMgya7lrKukRBFwuHX56STNlvb0ie
gZ2qOEJi1lF/Rqq33QBTrCT6q+wUm8mDGdsaGhSF6E2uJWKQ5FE6JGt5MT2u4bsR
XBYYaEamJPCX0gNzXn7ZRfOO1DHTRlcbGCBQOuesFcpG7k1azN2ZFWQ2xCtWFzQk
3jb8EtRKW4L9TFdPqkrhK/d30XApBC2NP5f67Pan9sL5apMervRm02iQswdjHZrS
+ZYsRaWDgr1cO8W+Jvq7PG5g69ACGBKl5AB1jECe1GUQMkQ+v/rCOfEygQj+623l
1/T8Ip1JBtdLtC1iyMiEeyjRZTej4o/ruxaLmVf/UJolEVb+5PKF6YWGy0vCjZYm
jVr8a3S9WOFnFspAX4qIPFQEsWG84ncASw9V9jwrHg55NZt5SNEeuiYOFFsWydCI
2ktbZrHDfOBHtGXrr1Jo5IPK8iotsNI+EgsPsIYdLZPWTkb4GRrFTvmHLte+OXCl
37Kr7fXP3KZX6I4jOsmLu67GMVIxFdE6e/wSEWX44EevjZpnHe9hCe0F7qmErUKk
IJhutX8zTcXEPGLdKGUMhQwMkbM8FWVMNkh6kWvFtLUfoHdGcBdsd9ULAtV4C2SH
FxwGOo7ByiL+gTWCc8ZQRXwkymMR7rzWWZTiuxsupZ8dbru3ybLPts0/W4Mh2aL3
sBP82IOVUAoZHn94agru/140ql+aXvgZijAmgLTsI/S8+EetDhPacBOO2nKedg71
Td+fVusgnL2dux0ZdV0uw1uT1mlDI748kvfC8S9KvegxMMmuF1RuyMlB68kAYLhB
p3HIigDLN0GVEAKKTj9dNxPQnK7wcfxxmbQ9POhKr1rWm1vpnZ1TBJXm12aw4FYS
SXcwLy5pLtUGNK5nJSjefLQtpuhd6s3mFn/PFju/GmUoj64M2Ru5ccOkQgewru7Q
1LfLhPK1S/eXo+P7WjnGP/mQOfBHAqbEw1iwh5ckzKu6N0puLbbtA8xxY5mK/JAp
4E9KxQ2pvi2piNg4KEEtzUJQG0Nl1ydQDjwF3PJVk90wdCAkW+RJR0pMhLNnT76H
+hAAPr4Xp9KBmFoK1W6juh2c4vZUOQawmi1bZ8MRAQW89a3ttdkkFga9mRskkUNz
5is2F2as8iGuLJS4iNHobUTurlxydn9hwQwlGZwmR71A718AX9RZdu0BQWPrqIZI
B3pJAYujBfQL+N4K+JEOi5GBTrHh4yM9juVf/CsWzbd2Bk/OURxST3LRa8hqBYP2
zpFWVvVWrv+fHJSk44cNpF6yTNXvE4KRIpwgDxlaNT9BXkA+3OW0L/5uA+SpvFoS
3nZmRxymLdFwCHn4/we48mdt1FCP8w1/DOT/IDZX+TWTKDZ8cT1oQ/LO/PGW2qqy
eg1GJa3Fa2kIsppRtv58CA7rp6M0u0mvTph4F1OkvZH3/mL8Xu3IF6iiCZfx1Svm
1wH32MEqmGsc+SNzD8Ew8bdWPpitE4lrXlP7aK3ZkNi7wDP66YyLV48HJPcPJQqk
imgNDisaEXwDU3qpgrVbSkW5JvW4muta2s+t0OCsc/WR70R9DHC8/7zyMluwze90
37QKlwmOdw0puTNJ+px2J0Fdxyic2hbmrWEkydTQYgc5Mp+gDSPawLqGjtyC/5Wu
IoZSRLLDbMXN5fQF5VAkw7MgLnRz6+DyJbndrBA5Sg0nbH5dGKbpOhKFfq5nYcP3
+3qqbaLmEiBfAqJloouWLIUNhYw5GLkHC1CVaVpz/SjFVn/XOlGtMS4B/X/ugu5A
4dwDDov2nWpFhGOufuMqgolRLIc2mijBCP7EKKYYlz9Y7nEUsgjZbBRgqPfpgmKY
UCFxTOEOBmUZRcLS7JSGEIwraDAhpzW/NGlMqYDgrwFG4is5w97EkF1bszjMWolJ
Mc0LrztzA3eGmPJWaAL6XFqTmY84iaMLJEVz1DKngzU5OmEXlFqG9XfQT1Mpqyos
lwCaNWXa7LlD6o4oOjP5ku4smPI0Pd05R9NaU2bQMPNsbAXbM1LuIswY2vG14sI8
cVxMd1F4wGnXWWAUsvqUaWQQ1JMHRuhTOONz3lLgfP3FbE/Nofq6JvGnW3n69ZbW
3NPMG5SnTHexUi5H0LEYJX0pX01/FkBnyp13X7yd7LZW+jbicLy2EjiWUQkp4Wgz
XhXP8CT9eztMAmg58l5/vdNoTHg/itETVTbyCM/nLxUgOl6SsWg5MrPOcHd9SwDU
gTsEQdrynZtd37T/MECuxI/kaX/x/4vcmVj5Fx5/akJpX9XfXsGmK75XUJL5glX1
Jelr7prRVN4wWNtQSZwuS2yO/tJ9ppW7JNwTULURlLYuR0K7DZ4l+KpLZwanRLCs
FYylRqQSONupkBA8m78S1DxL5g49G2bkwX9tas8G+parrj/jcFhIN+uJ2bV9F3p6
gLYF3aFir9801sF2LSigim9FQXJ5CKX5lgxyhrbGUu5TVr1LTb2hFQktj3+4y2dH
FMRcrqZncln3/kqrr5NcxYdoGgN9IfX+1EHCVNv+Xy8CPQQCKtWdUYcSFHJKz7JR
T0ASFGjimBaZshUu1XZHQvYLcl0LDFZ9HYIfzIroLREdydtgSp2GP30KboRSMYFW
sf92CpfiwtSaEjQL5D+nxUn7nob+9wQb7+0Vz8ekx6Znng2Osm05qsDXF6dmgl7K
Wxy9yzVyLl2B6/UhaMWzlNQPVVIKwAv44rOl6ULks/1HMvu7eOzJt6K6QzXVXzJN
xCIoTnJtpOMT8KY6K04Ia+k/XErZKrB0fgJqlOerZVPnWwwJipg7wOpBvLdRVBlh
wFN9PiTcDNPULxcJZ19P8NKmGRrFz4p7Y2NrAxV9XnC672NO65Yw1waNp6LPu9oO
+/TFZ4912RV8Zy0q8BB/jfDSs8OkZS2PzSu8/za8/ygxtl0kggHJSmMQfXqP5nUt
90eORc0m+JjC1pZHtPEBg3te+slhlhEho/sTFb3E3kvstXx3DNm10BRxt+9nwCVe
kqn4sWOTH99Bubh5waRnksubq3rykq7/DoCraoIgT+p5CNdX55QfmywDyEhwJRlG
+nTPjOhbswDY1ke51B9bO5mHSm+qW91yZrZm7DCq43FbxdEFTjcb7on4GfQpxUOK
o0DhlIfY5EqCMOSYyD5hko1j/TlalfYKvwz6WO23nS5fMWE64qZHe3lO1IFiKydg
JGQUcMHgH6ryb8RbVq+qR1j+DT+2v8jWiSsEzjVCCmT75AOsMeKoL4Y2qM5I6MG6
u6PWSUBDhHZnfuHsJ/RAVhkdgXjgUhSbyg/CM8QfDUvEEaBRGbgyT0UMctadwtHu
gifolCXGRpifsUgDYT+0OJee43/lSaVj5JFVnJ+QjFyZ8g7P50LayKhmxL+65pMK
KkWO4z4Gwkbu8LJRDUD4T4RoQ2pJzVOM+LwN8IHc8x7oCUexp5u1jYbtjP6uN3vU
40soWXoEb2LBj+0TlbXVMHF1K3c32GY0ull7h2uj/0THKD8kZWw8ef6HmNKctEoN
6zdaAfpaxQKCgxChXv5tvAg00knEI/x0eruBIy2lphlG2tvTa9O6feGfDgGBPThS
pRHlF0LcKjVuV1p0wnc5IOnljtSwGLxotODc4sLupKbXs0yYqJrBRmDi6eClZIIa
8IQfdsSxJjHMasJTgjiPwnFnIe+YGyfnVBjyftLWoLCjiwnM/dQZbLkRkmCBHl6Y
w9gEtoMkHDD1J0XdoBVxrnnv1bt5vd6j0/+5uAOUDSQSDUITSQrYPm303gDmCNDC
OjsZs6/uu/1XiJ43jzwJfNUw+R8xqvOlovSZGvfhB3WlLPDCrtYxZPaSkrH8DC+W
jKF3bn6pbxTgg/XoTGHKvN5/2Eb3+Gk2k3CR6XIHWx6UbfDriyzytLV5E1Q3JZfR
yJUYT5cbtObDF7roomKpPV1EEUjdXsIQ+D7RiWcCruhAn5G90i0mivrAfXcSiwHp
KW2FbPFA22CKDF2opbRaPwwQZG0QVnkcmr4a2GuW5Umrt30vP8FdUCoNF+d8a9bZ
cSCMyJebjlzwCANpmrFh5wA3Tg2wiftZMo76dYwHaw2C1XPUp8Zz67XdLG0+n8FU
6Vx2eniVtXM58+1rd7M7lyPopaeqt9/BX0tGVupn1lh++wr6roMXH3iu7aeK2kNh
XZIagO8p5agyNKyqZ5j82nKuKBlwLP0o4I8IgFnjQTsXLqVkbKwHrem12r83lLSe
lYcQ8Bfk3jnnCj4zPG2KlcCxJwuxboyyxFJ5N0Slh1Ti/ZVnhWCecHYj9hgeDFaK
BY1ghBLaLLuOfzpL0RqncQj8FMNSQW0Q0tmlFc95HHHSnJp0InBpo7+uGPd/pQRO
uVQ0IlPWi+yHOYIjU+g8z+ozapbEmzs8+duBtaswuj3xmS37MWx2R1ETNLHkq3JR
dI/5U9mLyPad/xsIgPyYB1q0pnYR7Zo6bsUDY60JyO2jcx3FRAEglgokl+RUJw/k
YOlVmrTMFpyHrzgv8EGVx/x4UUUtBMfjpgb+uWXrpNffetGYOJvB20hzbmUXnVPV
PYL47d6IIVaiZjDezP7j88+q8fJ2gkURGkQSehhA/hKbCKVYfQgjrhQGqqslTOy9
Tj4eyHWImVBTn2syka+BG3I/jAAR+pSNhOMBs4zE5aehHi32u854b13KPQUu+0Oh
IiWlkbJPVlKfRjLqNh1fsWS3kalTM8COiCYBPuyEQ4K8nxDAeFDmLyvbg456Omc+
TZEpZPoC9UjVoI8yk7LqvEBMSkhtv1J+un+aG2DpgghjtS+s8wxLZ/xQLJj+6t1e
Zq7GJYrApaBP/AbNajOJHjwNvDzMTdWVf4UTwqtrVDB4LtbGkwYsZ99Y6ISJAMi9
PFTBPYsYJRD5qe/eT04lXrSS+egQFUgVp6RobHIPU4WRBTZKC9VICk7l2kUiH7it
mWkdKYJc5D/ua0hivk/1SDfzloUn/tjpP82YaQ2hTwNjKiLxI9+wyX1o5PLBPrt/
88iK6CChrGuz5I4Ar7ZLCg/FFGHue5ABd1wTQo6e34nEoaJwqtZaH+vDhVrjEf5T
XdnMUz8yg6HXE6Ff9+zNz1GxSNhnwk1rneNxU9TQT7G3x1+W70MSabUmGANmMGbS
HQxYYFlpqhgnm3eyo97Cyyil6FFMV9eZSLOl94ryC7DXFKwBAKOyNt3wpdSfkolH
kCRwaiwUhRNnU5AAhXsnCzfBCfVAA4Xen5+HmBd6K9ydmOyqRaAHfZhk2vvOpi01
VyFgW7VARfjpJcqFMAs8yIzBPUscZVFNVBNn59V5sgovP5Kvi+HGx7s9b7i+0Mga
7q/j3k3zU4qLqgkp3NTq53RwwHT1h4AZQo/VuF1J3PGXF22yayiLs6X9HVUL7N08
vGBTXL2uPv7CBB3z2aC3OT0WKqbb9/Jy010h4AkA6BuSGcf4TGBoCAAcitLNB4uE
vj3Xd3VT119mO6GXGBAE8LftZQcWfNWQkZOBC3B87HD5bh0+KiNWFfYcmH9gpI9b
aaO9yfp9mTc+O04DQ7Z/7YWcMBo0izjFVMpUXjSADS3s46xThGvQcX1qccTDkiQT
iXzlGBl9M6Oyp/zS9jsD19z12+P+YVglemdhd/MJzkam1dyQPPLQZL1dw+s9PZCs
mFqz5f6jzK3ogpmh19WSDNRBfQdV8a0mZHJUoGGxndKhVfU5nlmSI78Y5fvYsBGz
lo9rI5IxOw20LbJhbrFrXgLSH71E7/NH0t6z0w6dWB9EcT1bsayWMl8ssFRZml42
SQMAJ6dMR0ccFbxLZWjJfTf9rkPf8ibua4Z7aaeTbIcCkcwIXXsy7Q1xfToTXiJI
OWa0UULS//yoHS9Alk0mBGYJeXduONfhlAOh427518f3f5sKgRANJvd8NYrzGEyy
z9spqjumi0r7yTZTsMlrhyzRAMYI6Tkdp11014WyJkp4kfrcR44mNXQlkUBqax/a
XW2Dj/nSsZzUZ21Ydr+xyVBzHp9UjR8KH/XCKdlc3ORBzUQGPEx9BB/4yKN8Xgc6
joZGZiOfSvwhyQDZcwXbVPUz6pq6CwWzKaXX5UCT4VipqH0d7h9RLYWvkwUulmzy
R9NzzhhMpg8PZA5pCl5k7nsPTOq9rc5BZYCyO3+inP0hN+6soNqLtgFY9sKfuvwE
S0cSxqoAxhU2Ew46tYFL/VSf+pxYwzkPARVQ2tNSLGsN8colurMowjzHiuEi0abY
FdJkakjp62b6lLZJEnRyCmM+wNm4wFFZansEhTLubiax7qdiyKG94+UK9dMdCDhv
W9bnCq07h6LRTMil2spyMDET76PbMV5Vp7ELEQyhZpklxDU2CUEpskCs49jSWpBS
NEoOm8ESzkuyGuDdKMO0UDIwQhYThiOhMQFPlCDc6k9BHcMTEYXdvt3semYuA4h3
jRqqLDcKRNZvtw7NaoL/OhfB7yPEZ7B8P/VJlzgoEBye87v39R58bUUegSAU9J4w
wCy8cM6qewfpDzibhRtBLLpqD5TtigvJI5yolX3LWkTO9g+f2vxeTe8J20eTPTm1
eSYEaMNNakFIpLF66lgDgajzbw1gtR6+2nDROE8gQijt+g4/yWu4Wto+JrQ8Kjcq
Ujxqr5LeyvPOnk/91li9OPWp91UQsU5CfCz4MeYQVOARjq4uNnLpqkJt8cAtCPPa
GhvJWKmkWaFNwte2fg2HfsGAoeZuqvLdafCKiGppu/U+jTdDXkGq7lz8V9CfJDna
pHmmsgTXbXpQuokmXsI4AVyuYrH0h9RVhGM+DmZNeP33u+ZPu6P86VI+K1sJAJMT
Gki4qgzihRYlJhVYnZkFiJo4+h+fcr6HEd9lwvjiCX/BNBiOiJ8nzyDPS5ZEHkOp
8lhzs3kjt6U/21ju54IiakSM+mtrwywvgue2TS46yPSnBBmM857nmGcypqWwpqYG
RPVlfrJvZakHHzr6Y+GfUMbaV4cpCY9XUX5MMmSdQActlvibnGiRURpuwN1hiBkG
xElxsbLPSKLhahXKGGI+U8+G81P5rmVEFmGt8Ym2FeVmdmkOwCuIDJlAZFSU4fIc
ikTdzt/LjMugJ6g8GcBBp3QqAb81munDazRZeZMBWgP0zVUr6ymOTWK0f74ceZUx
TXNFdVOnVOTeMxOPOiLqaqAsNYRNp2OQk0RJA/uw5aDGiSaw1QXvGOtL1ytsE4yX
jA593tUBZWC+lFhGfiZAWVXLbZCUn9t+8itsVgReoPLKLpjBy4/S8vJ2nLak1Wgt
WGbtApEMXavhbBPGDTKtuiNwVKaeNep+8pLn+fLG0LdjWnG3sPh7a/rkTgu1cR/o
dFA2cIAjDbwN4267y0bDu8Ut4PwI2v55GOxHMzR5KG7Tlektcn3dDhZOTB0bVgxH
0EfP6sqrYCl3ZEwabbhVT/bGrxzQ0Nt00s6GWPiz/Ix1DVwdf7pfMeAnF/ZCprbe
ROJe9erbsqlgfckIEn/lSUzpj9FqOVkXUSBGs+Pr8SpUvdvltGdLILXNEKQawZdU
QuKLe8yO4jcC9P7epvxdoYAK9OnvZt2/mwG1qaQcWaalc5GvLsv9abaA6aU8GYuK
pQhi3+FjgTBwVQgvfX3/qczEEE1ma3Xt9PpvCXY5xwwZDJgaAe2kMdTKuyhIlkyf
+KLQIR6AyeBgOViK+KN4TFXgJPFFO1lg8x/SKnYbyZu5gI1eJrJAQSuSOOIGcXDe
xi8gRBSJfqWWQmLqsump7qhTSF+3lWne8Ez5MVYOI2vQcLyuVpY6xrlrfgEnIIp/
HrPOxS4OYcfs148tK8koN7AFln9M3+lS/rLYIDZbBRH3U7SugJCDCKrSHC4dprnm
uzSdl4RThhaErTxk7ifxddmR2QyiYaaVXcHKoar/77sj8sbYCTpwGHydoymwsM+4
VyZShH5hRn1u7MAUdPIsIbk5Mu7E3o1giEbYe2T0dCM3lpoJbcTwoyz3ug+asbHK
Ii0Jd318l9kJ4jVwT0SZH2JnAhUZOZ1qwyNCnOs3325wybxrRRjCvdtgbOgMz1DD
Bi+Lz34lZmHV7nL3BKEf6M0mpt2+tQmpD78NizGinGD24ztqRvGli6UjjSWhnXaU
cH1FzE5RRLXnWgXNSptpGYuNyHFIdo75yCW8wa/fIlcs065OFLpyJ5GASXBf5r7k
skg4bxhCMU2atVnNBIO5iB/Rdu/vjPnZYU8DDdeAuCvvLPp7Plv4r0cItffeTWgk
Zwy/J7gV0uakvbEWRte/69x2DQnC1TIUxhljYf/lpBnAmOLpVQer/f4XTUJ2UFOU
ashlOYozmGOCk0QdwfeC3dhmXEBgtpB1vkChHDAG6dfOMif9pm1DO5CItiw1+64X
oeqJ+4guyWJKQ5iL6I+ZBT6cMtdL7e4/TgbB5jPSyHXX0myw81CuisnM9qWOjBmR
TtW1VdoQ9NGNsNjxbqknbcyGuS3ppJRK898goFP3zWdfbVj+NWDifl6fGKQbUI2i
weRmaJFNAytB/bDFC8ePPuksUMTjffZIYnIHMO3pXHYy9xUbed1T2yTKk93wOm62
LGIsEuNkJ0nz34zsvy5N3EJipVcA/s2uV2cnkjijib8YqbE9MPcazQePvK8gkBN6
WqZbpXbd3mvb5xVYigeKK7tcUe1wrSxLKYQf2bK5xTN2+aTDW1/mXwSeubjB8wDt
3+rVuaGm5PFIXxkXmdKpMNMDnx//42t+2N1Ksu7h6YGkmLW2tUoc17XXiGWo5vyv
B6UhoENkCtuQd9rpHsAhW+z0FgWlz8FlLcRxD0opI1FrA7zeoxoHVGOtfXYbjRQL
T95+Oy3Y+tjU8iw0FbE0llUPLPLuIpKSE8yJX519raG1RVPNufvN0h7BqpIMqaot
Pjc4+KjRMiwhUGJjkxXu6diASvC7FjiK3sgVLy/qtAtcPuu8Dd3fG6UvPAWDqxQO
x5HLDdc49lHL7GJK0B26SL5TtbeWnlO0BEYr8Ws4glTzmBBTzPn4GejDqvsaAAhL
WLemJbZfuRaPbyeo0BVVc4DJzVqqGUjKaEl2Zj+It7rzOYc8ynNE7337UPItwhw1
wfcfBTOgGlmREKDRIM3BnN1I2sjYiyLjCvkH2GJ2fAOOdpFvJRd+bv8kLq8/GoFl
xnW2zXCO6FmfiCm2qcPeGymdhEx/cqQrlwEv9XHv5lmdYooOLauQ2GsMt62JTg3f
eHGLT/ltZ1imZLlRYSU3e8FBwm3YmizPZ+Ya9tl0kIQ/56F01n/lcyH8/ORSaYbM
MxoiWlI9x2TnJzQel7SM5mv9EfWtxMRsF4pL9ak0Y2+AjS7/1fD7Crsx7U/QcVKT
BMQss1SXiH/kU/3olpFhnJtl0fAE8KsBtPvVUPVaEgBwyPx64A/KxyHt+yZ14CqI
2Yqxzz7T2850825OSgjEhXkKPrQ2BoKw5i9H1+yu9yhkicu3b6FmOXjHWwsOzq0L
lx+FHoJlBOb5vBQfXMyYUAKK8q8GImzwNCpbZ2c6jegcWYMG3rWZaMW67JPtfO9M
0GCYjqn1hTcIVtyTvE0MRBFhzKHXCxIHH/JjnBi/acvnUPtV+EF8MAm1zXmNrGLH
juesUO1ecHSNDH8SDdDe6PCVlgJDrpn4MNHWOwETVkGZSCrWQflbKfkh/KWdK6FK
py/KhaeNKCuKwTssxNF8t04VqHPxLiz9a3D52BoCuIgqUBhEAVAgwH7f/JLIpkRe
q8YwyvaL0QhB7LuO2vLt798FpdgKbL2KYhwa/PGAnl31I2YftpR9Du2dr9RjlkNI
je4srsOb/8yAlG+VC0rMTF8tItXdcbHR8BHpbqOd24OvnPpcP0K50qRbRJPJbgJi
dGhi1y1AVjfWoLx62v0kYm9IW1arbEyedeeWDya54ik355WrfjOhyv0T52xHk1rv
K9/T5ojzQtH7Br8WF3YABZVZPbtwebeaNbN5sr3ZVo+sMECilA3nJIXd7LOhGx+W
vnBbE6Rk1Ze8KjGtS4i4kZMUlb74Cw+9bgEezSy7LJ6mTdkDzVZWmCXV58JeEPGL
3igS3Rh5lYSoHX0HRKVitHjiS5RDQ9/WJHJpRRLqpBDaab7oCWaStKTWhWvEfPEe
3DJaoD9WlUJxlnnGv4ydI1rSqgCFMZhi98ymnjw6dheJ3uYMnz5Cjg68akE6BBWS
TT4nA8ixkSe/whuLa0qPUH5OVS0ccYVZ6898DvSqW2RhzxV4c0k/LtUXW0GIxyav
ztWYNZaRPw6lDvvKyCll9UZ/BeMtsyUHy7VKh3pWjJON7zXiwSxJBsomdXWfwZYq
0hgzP8V5eq3u6HzKHyNztfzOCIkPVie+84nD+izZ1j3/DA8nVC8I4OOGFMy//05u
jfIPWBF50dpre70U1NEyDIXI42Ycikul3k8LuDKeZVur4Ag7P1DWQ8NVymlNIv14
uJnL0mohTSTNYc6D//Q8Lc3/PTijDltq14WQKp7iq5qvjBgRflXfC/F7bmeBs2LB
qgjJ4t75r3NhLBQnGXfnHelqpXPA/fI5CaphHJuig5GocPZzFdX/0v9gCVXCk2J+
sg6ZZ0orQ4eQf1hJVUNfHRO5NWIgwK0HdexS/MaymU/wbP0Mw5xCSSHFBeReEQcx
0Jx4ioasIKR/hT8t0h4DJa9gOjSUsJ6U+ok8pRe/OfEwId5GnsTikqIcSNFEErQ2
ieVlSPhedo/Hs8+ym5RvOVZsAg2bpS8L22o7GQHFaSLdYolZ76uny+7y5RQoA94i
/OKdH/5HyDHeCu1m6Pr9VjgudHnhbGi8yas9r+Q+JnGSdhPM5XdlcDlvVx2ZOw9W
oCDhWxzqcmiRL/qNiKy1m2f5mgswH4jDhD+uxTqvW2faFDM5RypXqS6lmZfjpUY/
vPvsO3ZQcxkEepQTJuox2l/maIQqWZt6YQOxxcWt1wQhEW88hvJqPQYNya0mi3r1
QUoNtAMokwW4E44lFiA+Z1v6hFFQXzOAeyR8d+YbSMvay1mJSPvA/eF5uRyqg0Xp
9vLBTYB5gqSPzKTsF0NY2bp5sM0M61vrMImQtZekiflsv4Y96MkeNTMX2If4ErnW
Cuq+arUurpDEoJx2XBAGG249klc78pycKr0VenVcD5LRwfWX2a+aEh22uuXhwIbB
TrSXc6H0jv43idK9iRSkp4TSRKyMX5h8Ko/gY7fIQ+a+5UMrMnUYgHiUhsN1ua7B
qWwwa201pTPtVRtQFQcfOnKyXXHZSSF79HWI1cXiUno6+OGlsBKg3HUMEiyfXM0y
f4v2fzn9PNvX22dtCFX2bFX2b+PlU5g0EttJTdatxx54OsmSg8V0RPFQxvh++uSO
Q+T6ALRLEidVMdPVWzF0Jc5aHLR7ghEsHtqZYZ0ceCrfdHKs8WBTmr1F/GTc1SA9
7jaU029HOdiqcsUNwFYf09b9e4J1+KJIsXJJE7ITlAAiu0JvgxFMmzUB4NUhEsHe
n2yVPM2f9ghKkq3KpXNhrYeUdmHb3X2AQ6Rw4gJN0AI7hWxPmPXJgMzQ26oRYCcZ
CS00wWHt3k15PVURJYTJnzi35CgGHwA7+MTLtGHGKg2MUkm9a7d7FbTBDvtQA/dv
bHIpZBfe0X6aBOA7nbgk7D1yzUXajominyqCfrmwngAGymxnmYyDPF78plkIO2E3
RTtrlmAn0K2nHX7sOZpQAeANhthV2Vkrst0ugL0cLj0/fDtMQ35/+Vw8OHhvMZDd
XYht5JqMesNCw11d0I3ySBduK87660O7ntWFrMrMWPOu0v1kFHSG1s/kbBt0G/8V
U8kk/Iz4+yERs4mCEV+27kYL095qbmU3KFjLei7YEN2Zq0yddbm4ULibFqO9sLgJ
+Z6qCQR5vYGxIoYRKdIfhkf9Z9C+7K8fF4tga64pglHsYmbodbIr0+1ad8WFyI+k
EX4VBfdN9hK4+/RViZCkXEZtsVutXEn/YN7fiTrjJKHxq2lGGntJ0BHxsGJ0oV9W
cf1WUbZ8bUQNenA6DA07FH/A0+6KjJDqTlJM1g0FexY3eqSKLw/RCierlWp8sv5Y
c+qjaS3H54yM8O3RGjsb/UzWTRY0HKJw0qJ6jfX/UnfaRBKGgtSXuII5VyxeAqyr
AB6ari7BsGHecpRJLqWwpsG/+x/hiRfhh7PRHDzJmTOYaznK+TO/sCzFsiLem5C3
8rGjRchaZLdh+NfhqT5u7XmKDVGI2Emu1fLSBRSMw+k+1InICFGVexVofeB0UN11
v+ZyA5amRqHY64UKfmd2f2DMBhytqPY+aeOLdSY9tICac/UqLm44xCAtpBYwKUY2
qkOOoNw0YxEach3VNHxL8mkWMXmNYLhIbktFAm/t9HomvmoaycM+NiArrTwWfloV
nLeH7IySDMIvj7Le1S9RLPvK9Imd4UqxIiLMsFMgaR/20pFPKBWRDG6338qiIOyD
sdaUrE9vgn3+YkckSw/xDFf1jwIVE6A3cmW95ICDI5QhmhjL9OxvFXNgdOwueM5z
zpKKIKhch0S/oXZATmsy5NZJLLfqJhdjRqTgApc2EkS4bIEUhFXNG5DJB/9MNaAW
nnXQBhpwC1ekD1//rtRbzT2BJ+aUzjZJ3ahtAXGrouELWEtsz8/oeULRnsi1fiad
mQlSwPWhkolUj5O3vaEZaQZ2udgUvUQ9zTFtYvv7F7l9bqYrxbUzCLGXhk5lumlM
Ey7uqWR9w6bkmfToxB2tEr5lO1WB80wcKS4VuQKpeao9VHz2frfruGm7/msJ9I4i
0rRtudspUM39C7cx80c4aOrU4880lrFMxJWhrhy+mKlQURo2tIEvoOdt+dIUWrL3
xygFentfeiTVcVFDRXDnMKs+3eDlt8OGMET0OI42JTzg9q3sCdUERmBs+oB4VXBp
yy2H+xLj+54h0holE8sfVymnYz+CAOGNwOh24Q0JAXxwWXtPH91gKTSiuoNJHrkj
CzvK+DxNSC3Ib+qpvwCjf7M/QUHTCP9Yh3BZuOp3X5L4bMoDpFTTqWdljYT7g1rM
+2kq1Wv69fR9FCq9InkKnGzT6C3Hz9X93UCI7QULbmQj9dAkfgILy8wWgBwLqEAU
BXMMD3smel+931K3D094GkxtVo41PX6eLQNT5YN2AbYihOLHodUR6a4IFCGWIuW8
d+nrT5ftG/VLf9mJ9Ifedy455TlppMGsGol7ZqfOfxrTmLC5BOFQmqaLZRup++/O
Em1Ms4OiGORxS5lnvb+wcASeOZWHgoJRen+LmMCntMLdTpgXbOSc06geKbfOm900
Ng97ucRC+543xKd/7F/wG9O+F7vHiCZHBQNtAPMp91s96QZL/YWoBXygs7BA8Tu2
3l2M00Bftw9HfDo3aZ7JWdIPoTsxYcRyhiDYQYJ5YVkYdh8quCvwCPkeg4DFkK26
Y6jZa6VeFi1JvUy2nbyko6I/Qa/5K+BMmkapH+Le7QeXz4Ab9x8niVJtxwVIBH7E
N+DVZwc6eZSC12KimGBpJ9dGx3VeNsO/9akcbwqdEkv4DsUsVZ5G7WX51I9H+uww
c0lcIfYyKfahMESRolFflC2umFtu+/cUrctSZMXsgMS0M079haagEoIpvo+2LhVs
gbLWunQPqLeC7Y9AYxB8H0IB2DFVuRxt1V2Wl5MiFhnBuYVAQJ7kkoKquqTtGh6L
vOFd5TUzMtsQS09mogMCkWywjU9arU4+V9VXqsgpdD9RrkLwHpnH1NpfWdVGZcQ4
SdZ3dy91+TMJeTpCsvn3qhPhF6CgkjWf5Ouxul+vE50i6f8lU48akHIiJI1uZp9y
wn9K7gEOCu41nBZoyNKlTo4s+2sRZJhaDpGJdKF/ajQ5cUC494s6y3kt2rECf8+v
MRouEZ02r9B4DaVdUcLTD9dP6LyIOfAGkkiVG25bjbnQRbFniXIvJJkf9WQcggKT
65wpSz0J+3OuU+FL1S84yuJMsD7ozgIHNGwHuIZflKNrkI7eYoTmS13Kc54ACecr
s5ByyyWC7M63wvcJ6Zrk+joNkFN2gBA9RVW/chPyvjJo3mcFLubLzZ6hQNAowlSR
tKyhnCLe39NnMo4s2bGwL/zOscO36RAptAzPLBlxO5BVSkpN0FuXZdqYwgAqTD97
fU0SQLNPCR1ieAEJtb2+0Ro+RdPCZ9S+Xo19qARC+FcMqPPPWs6ZUqVR5iYv0UWG
oJ5U+xum/CgcDGeMcYVBCSJg5wjWXUgRVyOodkehFbwA+UhSdmZa0K7laCFaGm3h
/NhiZoXEWrGcMJz+JfIke22kiSRuxNBeOdQRNxqVJVMN3iGyNoA8l8BExfqAth3W
8To/T2Y85YrPQ0lfrCC7LkQcWjbo1JcbAwIknPIN7H2rO6wQ8bSsbCpCtUjI4bEA
G8SWq3NzNZyq/SWH+pAbznq9kdi7HQGB9ZnedQIypcSP3fZQNCRRK56K9k1Q9W19
9ncSr0G+EN+E1FFIMTESp9Y+PxhYFKY/g/SZDpBN+n8TuKMCaeFtmUgfaarvwvww
W1dMcAm4Ainjfn0NrbNnlu2PrSiXNx+xQdqLpiHQfJN0Tvv7Hn6QmrTO9cnViVqD
0BY9rhiW1QrImJODCiBRMKmj9hCfc52YlQRoj3e5DxkE+NmkxxTilL9m+Lh2Jzt4
H9quGqCZqCH1cxSISfoT0IR3xk8zBasTjhZ+8z4XaGbtZy8KrurTPsLLl429Cseu
bIlHRnIUO5f64eapUpV4hOC6nTphQOzoQBq2MNy5WMq8SNxESwcKsc/g8OvDPItS
jNNhGLwKbJtbip9XhPLsyrgaH5UiDE0Klrk63YMg/GHv1vNaMqoOr2QVSFP8eYt0
9Teq0/zrISS7Fismr5TX+16+vL8JpSFE9NNJfSGcASy+GBP1DGwVsuY/mF8dzdvC
appo0+sp/WqUA7YTslN6waquUHy+YITC6WKDLLYRL2d/iDFXNnbhxmjfnYG/lTWH
+YE6obcz1nUJ5WEIPxWGd5j0cj7ZIk3bGuH61bcFiOBjk46T5vZTDSw90YWTm9o8
OneY7bcX8rf7BMAmVQe6ZY8lO640bXe4yZIfs6lzg91XiAvdLJRHGWTkQjNr9uVk
7w++YIAUFJDGfvGTSagnZDmMDUtq3fOfJ1WUci3uYtyvLAIAC38hbMFOUcCslIlh
SngNLuT9+EyYjfrZxK6DeMSRaqL6jNzf6A8BiDzgzjvFuN/WA+2HEbRLP0prawPH
KqmhYhA5JM/Iw9yvEsd2bWwxWql2KuBTCAkBpEY9ZbgaKmZeIo4oUMcFBiyDff45
QW7/3tgyZ/G5KAa74Ltye8lFsaw9q3n8v6OydAfD6N10H6IEUO40ujDTBZLTjLzs
DETEOjwJ/vpnh3JqKghRbSLh8vUdN+WEfNPUS342LvpCh0LUmaIhUDwWVePAlLVh
753L8cz4Ca7yoeYmSMjZnvGvZvmi81IdWG5oMNhUuzCoVtGyrjBQ76aC5bsuoEfP
MItdaRjdgJc8f2LcY6IwYzPICa9UIhgQ4EavtRDK6PngZCiXuy0IDpBliZi2cnR7
NLiyQHQSilwCDq4h+5cGYDF6rVAhPwQq4dbPjXH4LWlck0QX3qEMMX1uNt7mcGL5
+u5rLPgiGhSlS/ieRpy64JgBKuF0NnqA8JF0maVkBfprRiJwNS4jwLMPYeQqfVUH
E/dMn2tfP7TNzegGiRCMfvZjbfJlERfyZ0kZSjieGH5eRKbvnzecUsk3NcB4r3kK
ZRvgX83Yj+GOsLNpZzJb3D1cY8Ibp7XcdQl6/c6gVNs2vwu++uK5v0+3/kjiyfzU
6Njz1JXlhdt3owm/CSxluXeTC9sQFSTCQZCPMORQpMRNHy7BNEOeJY1Uwv2bKVmU
wrxqOZxFgEZYRKQ76wr5v2HuWVgGr4IMAMVw+K/1UHORKOHbMzmCd4DngTblejDk
rZuSmthM0KQ34m3dPLkYUGA88Pbt6SMYdbBdSe715tPlA0Gz3wxloc5whZg0ik5E
xj6A3rJS/Mt6h4VAnXFZmAURtgK4FxK1LE6mUN9noMw5urgiON0DfQfaWU2A8uM0
KB/6oYMKb6ldjrAM9Jm59pW7XpQpcMqQFR4PcMt2+YY3k/wdIxmzOQQqOHqKdm5z
g4zfgUYAG8B7whpxbiTLRAu+jLEgND5dElpa5gNUla4zpN+UIV+8iW3DIBOkC6rr
/LDmMy0KnRt2xtdxTPboZPN/FUQxmTei4fi+D02nIERLHDAHARtD/qkxjcsg1YdJ
F1fzrjc82GRS1rIrWWMFsMn2KxXAIeNkyn55EMbNIqmxb2cvjuVS040/N/tmUByP
FqMX4Ml+tLIajl2xIIZeY8k98xxA8exDMdVCaMw9CvNpeizKdTo/oj2IiDASqtsq
GU/N+hvMPYzoYzb6RgpG81kXFKSMrvDmr8KRrL2j6g5BZE8E1uQKfaVWz+k5IgVu
thK48mPFOhbthYqIaH1UL0/eiCzy7hOC6icGPCKBJJEITC9ICUc76YiQ6UR9jnbF
6DtxlhNoJfkvZS4+nQZjv2KVjKFtiApv+qs52uCp4DJG8jIdKLoJTI8CWaInIth6
kmalAjZbGkXXwr6EXkFvD7+l0nlPManGWggO44ZZm+jSJM4XGUpE3kbOF/NWW1S/
UdL1KwayLrw/IoBN1f1k+oe/QnAaaHpwbnYUCHAM8B765A5xtVWVSJMCWroxB0i8
zM06UvXQZeXc8bPzEJSKJAd3OjYpqyNP0nU3aCcSolgpXTxojQ6EcwJdhZiD5LXX
GowcWhB5EmROV7HT6wvLdNbOui/pmP8ILwsQkHX4gjxXVsu+CcDTiBD4bt6caMEx
GJ69/IpAGEVODckYCk2Dg5jj+5kEqONERu6MTjz0NIbx2f/v4yfyGqtTi3qLhgC0
owDy5t3LDWaIw877GvEfNBWhu1i9KeS2zLH7U2h6YKHugmEm1nzeioMNzFSHTmkM
tlsnUUu8HQVaxCqk3Uq94mYIuqnC2RwFdIB1CGiqbplkFxfDmfQOBFLzyILGQqBu
5kXjArcEc0fkKYdpL39f+JyDSm/st6m33DvBZcX3+D0rH5dAqfeninjvBXQC+nhm
Ex06l3rtZGaefheNkGOB+2CoojiaZxedAjAv369diH+9H9fVspymeVhr/+cDuVwY
IxtqcVYTYfR2bsTfiSu+XdbjWf/YV96IM/upvsSKr8eLPa1HKOaX/YSGChCBlbgW
aobeJlt+LFma0xGbbJTk6PfLUa5owlsFv+TaZ7O9Pd4s0eqOh8Wi9Wb/k6BCdcGI
4NBo0wDwNrhgEkZ35uEINadCGIvGkdlfkINprqFTv0akYEALmf0j5UtfipmQOawb
UVfVt83ZxWt3ucgKSDbinn2XeGrL6MnoqZD6AvJEEBhb2EH3PpikA7n+hvWP4bIX
l+0NMW+3ZgdVtu6sbwvujtAe6oZExdPSxJPR+CqAvu1bW02otXtq9DRlbrrGOYv0
FZQTdIZ5+VLzoA54zTFy0LxHwK2QyFbLq0Z3zrU4/ufDM1yydpa8QK3ktKqmILos
dUGKWMxJybZF9BVZ9ZazKpLVZU5v89WY95Jb1xUQ+uh94k09Ihi6uiinqiVH4uhw
zCZuXXVqdMTeuWhD37TN/7uuFGAbHLOFSEOc9B+ez5qlxlshhJ7cE0FYIGyemcVA
1oeyUc9oGmE7fR2GDZOJq0SwsPKVgZV68Ix/nlbgfWBJh+6kQJlcMRNUVId0/sXi
weMlhQs4L3BqcJuBaDCMNqOVgiCllGbo4Ia4OZRFuGZkn2yHHjc4ysktpwTQ90Dg
es98ypj7MUl4p3duul0jmxgbJ9sUga96rnumvUUGoWK9DiIfMluGDf1dX1RIgURj
qQf0+713sfu1X5R5d9jwAnKV+zuFIHTBJkTO1KpCVuB30UH8TuhqN3aMCXDvDUYg
ckv8PRjrlzO3wtwNctHyNrsgmtGSSnIRxBYnbWlxsiLndTSHJe8WUpcAebUbQL9L
iE9W0KsXOZ7c7On9IqKIVjbCxNvmkMsOgDLwJ8H/FviOkACqFr3DKqxjw1oAABU3
YI5BxoskiUy0zmLYru2nMMr272aV4E6jkwzI9BKaAm7tDsWA6GGcQJn6KywtwLMc
9jE7QQI/1TWNlugX6q9aoLRoMGQm4ktrf89W7rYw18IXfhEdaMRqI06SAQQxfxcA
rgKwlDiiz9XhpQ0DuznuRAT10whVCAVOMm4z/lhWkr6MF+Qe5BGvb+pZBmLEvVUA
CIIUaUydmNngDw0DQ/lytyQk708bpsQ2ebDi/ia4jnDYtXyPTZFUdSQd8/XaQVpm
5iuxnP9mwc+qnWIAVuyUFYNwVnWqlykwXDfSmcjcspMH7fnrwM5uDgKzTC9guyle
wjIje1n7bLprYxLj6X8XGdZo+StXHKPTE39/2WWZjFyJOAHXAP+NlRj1kbC9RwQr
Z56aUrner6hKMod/jVYXWqC9vggCfYCeeuCO6CqI/AB78cDPItGYnKwwRdVVPYFj
YHozr4L1J662RNazbhaHIAgcjjPqzUQD7Hzl5V8RGloMt/wOLYDEZ1e5lvC1sLTw
FrQsgq9ERP0NX5bCpPcYBq/lBAR+C/HXp8uIK0VM2mZ45K9HIIEmIprOkbokCysy
/km5fN75lKxWLjrobKiF32edu7EAmS1hZXWxEYXJkDGGgxDB2BYcSf7I1RMXbWR0
lb8WUtXcoLKHKuti2PJ9BcVZeq/tjy6agz7u2SsQdvPa7F1cRzfwe7/WINtNfYYc
zNB8T3aiLeioZMdVtwg26D9RVhzPO3IRnSglqM8d4qf9p6dRhWmDXbYONqL+JqId
hfGaExacmv/LVQMShGs4NqUS7Qk1W8/SEAZdMkFGLPmJSEsArty1oqxyCnToWeHj
N6Naq3k/UcJkqgW6k+at1fKhZ3oy8e9UzCby3Z2T8SX/XOntlHOV1+kiqvgKyb10
mACWb2iy3gVDoC1VBbYgBZ0uiMMwxXKN8QOLUe+ZGeH8tMm7xMG6maykMw1jdE+O
umUVHzEQEr+sxUrABom3defaL4I7qSc5BskjL7BF+Ddhm3QqP5ogd00/jsTbrBfe
dnRneTnkqU7yA88GDiw0sRSKS99+D7TYK5WDCOL/vMye2agaPv4P9laS0fMoqvws
BlLREglHCo4LK28bAIBWAPRzoTUEc/mADSwQh+fQA1sDppH/IEh9aGih/PYCCWMF
aAsYIG5wXPDP2zPtoGfDKq9lmzspbKoWqg7+K6MknFOabC66gcaQIKkBSrf7aBNv
J3XMGf/Zdr9SzVsaW2Y+UneXxwxT3qgazwnQ47BQSrOcwDev1hJNgHjKA4lvgQGs
9tbK19JizKGGe+eFltSQ+hxmGM0kSK0zpSbr0hFRzEhsv1Ll9+MZCJrx+jauNg4r
1b/BrPfZmwvAjFc/B9lWH4nwhryCZVgy0ioVP43hUxcXpdGK2lRme4R92nICsm7/
rbhUgJ+8NfIhGPdY7KK5f6IaA/XSRHOpDfTsDRDIXjPLONyiJJPIOGuI0w0VfbiO
XT4iyUzL5NLGCpBSn7HeSCuvpaiO9j7/jtcSt4C+DNaOSo2BtM4iss4dQojqoyQQ
sVjCqDBk71HQfOgW1T+DFYcoLTmxvoD5jMtxMtbGQq8JMurcJWgFOkKxrggVGuL2
aLZC+1ojZFnTRBmno5byeG/SdZXPvxpmTm0niqmX8QjnARx4CgHV2BYEKez0U6VM
V9gFTKWRmSescpHWhrr2Jxu30HA+9w/b44n34qs9brufJshVmTrKQ9sZLgGfn0I+
H4wqOavqFaUshtSMxqrF2TT1dWMDBGDwqeZxyNwiOJwbJBoDFWbiaQBmsTGwDhjd
sBptVdY/QiZS9KysiYZD6Ku2rj8q1ag3+T/04PkMLfdD4ccDF3q2NVexuMP/XEec
tvM81RPwM/IgsOtnQ/QJCPn2WGDgMvUgGI6C6wflmj/f888+fcEFFoGWKWXqQoX7
svvygYvWu240J67hPFFKDg+ZbHrI7Q6zu3P55h+dG8KZVEyUAdDMK2rQmabvqXy2
+T0iGOyzQH9k0dd5lRDxGKlUCfV8W3/6dk0zuQvdqfFaQPr8CRXGdPdoGLbSDzL0
m+h+8nWESaRe3NBi+np8/HU4kvHDkwHYIyX4TjyR7ccKbR/KvV/sB56uwc7xjTO3
S8VyvfL3f2v8qazFI/PW4UpbxGfmfu1cPRfmQzQ3hn1DTEqlvYTrQt2D+HkH3Dih
7w2kQQ1gXT9QRrnz9nxvIKDdWK0pwZrhFQ/hNlpb341Nv6VzSngSZLG08xwib+bd
YVJuEYXWoJcoH6bypCqksIfwtmBtAIYXs9GXImyEO+zau7O8AOqmbTku3/uVd5Qa
8rk5KGE2Hm3xFJ0tTP4k88tenp7f+opePzHmpBkjAf/a/3bFlp9wLig7VXwKInt0
8c0YRtDtFhUsaRk1nUyjjLDz7/vxy0l6TKdDTRjgrynCbMskVsmDl8AsPh9ygCle
WvUotszsduDfDDhAaSIJmLgF+BHYgiLO7e3pS21WwZJUr/Z+0WD3zkAwB03Uq6vp
Lr6Z8q5OsyJQEAZ9X7sZJ7ZdwllaB1ShkeAAtkoqAoA212j1Va9l2F0pCNoVxwrv
e01h0y3Wa6kYxgXY0xYrxAmT+aviS+74CA5k8GOzdvapkJM3+qtrfgtSpbetDj3Q
mjIH4+cfDkyRCeegfmgbTl15chKuBYv+u5Q9dZeVC1Vx+jqVs2X8Dg4X2T/2132l
V75a0WlFoNgDalUKQJsjfdTndWk0siTe0ECt5duvqXIji8cwB2MlKrQ03fHWEUHw
LfFvCR1V/vsTX5h/ccvLA2oLbexXOYGYuRkVS3DffMN+1SNDTt3wWHNP/ni13yyv
IwRlB3sTo242gFTvr2OtSZi62v5otcc/KQZ4q8XnosYRY/INIPZsgwJFnDrhCG33
FsD1dQuBcXU3HsuHmi56Q0vG4U+2jh0E6OE5IU8E8QUFn4mSaIhj2LZj6HJt+S6N
nrniecx2lHCWUkQpd1haGLeR/Rj1S2PProEhR3DrwAJh/BALz6FXaI8eI0CAJX0M
u0f/dbELfUQTrXkZlT0BAKJLtJYZrMSN9BeeUZ8TWiTSc1vIkB0JyXOpICsM8kno
/W2V04OueVYP2aaA6SkkBYwTOX51nTYehRYnuY973ia2HozoyeS28Ql9mEGlcTtM
xnH2XVXEtemM+9RWm/pqpqhCJOOtnSQFm3taHRhnW4StgahgkfuNjmJWJV60WLZd
exCe5BxH9BvAt9vPD1OmababHaT2sfDFuOEvFtMS6kxwER2LFCdvbJtXw/mawbvz
ci6IVUl4sFloG36dzXMfaAJD1eiTtcpRuvnnbjTzdLHb1s1l6slGGfIsG8s2pVfM
EafSXCgySA3x+4EkZlE0Chef2+VblX58iULjeYxA2ZrWkLpmo20eym7TYgf56/o0
blUR7HqjH54req+i1ofYnxjWKmD8dqsdvih0Z2Pu+jJxodEe+wPdGC3d3Z5M8o22
LKlEgsHRmgiFXPV8A6RyVRYGjBg3OPOQw3ekzsQNWxHTl8dz5A60frX6czn5lsQ5
ibRgiJTYcClg8cBxMSB4msNgALFOAMbod0UKP3osK5pfsjr4In2FmCufoa2jRJx9
0kDAD8yYfA6Cv1FEqL+CHbHP2bLgOv3Ecu4bEPly8RchIkUGS1391zsNfUxja5Mz
deNmjAro+0uWrbecKcq65IFANy8C88agBCh6Wmjj+Oeb3D1EqjKKLco267w+s8UG
e8XbZWMMpKOGLj5vG2OLtc6i+9AzR1A8POcmq3fob52JdUEUycdRM4vH7VslBdJr
wme7arEnRS7oEtCcA5E5hmzu5+kei8hT3A8o7ASy+ikvB3+v4XL7hnycwIjuiinK
T64qFLjOkV9+Y2q5vOGVYxft5wRka65SU0xprSDNNE4JHw3LU+pxke//RKiiMaK0
w+mI6sG/PWQkXaNT3Bwq4VfDQ1YvDfe3G6zFUt2LegtuRAJnX0qP/iwBPrUOvnE3
FpUznn8m0WSE8uQFcCiF7EOO+++Au7v1yZf9iTx7oJjx7CuQTFXMAtELMo1pfAZ5
BXbJ8Z/2E5E2wY7sbhZ3RgUI9xwayHvVIuBTMd7ql7bk5C+/FwTF9hWDFwMK86HA
WGYC6qCcTbJaBL5Mf8v0SxGOB1C3sp3pLM7jNQ7gt0lcURlC6G3+CliKKsRmZcno
hb1XwNl9GR4PZusQcn6i2BvLW8Ut04+wgZhEDWyRowhNcWA5Ac/3KHD01Qh9vkWS
r8fbw/RB5fNDpbjSyDBPdaTqIGd6pGLoqWbUEj0Bx1ilE4RPd7ZRW31GxWW9li+L
Q1OCekn0bQvoC98ro5tnwIteHCcpaCy9Jj5duod4x5Tv4D823fs0vNucaHpetOAR
Ybo8cgBfWz0Gh8rSYxR5A3xHJ2I9JCcVrOHC7Iz3LkTerWMzkObRCY37sMfGAgE/
45mLq6FK4s52k9VLO0JoI6in/UJkVpwPuHMiCP/VFlgyhhi4QPt2o8sXA7gVUZhr
E6Kx5I/jgj45giRxbA5F1grHV/d6a6NePLoOz4/19gDmQlxU5eWXfFBvZt3GsqUo
miFazmGpZXnEimLseosaa256JEDmR14FCTEODls14rvetw3MnxxPnjijMdlIzCVf
zn/yjkQi45isPxZhs+WY0OSUy7pijbnmMSKNE6ey9fFd+RxL2Bosn8ilg5icuJ+W
0uWHSQ/0rdtpWsKQAqTldmcmYMmWhxgCvQ1+xvCKEIOBiAd3CfY2tg0d0GCR6Cb4
OxyPg083QVHnwyNa5UDogJfnkmWToqPu3WnVrCB5KNT/d7czNbmH63o7/LZ5OOPX
s3VSbMYdEltr2sDRFT5/HF6usDqlD8FR8JAE78vw9ynQY0JfnZ4cKa44c47Mwsqo
S6bsLjYVqhzKTnsjtF1/jxFua30gm+qOA8J/+Hn0kOqaBquHbn9Ieas51Jn2s/tc
jlYyMHhb+BCf0+nzig5n7QeZK3NWLodT1XKR0KKg+G+sIwqAIgSyDXyTr2I7ZYin
D8EegCCQ7eTAq8GPyEtw2S6uY7zF3aNnVJ8UERiuzOu6bPKz5LLqZqMha5sKOK57
QEtbkBDWZZtXcUbm9piwTD4Jrz1LiBkrpXMC0v493UVlOu+epqcQLuWGlLVgpN29
cQiH6tvWmRS1QEz1kKteskTiQzP5qQ6bYkJPP+TanyfTZ3pVUccp/eUWh5UjeZn5
MxlZi0aki4KuMsY/Py+g7HI9/KerjgH2luarf49yNJj13kxEBjEranTeslqx8mVp
ZfzG1KaeknZWpVoMY/wpALXAR9i3/6w1NoAZSeWOn/hBn+/3ughE3cqFYHBxnprk
lsGGPekcuB2zHInLqOhG5T3f0GsYaVDrbPI70R0XNBNsOX7g3IajnXj3OzN24tOu
LUpLxIrAjTHTPat6o7co3EPh/ytPTRHZoJeiHaTX0HcPf3xHlAqkA95kkXP3q7Nt
o/Kr1hIMVEqPO+toAXEH2QJxPGyQobPsuFrau76lsdQ2dwOz0A8F330hrELRrgw2
FRUFTPSlOOFQZJ0eLmb4FpnF6kS888gsCDcyZXH6s8xzR5ZxzmJyflqzzKH2b8jx
ZvGza6yBkAfCngeE7d4JLXamSuwJoyaq6sEVLzqelwA+bW4aktCXNZkUJEP+t4+f
SKJ896UOEIoR9rE1hTMNxzu6PaOTqhKzMpBHnI6uKBAKevmWtMAqQeqxnAlsYDif
b8XU5RSEziXBZL/s69rK1WvnofWNgbq6ldG+DXKLfJ8FQIMbgZFG8t6I2/QT9HnE
urQisTyn0FtMuf7+JvnMbTRRMzc/BApB9oCJ17fTA17GSdTanyKag00N1oZhwQwj
94ggQ2jOASdCUJ2gefigdd9gyebcvavD4MzZqtbmQ4E2hrtSsxJ3Nqv80ebj/C1v
Qd2QfpiOyE4thiKF7VAgooqFBh4ik1QlFXXaYRq82zLvWgIU6+P1YSbNomGfYj5i
31ZA8dB8nQTgdKGB3KWPvnGjuWvXYIepsm+Udd8JND4+rsMGUgLFqLsXOSyYty0q
yzkRdIhnsfsB2wNADXtj4UDOtZeE1wCmb4jP1nnY3ZoHHkV1k5LD/2kAlq4zdLDC
WTVCQfGOWAYDWaNGzAVADxiv/QSpz+R8JDinQohM/23k2/wUASPlTc346kaJE0a6
onNgE+3OSscG+szebPpPjRc2oFzDEx7+lPZocJQexd4SWlWbbtp+rhOLzR8QTwRU
nNe9gFaGpolO0sYZj7xwGImrpRlnBVlR2OUIMkcyyVEd2/9dz+/K/xdHkDO0O3BK
jQSG6DZkpgIglVGS+0LpC2fKoZYAqdotEVS1qHc2fkZWcsu7dic4LreACkDzrCbY
carTT/08ZDtfp4CzdzQW8MF7Moaq7qOWTs6blCLjN8o7QK9i6kS5gweFhCFnq3eM
tc79dQDSxxxOeQwVrL1ff8D0BofejmJ3seOdh3/zTeiY/SfOXEa+fay5KO8+Zndp
lZKCHoEVdlZ6CkXy2ZYKvDS+LqmrbSetUWqEd7ZDNI/VftIvBNZAao7a97amhQD6
Qp/yw4QzSI6MpBcaI8FBv/LLGjtbo4vN1ZDKfyWdT1BXBcAnodNGpEjWQSHTvOb/
ibqO2OChKsX2K8Uqy9hYv2be9MpgAJiofYpAu4aPY0+1AS5r4AI4AiN/EOgingpx
x7aSeQH/mw62ABap1V/OxqP3lVVdQw/JwvF6VbKoEWfWahhFetfelEvrECVHfaSz
r+9EvMtEbKLFRlKyhD1jfPFAZpB14vNOqdpmd4TbYhNYJHr0+El4340a5eu3LIEu
1pMKnUHDvVyxk8AadaXld2K4OVu0GKMpfjHwJxO1dgvsVvEK6ZBeEHWO4LiOasy/
G5xAt/5dJsYyDMz6e+NggY6I+bv8ScyLdsC2JKD+GcxOxmHD+kkrO7ncm/mywedZ
EU5922ezLT1j+5yoaOZ0ADabLpbss67IdDunafYhqhFkZTyrhgXyHe+/421DaD2D
t6lWb5E4dTSh6EqYiCI6OuWTrAO+ZrBwx6Q/q+XKytJZK9N+Ah7bQw4DPcRSajc2
L0MGHi13jNzcpr+WO9RdjGz8yTUvcOviLdLvqqJGyQZJ+FiPTXVivQErrabqdqoV
032S6fiPEZ6cQkvYcsRbTUxhGJB2LHJZNdeSgAdnQnMSe5uSPCuYlYaZt2NyPqGU
N/WEe8Rjxd1Hm0ig8bVmgON18sUfcMgP4bDGmZgSxrNOnOprl3tWHKXwnt0fyapN
VzcR3Lxmgh2Hh8WQtm77k+380OqerE1x91Zv2ZFn4zAkW7bMExpEme81ZRf+Ms6z
8FuHuJcwYUEjFLLc3OydDs9KmXCfWCQqhDY1QP3Rz9s5YrIVPnXNH1GVTDWAlS21
PiHpI0BL2RcoQ7EFx63qIyUcDmMzyTdT552MbZjsZwk1cONF6NTCsCbOK8LplmY7
ivUV/rGFWdVlSxcbz+IE6Pk7vbEB5zBH/7DPgDC8/Gp9JJ0X+VIHLi3VthUH/4Di
7YmT/68WoMk9//H0tvtbe7zKtHRiV8z1uWsjmo3/QMlzf/ZOyaCu2IArp2hegEjv
p4wh/JBaD9+gi00dFTfwKxTiwtRa/4zUZcStRP8BhqV3Ls1ZPhwu2TOHanu47HxX
TAMgn4Wr+CWi88h1KpzYVa3Bh5BKV5/0I2kYvUwZ0cSBkrZGrwXoj9vK8+yu9LwA
UUmx+LnW6NdMF2azKVWmydnbrQCTVaxPf0O1OM2JYXjlbNofCk8OamtYpJaiTO9K
Mbgs2wcJFBMw4YLznj0G3Gzamypm9SnpuhEMq1wJ/qjSJVjieN4CsYtjHLcAPbwV
rtmUT1dBriHE4IK0z7VnfzZAQ599KJB7qfpAcpkWFI8DQuj6VaqWYsuV+U9yyzIw
9utwrUjzzlV9PHmx4bjTzY3+6fshXbLFAhi0U+euqrFthypgx6h4DCU1KMNy3QuB
uAKRI/KgHFBgw/RmkLwIr5L8TfuSW+bRrtVoNzit/0ZaYpoH29F8nZcUb1RVPvFJ
q8JmGfVZdyzNXEEhhWsaM0QlJ/Jv6lhKG30Ilg+IYK9iiVi0IEO43sBQsjVbv/Kg
3hyVd4IYSEZMzKPHl1kqJi8e06GAfb7N4eONntu1Rcapu+PYlHDX+D6p1HXdpfjU
hr7ETNUKXL86LmTHergluKVpFCNMYT1AZTQLUb9n3TenuyHgeCgaQxTlHCezIhP5
DXe9if7qtRqFqGKibVEJ6ux8zFodgOBD51t9cfznf7I8aaiUBSAkYHShkueNjZ0D
L1yp7ODJRwyKnYPMm1Eqr3mzeZIwC6iV5XpVZMlIEmkzZR+ST268aiT8DRVw5ACE
g8rVi9FKsNyD59e6eGVBod4QH74dggNRcDD0GgqrS5g5mwKyZb4FfXQKDaQpydY3
iLHiDXZCdZqN02Qz3LPNDkDGwrJDH5/jk8m7Dx3nODUxNFKntgfD19C7MkGGduk+
6BHC6G7vjW3YkGjJ8zlke37sWbkwmE7nbAmItGrq+s5l9FXp/5vEG/+x8oGwvSc/
TgZV3f/C8nsmqE2S3CIsHqXJUQDA1T3GTOuMU1yZav53WHxl1ZHxNtKDGBKi/A9U
IOa5+JQeR6uCgDZbgcOSLvyH26kwNH2iNxwX48alx7vHmcLjcava4L4exEtktNoK
JnqVPg892JMn8jTR8ehTYH2pOoOXA9Lu4Xe10xsO2XPZ+qKz5IwRCk3umitpz8xy
0Jkms0NkM9kiBzMcuNhyNxVGKeSFR0IdNO9JAn+0HUUL3So2HXOL1BTSPrjOaaQ1
CMEZ5C6OlyHFQjsqtOBX7SVC5ZIlxDkP6CVtqSdiGjJkfMIiDO9KPhWpGkRhjedU
sQjArIBUgSk13/g7c6ZCzu/xDCJtTSsEZPM3rSqN4HmNgR1BXBKvSHDPMYjykoFf
7TrWeMh6UVKJX/Ls9CmNKzr0Hb6rMpXiAaifzIi7XxOJZd3wEPNae9jatwY9WeQ8
3ibmiD7PmrVCaJGMSSPJIxOX0MOkOBxCVazPBiy20szisr50dEfoZZuRjZCsEB9A
pFd2ZS5HhMWegZkonnBtDwyxsmLwxdHjScwEsTCT+hURyVlzSBu/hRBm4MLHjLjN
fzH5uPdz6zmr47Nr1SqiI2iXs3qxSYkGQSCkN07UEcO7HTOe5jzCzGa+PtNT7MlB
TewtlChIb3B3eUkrPOgW+zXNYuTc0OCUHxZND9beRS50OEXNvySWF/h1kZSPg2yF
gD4MqGo1OukiZ485hOusf0Ri07stplpN60K+dW3Y691XyNgEswG07Ve85C5XdAfa
QuZOZCrgRmcqEZ5J7rhZSg5mlQIo47nKeY+5Tr5AfcyiffuHILNdrKLVwvYzTPp1
ETs1K03qZoBMtezn2PAHbyceUudLzbbyOYOl8sP4rJJ45tjTZPSbiKufM6vDo+rD
A4UtDNHxgU5yAl5oQWuXUcJiFI+qhke24A9C16wATsPJx370tA4GlagYWGUvPbPk
2jHEAt1HNcU9Lhw3J6TmW4owSNs/o+YX/vVT7vARPwC3TXcr7JWInO7pHpJfsEDs
55R2feNfDUFLbxYJqwCGSdnlT4oDjVEl3JgiV6J54GoiWuafLul5DF5MwFrZv3kE
JyFkAqcs69fqf/KoIGnuGuW/pJEuhsKhl8NVTeOLG6z4mDDQhGMFVbMC8HjjFtCl
p+J00+LK6Ddo56Lo5/IT0J/WkxJ/RA5dBX7GfE0Qv6I1ZmF6nglIu3nK41sCkT4F
jhFcGBz8bELPUet2g187obtd/Cu9murLYTKeSH28/g8FD/MJ7MMN1cz4C6x+uaqI
JjWP8fzqAbQHH2ijLBPDcAbAaj1vt+27E6uJEF0FV4aDRWDmMxxQNuJyw4WzTAOy
9WUHMIPeMeDwCHQq/UHebagCH5dCieCf1AKaPunH6uS+q9uydE5CTtIHhF3OGOOh
9P4Y60vKbezAE6r1px6ve9MyGJNclihepmY79FHK6LVjdc6PmN8awxt938ketgtO
oZIHQ8rgHGXJwB5OZE30F01K7zK74+pV3g0BcAw2lJMtlE/Y2XiYe/CUDzXGK/NP
s9Chebqp+e6Az1MtFp2ym9rDU6+2kUFriqJQ+6Mlnqz7k9PfEgZHTktrY2EgMqmd
U6fjVkDXOGEsxt+XoUG2b/7C558HsTAYKLEhqvtZYinY6zYKd4qtmYircmDavx4d
/0fmhtItvpAtbeFnw23Tdhba0QFllljotee3KC7Ul0V0ZK7QmZGe+tNKOzrq8j+L
9NAFW2k4Iczgpg9VSYRT6usY2kbOLRX0UPrNwQgQvmAPT2C2CG+Y/S/9gWUQdXXg
V2RMYpqmP2l+gPAaWev20Q36M4iVz5ibaadJHH5eJJ8LCK1CBQDFFE3U1YUN4RtT
ebhc4SsjFlrJdoq9eYpwSBxMrcbUElQ5NcRxk2kkXTfWOlMUejbCyArTN2YPREVZ
PqGaz0mr+xeQYyLtbOau97WF0erkxSQ3zOR3/G8QfoSR9IhHbS1vsYhWCTBUIaYz
xUAEqtH+NMmOEGZmsCSTtDZpSFVkLnSk7MlTu1/AzX8zn6rf+vcyVC0k24WZgMSg
NpG4vMTW1SoeCSPVWOWbJhZSZDpBpsiNYaF19ScnsFQUzpvvryuC2r2iNOxI6LHx
5Vr0M0BfgG76HgzG7K1XlDqpHmuHxPPzjJQdj03tRkrMdgzrwidOIKSNoD/EgZj+
bGO37HGQow1iBb77/5G/XPA7lUexNxa4etAs5Vj3QYFiVcVhi9t12b5GWeDeeW14
Y/4OsScRm0mM/5LAmJ4xS/YHEbnDb3Cgb0M6WF+sN+qZuPL8orR5irw44jXiduz8
zOrQDuUUiT/mY0GM6Z62NdjbvFnRYnjE0G1tuLLCkqU38xD9L42GnDTXUyyS7Spp
XI+qNMe+RupxA/kfSn2OHZ1fXVfdcSbca06FK7ap74HB4SWIJiDda0RxfyftsP6F
2esnWPJQPq9pLGc/1zlK7iUt0fjjgFI2AetQEKxp/L7kSyMR0pGs+qapE7JVkWzs
ZfQBLrGO78DddMZ2IRS7rgUcRqlPBfS+43vs+XcPRAG6fcMAwSNvS9pzRrVkqMnx
r1hqzrrPXtoKzItAPpxX+0dgwifV9iIeNlGJJfyPGfoCFtBb3QlYXNjeUHFN4Eny
0jae2iVy0+bVf9XVsgx78N+ivbr8+L2LUHcmmWdZCBjqmmsTOBepFvE4Md6Y14B1
gguyiRG960gj8U3TURRYGRlxaplrR0u3YvJeld1irxZBZ+N7W1RmGVsWLXavQLBs
t/uAhXvXaAfFnljAgy8MNZBPGyM9pH3F7Uv/9MF8v7lepJ/fDYeQzFEEFOsGaBjq
2ST8aXZGmOReVN42zeJUzx0dCcsgDUONvlP8oCKt9fM+jbaaNAA44cSa2A3pz6oI
vQ3/ztyxhpYiNntbc1wbqfEisj4FiocehqmNDN9Oz29JIansPyk5q/WW0TRmSXU9
U3b1ZXPM25GjP5dV/Yllsjq3Vl/cGyLDWOVrZ1MxIVB8u3dl1xiCbi6LGb35abAL
2SiP6K3zb9MD8CJ7ijyBCy5c4UX4JGlD9is6sol8WQMCkMDAOKisIbUr8ZqyZvJD
Bs1q6eu0TNogABdgDuC7JlKx1OhpY+qFeMAebS5EGUTM/MS5vytvLK7NfAodRyFt
AzWciwBkpnXUhxuMV18XJynZhZ4ivKATtS432QQSnNwatztzObGmqOL+HzpVoGkC
+HuQ6a90jck/egziJRfAHotM/E4QP1SQXyyuQlrCvLdyCXsDhbGwoTlDnjCoglFE
spcsElwKrQFy2ql2ne2u/W1JWHWjJHz3QC647fg7ZVlq/1MnpbpZNid2fcQsFeri
uOIJe6y5hN9+JXEK8W4AqRsfhAjRf2zS37HCKw1oXtSLSntvWacumzb2A/ymUsey
K2POHeDXqvmLZiXINozz4V+Ofa4ChX+55/zLSVeXmHJDiMjB/9ON3v97kcAcTB3L
M6dCi0XefC+rAMGOo8QVhuUjQkkX5zGJ6fjGOu8/mkPleAcm9EMLGzj0tNo6MnqE
l5wk8tLQR3WS+hWjtu33rKO1JtqII3EaLHYM+ogHE8n/6GBme/r4owc0H5ikbSSF
rz54VMk+4aqrJOWwb3E/xjsKz1O3F+NHiVdhGRvINDx8f7Ky4AWFC+92O1JKXNrl
RPaEA4cqlj2IqCALYJtLwOZGFkaV59syIsuq7QZ/5VqU86flUiRCZtz1HHy2dOiI
NawlLclbEQR3T2GjeCsVtuR0b3yTOirP3oVKijuxOWlMXxJErzqNaYAGpdjh0TUk
GVMD/id+HVKGYYu0lpjpG3Srxxt0bRP7EFQrBKr3JGhQuBmAZDurmPTdkM4X+7Ub
xkEvogUTYvY0kgevPeXZYmZBLhyU089UOP6yy3Y24bUwN5UReYsQwxTu/BVA9KqP
OWqMZ9G5y85qeJFyg94+HY0JIBCXU8FMk33RbvNlZn+6IO5S7ccnQRohMwQi0uo/
jw14UrurPnTIhkjtJnUp4adu8Bl+9iJ1XPyRRTdjO3HrMcNIk3z1qRoBi7d8zUwl
V5uKNJlhrpt+JZXFJcy9kmz/MZYCgjRIoEOmUsVH2uHPyJRCw6TEBHKiYAtR9Rd/
DgjFw/WwsBK0gGTs8od4T+YOVfslpAhcrLTGCFWypgfwltHDQBWRcE+SnPn18HX1
oc5eHLIrMNyk//gGr0Wb2j/lNUTzcDtlOlBQdeEV1P1bthZHxd+x51j9ZQkddYtw
suI58qwV2to6SRBj20eftnMnAYK2F9w1c2LhOTJQ51OOcc4dpeeGD2IfOzDe2WsT
4jJuXbBWUN/RZGAy2Cs11Yt1NdbUQ4eg5m2G0OgffiY2KuatM9TJaW4H787Gtx3g
8py2vd7CWF5mOH0ea2CTp8oTE3pslUZOhwgM1ouN+kg5lAaLwgU14y0V6K7mxQyV
lYkSqVl1yhOohve7w0+rjQZzeLAzDrKKlkkyb96h9ALuwd0GOFtAgNhjYKyr773w
Z3n52FRNz6dB4XFz/4Sq1cq8vY4qBEONOKpiZ25cbs43Cyn7r1zH2pX/F3QodRUv
cNjg0NKR1Gf4x7jnKME71wpaERFQqvgoz5uAoEEYilkx9RbMluwxPo5ZdUElkHmb
NjAtJFVul6feplHy04Y61QqZHur4Sm6Q2/vge+8XOnOcPyquuDWEVyVZnSwywkkq
mscwQpohJr81xhoLM4EzOGzbKalhaeoe4ecxQNImklDZyiHfCOMBVEsfXd5zQr5K
E+pPd2rRkEuv5c91gakpEN4yMJ+2mPg2hFCmg3K7ModL680r1uY+wroriI8hqxF8
leGaSuaD8fcT9TH2qzydj94WkP0lkBMz1UnV3nbn9GwmpXGrHIEjtCVR8hsKQHe7
o/YVlZeipo2iPUs4b5PBJXQ6TiiEZNF6AFiIJBupoqqj1T/ohWdrG/AKri5CuQgc
MqqWBUmcnDf0DUhldLVdMO0r7cptwmn1EN8iznxY0lJWFhSig2VhUKNJ4i6Xs4y6
/QqvnuXbn76lYrnss9/O4eTL9aYiE4EN99eB7j/lCutAF7e8Zp61c8FZKGFtAn6v
sN/eUwzPJdLyxhn6KHx4VSh7yFA0e0N/qHwphH3TumOdzr/FoxVHi5d6y0DvPBN3
b6eAFeDFExV7mGVz3jfkCtnej6u8f9KBZlfZty2ISUuowVTFiF7XH0QIPfTQv1QN
ouU6OqU/kUd4nR9ujdojZUpoxO9pgXlGkFkOvk8czNw6GZGYK0WMIAOOfl1pegyY
jtdIn/OH0B7nmTBtx/PBMrfCx7qtqG1xA06oeMQsw9pCkdFNYTVCusxopG5cKAt3
iHN9mluOifEBglXpZrzsFj0eBcsbQcyKmUFhqd+X6dsV+wonS7C+qfbeZaP2ut6n
lt7NO7PFkkXIBdTaAVUXHsQL2JRHcaSFnG6xw36fFUv69m82zYTpJ3B0aKsNridl
YVhC8a6C/X/PegLLrpxk6M5cK6/spBQj2kw8IKmM9sWnhri3omGMwSPBNSFKAbyS
DtYDTHslYey34FFfgLe8OhpB8BarEVFMhHjAMn6XWhCxpOQh70pI6uHpz2VlKM2N
cizIwmFFxn+ahP7jpjo2NBiwareZ7Nv1yRwbYNWDARPdHcTbDpvyi3kv+Tv04Dyg
g3FY9OTPAxgP75/5DN+VIIrpCscgBMDjOMR//jD/rLlM3v64j47YypTFnpdnxanh
jiia+vVbOKzbKaHXNqMPpXUcAXhBsPa80aSqdZRsCuD1jBttWyUsXvhYHb8vxkfu
V9QKLM89/AXmHPfcWVq4Pqs7azdg0v33wzSz77XS2BXQKuR0fDVS+pm3lCfgeYg0
mEgaP8m3FKf/BitXtLekkqxphOASd4DM8faJdw9Vfx0sEJnVU+s3+TzuxdAFqC5/
mNUKhXHyuZj4oQaa5mbhcaUP3Y0S2ZN42kn3UAtZVQ+pr01W/auRtxr6TcZcnuNZ
ou2Qa+LSMDfAbuj7hn7hsixca2JcSoVj29da1RmNpeiTYavIcsadk9qLmrB0mCbZ
eBnHE0N5ZcAG+ZR+VcMQQJVJsvvseP4EhWPUiXF50LsnFJJa//+hmKSpvAYHbXXq
NSDtFh2ffQaWMHb4elpXzjDbFuv2UUd04wsKvaeQCvBJ2LHcCZ+eaMincBXnI3zb
VjwCiha4cp0wGSo1GHOJ8H652NfMfnBFd936wDI40KXT9TQxOk3360pTq0GrcuYe
tsfqW6/zxDQKKGI+/owLSoYm4iXvkjMVAm/mCTspd+AZFXhDMrKHibg4AGcVAjsj
QYdScpKB+Jie1uoP198JiA2WtM9OKh8zvcNkm1j44Y4mVFF17wkggn/n7ul8gMP1
BkvXVENKdqS/3fj+4vK0TNT25QM/53odrk0A443W5N/5ayKrD97Hdv0UssfscB5o
3BbauyZhoTr18gl54iyuBKNUyKc8KDhK/j7zZBTFY01GFg11ZY6jWQXfAGfYKbWg
x3uTbznJV5Y6G+deaKeNAPMiQvhFYbaPK7EmGTE2PLQfHWGfbGuD8WMA+dyFiBqG
aoCbZzKxRSe/c1vwA/g0L5JSY51EgHPCz5F8VkGpFHxSmQOIWJQqiGui3/K0B6co
BwiR/rq1CgLemTWSrcLJpepAL4lMJxPFTI7LNiD9DCP5hzWebW6facQG78sB9XD2
Hgl4G6aojUwZmz3tQoKD8KGRUasOiAGQ2LrMLSvPkCZ+9YHzlcPhhA9kb0y2Dk3S
2jmRLWcZ1AaTfREAAs/RJy5kGMPd4dKL2qsp37JPvSIK76kt6Bc7CA/2hUhx+LW0
7Q8ihToky0nrrBDe79BToEAnqASHmDtOC+U/8iMSY9r7rsKne5wxxDvvaob7Y7rg
wsotCncw8GOvB1H23NIIxHYeN18Nbt95k8rskNyz8eP0uqmcgk//R6QvJ4pDVvLe
gNBjssdKOlZeYau/dLzRIXrAZKxsuzuU6VW13FN8acJOmcqNDmw6lq2PQdfvLu5v
luR2jNBVshhe60UXHI0QgEJaqSd+u7JbSxJt7BZesDQu0Pt/uNusGrb4RrV41E/P
Y7xuMCXTwVgiTzkta1X09+sJ41MR+GN/Zm1pnfglVnw0VhooBqPwB7HRKR/Qb9o7
pPVrKO+BUbMux8YLxev29A+ob1m5+Y8s043kDG08iJvy38BK4mFiB5ucAEoLq3Nc
1Glhlw6wqcRqILy9YIx3QZIXoi6bCGdajaYzIWPMwnsXjbtMlJuCNOrlufJxpY+b
M+NvW5aHVAskkCgKtFJ5i6+fZuXJ5Cg3Ke1itRkeIJAYZuKF4145sqpqKCVdMq74
icKZFvxs5uehM/eRyCzySn1dv3lNBJx87HXrwcgVTDxKnfVEc8g0yCVAKriti9kJ
G4JIdGG6JHREhWS4W+d9KA17Q74/pkI9ynFCbZrp7rqvV0rfMN+WLhAh58KxaG1D
D91zY/HWn4+tfbQwgWAVIgQWiJvzQl7RmTCjJsiKYprME1iuKoOmF6MIFHAMauvY
Fuuc216zTHfNPF+p6LEv55slMDdVbziP7kD3Owu4ycC0ohpS37njAEfBNPYArORC
HuuR8D+I2RPPGpdTopj41su5jV2yEmM1xWtM0i2CQ4AruNPYl+80dJtf1QlJwWIs
+QFU/5b+Xz25oYNCOplWSR1CV8LqfiJfmwbNoFCnuN8U6GMWZ8Kjro2Wjm4q+w/E
otz0UQxC2ZZAEFf0TWj72PeengEDI3YTSYohwrPoSCtsMMVIEFNHgRUSbBpSDMqr
vjlJJpIAxQRNHWDBtU0zwAl6q+RVseFH/RWQBfSxWVqhBo7aqBGS7Mj1rdFBDNCv
AVbX0jDBQ4PgdqWcRhvlsk1wClm5Wf0hK/ZW9VowqfXcryesv4I6wz1sEk5cAiye
p1U70L8SzcMZGcswuaQn0ZQjJQJmvUCxjAK9aJWw+hJ8EF10Ld4CWnn694ZXDwR0
af1CMxInInFsetrMT57REp1fTkxFwLzozOhN1ELpgJuilmsokBArtNchbPQslqOZ
rOD7SRIrh6fWn9ooHKrEdzZsSDx25xZFrMeK6jf53sQYhBdwJOz++TvCKAAgGpxW
k6++k6eILzHsIZRVouZXraF6OHM5pFmQcW4Jt1m+O+Bdop9BFShL5vEwljUv1+uV
3Ph1+4nDLbwUeufOTA9KZgQIbgpkKm2ldwQg5ZquIxV9HnwHVzo5H//iHBap/RDL
mXdbiYAPSDJRjjuIIhYmLfE50e26NEAOXhaBBZRUKtlArBp3hv1gT0ryQAkPmIxs
LT3Xl26WZnL8nV2TfW6utVgxRJk7VELQhe3q7xTR0db/YOr1bYW+lXcnrukf/lt0
wh/WeX387irCZC5eCoE+GVly1dm5r518lu7WPgJCxO/Yisg08KCGG1Emu8t2/22Z
hiQUXlqukRJMWSLIpYHfR7JJQBpN+Nexl4scBMm8gCbt+AboxbRxE24WRxR3DKX8
EhesxB89EWPOOuUcH+5b0fgsUcnmIvX/v/v2USz1ng63rqzgJpRmfeyTs5Ltr+IW
fyaoIh5kJWnwBsM2k+1DrzN7TpyRHCW4Y/nBq26xLcEpxnAM4cerdrP0NYltL4wN
PxHPbSYIWE9YgTShC1K9+z/DZ5SpzGvBkbHu7H/Rq+7TWo9y0UJckkhBMoBEVOw/
XOvO5IkMxllpXIPjv3crXN8UpL8smifhC9fQUViE8SYQEbt7Va6g4LuX2DtkNAHw
7plsSnv8PFDwgW+UjapmSTN+D2T5SFqTe8dCgDXXqlFIwF5BjvstGKRA48eC31o9
r3nVl6U7/351LO3bwG3VwWJcqBuJuzGbc0BFFu/1Dq1TaJY/eSJHO9CMWXGzNvdY
m4J4+ETWfHLvRrMsg1Mzqk2x07M0ykO35xfc5oBlJwMiyixViWVJmOqb/OIxTbSc
OePj2L8NEUbMm85aprdxrUQLhzbecwK1Jsdbf6yCDWqnA1isOsOUVQ6m3wwcS3xs
fqEvbfUn7ixCC5m8dQlILzciJq+feA/lcg4IhZQWEa6445HnGiVUnFbNh/1HDkEc
rb+SqCXywrXy31EqibT4b+9aJhSRa3nHvt6gCMiE2Z2Ve+9pezEl8S125WXK38Fp
iPHfF+ysmrJjFQvoF2k3D2QlpIPUipzWwed5FOlussTGLMZDwE7L4qY4RONITn9H
1Xu0H5k0hENLMtPYOZIDdWJRgpN8QnOquzFAsN6sIQ97tzYiN9OsGj+ywdpxfi2n
6kz6Qk9phMWwrsE827r1Rb0W1bdTORrTl+xJgg/Na0V+uA+Lpy/8ksvsdAumcXEO
c1894h/K5u0gxYzJ2+m5j7hKoBGm0mE3kD328QPOQsAQTcOimEiLcIHBd+iq5suk
BajmM5Uhxufd486ACapSubo9fopBXHw0cYjHS6vHb+OHkBOgxjdevG94sm67dBjt
N6u4UZVm6DZyViHwSfjUvjIhiQxTLTratcqMXx2SX/REoTfh5n11XeTChpDWFqiB
3pi/wJ3B1Ykw4+63/qItps1cWy9ViaJXkSWu9J5d5KOIaiT3pyoB5z7lYCRBQZpG
SP+TihR0OA2Ji5YmBnlrLw1fST5I3XUJ6F2zp5GOUZObR4RHdAv5opkBh7h329lZ
HCqejxNKXDAT2D7+0W8YeepoLmxCIos/aPjJI1x6CvlQn+MHTVMmPBYzqec/uQU2
ngnyy/2hZCZo9OFm6uXETYveTj021bckX3QUpm9P7H45ZZzyaKMZpaOaaXIQ93Jw
66bgNDwXGTrRo5unZRBVqTb5L5Gxhb2428Lig51lJ04xMRZaKdkK/rJSeE895XrF
BQArtgAZDXQNxwOuxnJmY/24JLuZ+ciQvkPQkDdtQxaWkSuzfkxU+YeBbSUSfooG
pwbIXv7NMICXnA1hyv/9uLxChhL7/p5tqw5sisI2pnC6J1n0X4Y6KRO4ZQqhVVBw
w42xpN9fGQg/I0UImqK+Ca07m7wOL0XwqVIwW+zYDXhShJttAMoNNzHbegRf4p+0
jFUgYoSSXJtIIYo2YBHdJ+27o25g+lLWi5YeZBd5E4JBCuW4eBC215jEewR3wh36
qccRODi1+TOG0XD1NA12Sv96ha0YxcQwvbAv7ulOhLPJRNDQLb+oiQtO58D5crmx
HNWWsuwD3qTfiI6VzuIyWSd+MP1Co4NNA0Rvl+adlxazIzSZNd9z/EYqKRVmRWFl
pL/uKXjaVjFbbYvkI/+CiKplrMP8JbVelkx9IanrKMASamB7kOJB/I403BneiMv1
qTjASu8hzXa+wdfwOlgeT02p0VNFTsDP1iA9gkDtnC0OQstKUCWb5JnSNeqFy3zV
j4JAXqtw7ZfAa1DInZaGmbWnKMII5OqRkgMhE8TAL5oq0NI4Ywvtp8vpxa6rJkce
tqgqDVAa5ICOCDmuHr2qgNW4p4fmaSENz9ZsWVKh/NTlC5XVH6ov+PU3Q5DkEuQ+
3psNr1EQwnHvDi+0QwCJTuQ6/fH4Mty/tinmFw9qL2qY+7RbRxl7z+RTGLMXpKHw
WZMeJGJ9f93JxOiEOFeuImqjlvy45jvTO9d980JWUN2gtCZsorwl2PH7TDUNi+90
HdUFD/f2bj98SgZ3TitVkiVavS0w+qRgZE4DTBsd8cOwyX4strJXa4y5bvWjG41V
2BHY6hCqKlxzYWsESvFRrJrZpLzmQSVFHQmNoDo/YGVpQDCGJ0H3lQZ1n7MD2ev9
PhXfps41RpGg+lZl8NFKzbWC6gSEpf1KDbAkxj0fCGu2lAxVnmKeXU4gXw75rlKF
8NvhSAzt51XfzgkCMDPTJURZncPMIsykzDKPJRRWgk6DqXKFbKbx/tibJmaYbzKU
fsQHz4YFmUW4NTbuodD8+hXIZCmB5zf1C0KPj4KdouICqnpKx3FIuN3VGIn+FBeo
DD5mztGgis6/a9786Y6DQyhZlZj62Kp49ZZcHxY5IFn3cop54fG/LzeLm/saFz7G
EDDlVKksATFLsMY3kPQhyyifbrN6s48VgMdiBbrJbpsw3bB0KoXQBpftaiPxdzne
AYV0ohvznz7N9f7JvWGnVx++vkksrMLIPQeOvKBk6SdlPYCUhxRkwGupd9p0fUpm
NdH8cxJBi+UeOVvdFjo4ntrvt0mk8S/dfuEKmjT2cexB5whl00A6jfU6oA97DynK
r9VN8yFiyFINT2Qi35j4+hF8FbmSrUpNtCpWgUxQu4m1SRIzm4Wx2dAGtFPcV40P
eSzIFwMQ7VYknpF5TgCSg6uz2tBOETAiH2eKQyXd1kk6kWaH7xqMq19RS7CADFHk
0A5tnzGcktmfVYrqk0HzW4W032236JtpqbKlvfv/qFljLniyiW5lw8EIX8gUIGEt
ne/+COzvZBCG82lZaFFxyQMKjpZK1zRwuffxMrN0nCIrayhYQ06Q4rLDiBOhfI/b
w/2n/fDl9kdVps21XpOePZCWgSon7TFs4lyyuA95CCl0AjDSdGMFPJKtGKQiw54F
SVLzXYjFEDsPU7KXMhNBtbcM9JIqhi412Y+9e1cy7oecCkP5slXj7ELjJxARgQP7
fG4giUW3qgMrBJSq7AjELu0kRVN43aN0NsX2YzcNbSjYqq3BDdEn3g0o5NA92gB1
hJEBxqWvpOXSzOPWXszumim1Jn0yLu8pX8+hFY6hvTZe/lMR5BThNi06iYO7xaWV
gnst8D7UtFq/jU7GX2RP3aKmHGVBQsv286wOh0FhdBM4XZkX5noYELd3S7Pl1PMj
waOO+jnQD7UDOM/xecx4EGyAcWEBN/7vAmAmdynxeCBdfCloAEeeRi9pNPruMeW4
WtqtTP7n5XfP8eVk+uhs92Fzk16LL8Wlsw51WSd+a/xgKiDUT908PKXPqosV5I9W
MNbazTkH7pwg9immlVfxCpqI574Y5XceB7ul0ugIQVdvo15viM/+hLWIAy43i3ni
h5cp1Y8N1Jo7m5w/InXxN4Q8P8v9ZHVwN+LDXpd/9+kJRzKmAyx3G2NtGCowUGym
rOPoYgDQh0PaO5cLMJr3DJQ0T7mI/d6bgxsIiaM8ykue19GFCEbnusDgp/q77N3T
xGEcVt3UA5m1RghdfYFb2c19hr9vqOKEIzuzoT7dYhFADLoOC4RoemsNZ1DtjY6g
6R3MQtwOXbcWvvEBVKiQQJR+WABYtRNkaCsK35Sz0jhmbSKnplIjhELByehpCklK
IrKPm0rWwVcFW6BrO1Z1doFAHxHj20Zo9l1UFatkXWFpb8kzylvgNpa5ETQLJ45B
mn/nezG0tVpF00DlHg4SufooomqvP5woW9ePOqx5TzI7AV5GXDbiKFMTfqFcFV8L
z4sT2sG8utMu21KAoTNed7Jq0cNWwZWDU+BzVx+JuIpJHY3nRfKawa3tO+lgx15z
+oYHfRZc+FDe/293MdhUABPjRrVvAInwxU/q88j1yn5+oljDDIm+JN+ZuH+dsCse
lIUNPNMgtRywb/ocEjtWEjH5A+6q9lgc/wUYpjHhBPLkicWT309A0+AO2Ial1jjj
VU0ae0osKzB0o6T/LC6rPQeWy65jobucwsOSwvvwZnADClpeeAVEPYi/id68h+9V
WPMQkACufrvlsKFbD2THhKJgdsOJRxQ/n5jBYex3e9mAJGoxPHmRIspXQtGXRJ5T
f+I+gJlSvg3Prh4qHzN4ZWfJX98nn1gMIGY6n4iVaZLic2+LvUrn2NLJboLc9tIn
GDMypjGSIilfBxMjrJXtEyDxjYdXhPp3PtN301fPXqQJi0Qgj9EICkpZu40daENF
7rY6UIAUPkPQQZi3C0LvezoDyF9JUPvimUn5v+8bAZesxwJqpaOGQ8RXNrQoOlOY
mN5YpWkOx9Jhk0Rj6yn+ga2/DNl57eapzePlWlZEGDR1LY8AR0WonBTAtHlwINdI
HDzkMrrSrhLbMCkDy+wiXtk1SXbD1jhia9cimDUuSIth3ArktV1VF5zYYXzd1IgL
VE3nhMQ3Zj6WGaxRmQvuF6oasQttSwgzyf3lkctMNzLO0rE3qHECpdvZKMX3YELO
Fo3x07fH9Z2RzCXePV25x47KGCwHq6Susmp2oGVJyAOX+iCXKl5yCI4BRQ8IPYmX
q6vAsrLtQNtUVDtTUrzxW/rtlfUZlEkUsmMWQ8e2k8/wcMItrFaMZ58elCvj5ej2
Gjca7KEetGoZlkJzYb9dOyLG/uR6n1ert2ku8Tecajw7RqU1z+q1bM3Z7IRJcSWt
K60jf9Cgb8bL41an/QxqBjQRVba/A6hfPMMsemMhjTDTyIe55ZC1wsj+kGJ5TqQO
r2mX1GjYr1hxfevNrj46zlCNZ5aKYyGfWHu/G96bcXogJaKrDcuuuX8eNhzSDiBa
qq1cQRSXLLJ3NKF6+2s/FgWspWu7FWtkn3CffHMU2FZVb/FBgXvwILN1+MNkuTwO
/RfBIS6gTgyfgMrByJ3nA1osqq1U0iD8E/Ad1o41ml9ncvWq1NsYCAbpKsvxqPcc
kEE3KupwvMQEEcyr44jkJ8d8XimwvKLXsxVTU6h7zXyJ8Q5xxlWohVhXV5rR533/
ZNCwm/zg/GxJaq9GBLZas6mdt3GHj6GojStoeGv7U3IU3qBjGtOZ5y5klO4kx4px
EtRda2vCjfTeLWQsBGF9kZVDhQij34G287jdAlCtN4/XHiwVZ1di2jy7O92sz/+N
GZyN0zdgmbBDjDPDThISMCW1ve7tTA/+KVwbn7v2vPZhEYONbv7PJm93NTc0fQ7Z
1eZa1LWkKRdpw+ia8lM/GOEQC4WZBEyFZ7ccElvCiJWVn3PWUYNn6iT5+60Sg+y/
05K35ChMNdVeKF0jgHRpt1sgJLC1DRmSCIqCgQivTyyWQShnIo5pIyZ9yyjERwZV
JJylfaUZb8PzezgH+JD+Wb5YHKw7zd5ywnvaZm4g0aM/3oUc8gteNUR2kBFsZNfX
NNfJmkhaUwvuUOQct0V+PJtfXh1dGhJLupOmfjRdi/rjefwgSTHUi90okYw6Dtiz
nVRN2wnxr1kEcfCSu228um2B3f5YrMnZmAsV2kYMBqPwpiDb4MdWSHq4BrBqrXTk
vtW7xYb4iMG+ePBbLW8N6ZvVMU4RUNdOemdB13iS9kbTzzhTOwjBnmg0PeMMP0xN
0RqqMxMd8x4DSq0TxEcrLrgjWmLuEJSm/D1eIVLjnsfw8dXhl+w7e5QkKfUqsvBB
1VMU2XyfF9RWMIwBStDByNFD3FOmwIvL50B2SpoBcAxx7rUXw6utyKKbzQR8WGN6
d/sx7t36hmQX5aESxzkRjmNkmtL+e/LFPyBIGggXnxQBhKtdP1i/e/j2WIPoNu1E
ybcSDhy5VWpIs0DWZ/kAzw/vdw5y/fGf6yoVEEf19qkHCtlLn82kDR1yN/BcCiFh
h3mmXVS+7wdZKx8gvOO4AIpLsgCarpenF4bIJnAJpHkCzx8y4zsovOlnntPArsKZ
fWqx8VoOCQogBPHtMpXOKftzuDoPOrG7PpXULs8wVFHZhJwR1qblA+7i3sAZLXzw
aNVdTcheZ/21FDdRMS+nw2lVM9q0dQgjxFvO4XGejVWYt685H31pod5buqxAh7JU
0VDjjaVB7KGiLTD+6cozbGA4Ca+1erhUp9Z2ZqhW4yvcCV3pKUt2nk3SRIZbyMgV
6aJOujQyBt8H7vTZJBvH32BAJ7iWTTUcYKbv++qCYN9Pw6o1gs9kD+z5y1MA1zSK
58ZxIvtxdO/3I6wCOE40ovlBG/tHCfp0z2kjlXDIZjPc+oLnDbbi8sSlhvfkBy+w
AvnsDaDDNMQ6UoDt5rJqdSKEay9iSaQJknBPSESw2QxEXXJs3zQ5X+f9zm2ixifZ
AZxBu5OnOYnGS2zwU2qO3vVUb1/SWPzqrr/WCRENn1GZEWPG9ycJaBkTKVyWx9aK
AZF5+XTW6xhuBzjI8MVXaYa6vhhMrMwp06pIYFSf5y+zzMCD2zldXuCukBmvzjrk
CTHdaGTj3emNVZJ28MPbelUNAxG0OcLvKcqd6fDtlYoroYyVq/XUcGszuICDM2mo
U9BpgCy5+519AmMLYUkbPpsVBMSJP3LrRYSY+ga5uSTwZ814WuOZxJYiDjZWeIiI
OuFOJFD0Z6NMHiDj/162pcIaO13rLRwVt96U7t/a9dFTVnqvpdpS9SCgpQt8+lXd
ZdfPeGoX0y0uDEEkN6Nt4tJuaRQvfGdbNRR1/QbEBkDU6kPlnZe/NkgrLKOhZwJP
ZoBKJiVNPDqRYJOewNNTcC8AnGdNxH2ERNUKIBippSwiRr467DEloRZmMdqLSCiz
0DU6LWNyff5kr9wlu+vHR1GKQpabNOVHKQwT6TVnM4locdWfDDMU5bpHfosOSHgL
tLvpBt+EotMLDUctWRGoegPLnwyF/8FOlhks4CMQn2wMZck7j7fy+9MLvqOlz09F
zaQp3VXw2V+XpPbBQD+OvF4K0uw9U/yHxm5tJZFz3wADzcPhAOKNJHJ/tIWsMboq
8Odgl9QXyuGuBWJ9DOb8YoqnH8sYrzB6g73SGFC2nR4Bz2jIeVpcAD+xmhRbuJ7/
YW/QmNTdaPFTWrX0xIDXS6f/ZYKk1I4t2BOt2VrbTQuihKBJ0EsddxFbhp92xPNm
cELeM4vZW5mj9VkcURjzvy/pLwkpj6U6Knft9MDVSaKtGxGB8k99DRM/zhuD6JX5
wkHndd06TtQ3BpuM9v81VqyyN0wv7ieEQbJq7YLX/QEo+hKLQbtX7XQUFTjcCYLD
BD7EwzPnRiuJg5en6MUmgdB38KStPZpv2m1ova8iKPStHIzgY8gE14Vi0cnYvPKk
d7219NWzzTZyW7CJMrpnyQiw9cvkNi0Y2Qf8dPZtMlZE9uMnxQu+h9QdkeLYUUEd
ryzlEMg82zlOkdUmqwT0Kte19xviACb6fK5hzhfG2qL2Ri4NxR0p5C1K1QDd4up7
T+xklsKD6xbKL4w4wYt4TO6R9i5Fe44JyJVkYTGk8YciMEdlOD4/lawtudGlaBUI
xzRMijSk2kwfdMNyyvFrC9algoHcIY46Jc0YvebgYc2kz7eYNLON8kHgUPiMc/GP
v22xwvZ9lVDbWP0g0TwUHhq0mk6dWdxHUSLdh5p2sQDro+q+sKiDAMZoxSp9bXqI
a86oMjAjzUU6V2d+L5wV0K970zV3lerHx55FrhUHfEVxm63p4dPRxydWsS/stt4H
eqEmLHEnyqHnKupUM4QcCZXbpUQ1uNwWViMsRDxIFqOWHZP8mUtcc/jYTqGC/yCa
403Wbaf/F4eQ07Ei8UY34B1kVR7JGl63OMCMdAra6S55IIWIBD5iHfhnup5bMpZR
lGtCSwJKrfYwvEavst6Q2ur7SfwLjfSHVjwMeDQ2PBvPERETsJcySjJtYr9TZHts
C34hWVYq/hefx7aXIKo7Sm7cc/sNkZmEDyJFeJ7RlYIgvW5cUfSxfBhE3SZE9LND
vrlmzJcbDiUABV4NLRW6JfJRaEC5KNSObCxK5iCQBstZGuEU7IBA/Z2xLAw0IlXk
NJItN8ZPQAIfqWq5o+GTG/a2K8GWI93GNoZATdrcxt3Ct74dLLqiUJmVwUOuVnO1
fQdhvPIHFeHOpmF0cNvuS6+lKT/Lb7hXqFksaFTkKAxuEDqrc9Rtukg4/+vdmKxU
otRwl6zoq5FUUXhsJIUHps0dqKw0waJuX50wD8Nep52h+YK/8a+N1zVtLX6EYmJP
HEit9grIfur+gHL8qg4+Ymquj+tsXgAnwHlRyURYCXhkcaLDQ5RcaQSzhtGm7Vuk
REBqhAIFZr6bb/jPaZWUxjollo8bazpx5xgOQFBAxANg46l1pwnBrcgiLrDKWLQ4
+6aulTd7X6hsxABL1VJO2rafjNhY4y0CUGzCocIoZVUQ/ZRcUpP3Xfl2KgC9Lhu9
UhMQ5k4L1s4ZVdR7ix7ea5jwzUgAG1mse3OHeV0FKvTwNV3/b8KMB/KA0Xo0JXr9
o7ca+8jtgXo5aSShteWuzbTpmxKofUQ+n9GJvuwR+TM4SbqlMc6RRRSzmbEK0Gih
j9MmXSN7SYJYPeczPBqDiv0VFzQF1w1ZcrOVaytSCJg4jIlU5NSPJe8WR8erHxjN
EDE20b+zOui3b9u+1n9FfAWu13vASRAem1d2RjvZEu6Xq08VNsPlMjPyoB9Fmrsg
Abp5UeKO1+gn28dCEG3pWZQFAWWYSERssCz009k3dUwjBGyoucvLQopmgmL+XrxS
0lqGbIBR5L3cvkDV2Vo3EWjcCFjmwXYjVDOB+h2q2BQfgcB+KcWxYgD/Uc+VXx7b
UnfNyCyNSwS6bDvFKRRMgVO8pyYFXFkBjzQ8j7HeVCmdhxj3VLMwvPnDhpjGk+hF
i/E/vVW7gIEtHkQrKsrhbhZlWFhTWqPfRbp8TglG2NYhhOB0cKdtQ+vrn2saeTGv
ga/uYYz9Yfge5ngqMqi9eW76kAQv7D0QPeIKyKyI8grKqcGE0ro/4bhA0a3byIwg
O1kAgYnMyPJxHIJ6iOaI4lpiNCeuWEc6Ai8afTrAcaC6t72mCCUaAf1tMXRlusXP
iFw6Sfct/uBIGdrjn4QjZnPp/urSJThoEFDIYLtVPzxV4qyE60C9z3dIYofeKo07
K14E2lqiOfZ2nEz0rfGsrhxMNc5pG6iXhFjcnCOWKF96DKKLnSbFOgcnABllZB8f
yfG91l1NaV3GehARY6DOLUFpb1lupyJtyedPY703cH//09Djs/Ph+5LxJs+JcaLV
vL99HkiSqXHBYUCeMi6VD5sW3++tD5rTWn6jqJQhi3QiInb7vVAWXks/NnyfVy9M
kOTqwd7cVj/ZJiD19W+dpvlIG0S4lv8LUeNW9M9SfyWcs2AUempSTnumQLC47wFk
3jolcgBO30U7kxs4t2kO3P4Wxklfq7HjlyebhbgrsSJnUn2/Lma1Sh0msLvmpgjF
hHTTBq7uv8QT0I7I8JbIhtrGyc+ZEYEdsnj5wW5iCXsU8IhjSgcDmkHTfhTlLTzC
6BhH1VAqG0MRDdPCaE3gk4Z9Uz0rCUTPyvZgqI/3aGEqSrs4n96RTrV2moWYYb1H
dORpXkGh2YIqO4MqRc6DrEB66jZGgSUg6diuu1rBIqpdgNJakbB9aaKnHwDWkiBd
8QlNov3p43x95CBC8xtlrgf90nqibkP1E22ZwK8+/gOx02DoZcv3wfFlvLRuaWpx
J5T8jWURXBWsYF3/Uen1lyLl0T+U3IDwIX6mks5ZAttqtwSNaY441RH/1xprGVMO
M3sSM238oElPmIwDfRsiVNMLlvBk5uWTFlAL855qR6B1cKTiyVCcM2jzEvU/xn8D
HtxufFvhz9AlKhMD0QT5dqFlX8mwW+4SHlA73P6R8h7L4MIg1+FL4tczNrNlv2WW
XUvqut2KMc0C5agrk5AAIAL2VfDruLaZEPRjjE3heuuIRmMK7gP6+VPrlg+jWHkD
qiB9kRyw845eKHao0rc1uboFTHPvQVzoUHF5F2Spg1VvSE1mjYmED8+/Sh+5yo/A
fbh4sEjPKFcXT9bJLdyi6qaXCiTSS+a1/ofFQPPZNlIVh5CspehxY0lsoWtYyAYg
1DW6A6e+dC6wwIyaEe9esiENl6BWB0Ka8CM8z1zwpcB30V80X9Yl+ofeTRQHTG9r
uzpytRgNibeHyiDPvOEmm1SIqCjvtgWgsnofENAYAmxVZsEUUU6UYo5WXUqPhcwk
J9MJzKd6IsmLztXF+x1cTqsYcO9criL3DSDXaiROLDDIM2qm9jHMBl3M7Tq6SlNX
FmmLjRVjjrSkVYLL18UOD3n5/+c/RrLxWPgZKoKT08EPJdVmrztmjY1l+6qe9qck
ogar2QLNoAO5SXwkyzQCUiA/OcC5VY8Go73yK0iEWEnlTrRvSyVbH7VR5PgUUkHf
lcK9Y1lwA8raP9y0CC1fbxTOFX+tKb5pQVxPGeJoJGmBU1lJBLDL+6bxD8bG5brh
mQBI0l/aBCx+Q7H5BhYrXagAJ8qECJOWX8x5LzDmOVw/ktoWSkq/c6CBGM++L+Ne
2+C9FSyvS4TcqHPotultCYe7O9UxifVoq45zmXVifpRwIkAbKqiCJdk86gbCGp1c
lW/mIV4G9t2XeyGKU9f4YQRQXx/6/w4Bs4QlIZKyEAYnetyWeoO01VwHHhHuP7AA
r50FCa4TgnBTG3SMrOGTGGMDQOFgI9+hq8p835P9pUS546t1K71E4QDrA5pYVQuj
940bgDLdgdQwYlzVFf4NnE/yiBS+Y6j+Sd66Q1hKQa59baxjG90dQPgFWS8H/Ju9
qeTf3PLDMgP9GkPZiKAGlC+Js5NEEj3uSRwnZphCX6r1vN+CZsDaHRRBTsrovbL0
a1b8ylhPOuwuJTkeQ/xomb3S1u2miJE3awyf5sgX0ZJZ18UfqNkwxH4OIma0cSTC
WF5ly/5RWzjMNDDfNScPlYLt/WYHBWgBSW4zNioCSYuKHO+fDxg+RH3KdzyzGJOZ
sGrxWt4G4fSAXXq54+rs39ncUk2MeBAkcCMZ2FEo223kztcFkkXgBC5rHAxe5e+0
LGDcM/gTVY0jz7qxHYfCH8MTVi5woUGUGBm5FFhjv40Injg0fTAkNlrh9euCMht+
HoZ96+bvoVVqZNExSBhf+VY8RS2tN5vww5uiXufJIJSIrmQ75vGYZtYzztYLUDuj
SiDZGDJucR8R4YD5EhbaUIZp6MPR6b3Mr09PoVR+jAmLNiVXyS8hEfByuoFxywow
eSvmLhR4YsK7NfZddTNbokPI1/0Lktq9Rw16HOVT2F0cY3Xlz9I7842OW0T5u3+H
39LZzQAajlk2bvFOLmR6sBcDulA+8PT+zWJHTW8gQ4pJa2LMnm+QHOjWUh2Pf66L
LXsGxsF6e+JPDbFbJQ09qVP0nU1V5SDlOB5sLqxAZ1X3SPatWdBqtXmDinQ2+G+Z
RjmT/c/ScZBgNLP5+zAm8h9qsdEy6S4X1MIFDIhR6YjTGesSYAi17jriuCooW8/2
TU81NjRLyKxr/MRLA44IsbQoSIlNxF+8asSgUMHMlBSU36+8VCsFdZS5p04ZTH9e
fVUwogo7Ip6cOAPZgykLf+bTlJ3Keo2Goa0Dyy8ihsVx7ZkBjCiM6wIXsvBAUIpI
JuDM+1ORM2ywdivFIVN2O384B4Ts3tvmZiphPZ0h6JVfNjLaHldSW+jwJtVDt0CU
kbLCTzbEFzZ0yxS3rzWBF5chAU93TJfVYgvGwZpi7cD4TKcEXiCzkwZUglyr1mUg
8/zjnADREMzlzpm7m6RYaUVP9/4aEjpM3YbTYZURTfUlzNy62hVFx9aEDbkPVzUU
PSJhlAo0Fgsv3fC/Y/9AyfwImyRstiNYBqCB9mKxXfHYtDg9GEE37hdllmXhtsZL
x6nh1xs+/PKSamDcTNnVsE+eqyj5wgKOl0opGEH6LTT69+I5EfgSAcatd+w7HJTC
i8lFDEXEC8cvHAg8Y0TvaoiDyC5ju5dAFHd+pld/IxjkvGxMVRvZSGhXIPWHYeFk
uH/psAcJgANYjO4ALWKpv1QNCRS2+xflFsk5tQ0bioObcrsoG9qusQIC3dlq+IsJ
aWrjZ9or47mK9BkENve3o4WbztWwh4ZAyO4ETkjztHw6l4QLhnaeaIXPvtddOzrr
Lg1LJOmU42+fT0DaVhlDnj4uEpSe3go/V9lc2WJnFL9jIFNtz2v37drGigR7YNja
92KIKpMH3RKS3H5lazjJlkFRH0jCsg/Y0opKutj87DzHESTRyDzGqrWWfRtA3h2N
Nyse4/WaSyzhA2a6mLEduijP2BPwemZ5vcz/6kbj/0LkTRli4NTcfws/vcWHWh4L
NK9Y+EjA+opifjSbqPAc25Fm9Jaf8HKzK9pZ3AgwMk48y6GlqAUEL/ahgbaImQfQ
OlvRtVpY+fXy0w+wDJ7Rtk0zHlIWJ6rPpS76Iqevl1vQBfRc9kTAU3Ap7Xp2QtPL
i6VkQ7iqe8GcJkoqaEtOPnA4ovSJLjzGILO7Tgj8y2kom+neM8iAggR/zhNHv/8m
o1HFe91891J88AO/vF591kF2Lm9V5wR6xzwMxNKM1GLIAojCm4u+KO0bIvwZp1K4
6LFtn2yB+tQqmKs1NC2Jv3eFxc2+uEEd8JBeYU0WzCYmGHYibJcto6wy+WJridKT
35ofr9GfEj1KBE80Hgafpjn1S2RVuxqg4MzdZH1XCcA1mTNwLSloPAseJzwpuXUZ
hd8oWkvAnyEzabltcyIrD1XTpJV5UTUk2nmWFDIXamPwsuoY9P91kBk8NJlvzXfY
gDcS8jsO3oANYt4zr2R7jTPsSuYwdyFti5nYv2j3KC0bNuD5sbjLOmye/+uJTH+N
Q8vNp7rKIETr2VGj6hr241fN+6OADTPYoHq+2xjdkUtmq5TLe0rdv+SdPvGzgfbV
7WITksL7YdM3uRX4JYOKjw4hAXA3GShzbxfmb14pf+f4x5g0xB9yl5JqKro++O1F
NYSymFTbruyx0ZxH14k04lEOGx1jRpaehnaZS2K7n8TMRdTq873RUSlzDlbX/Du4
0pb1vE8xvzBQJZnlNWo47o48mCxgNMnJv5JYNnT1SXi5ECtCzQ+0mefCzA/mmt3Q
ow+hcgzl8XGCqUeTceJrEPCwnFsIqnV3lmaOYLoIm/9Jlgte9MygyXj5MsogE1Pe
GyoXbwQMjbpfirDRPkgjSnoMq0lT6GmJEewvMv7GOhHHcUmhgOtW6obyFS0vt25G
ea0bPGQhRggOtJl9E7CoI8c4n989XMezlkpQFHReJS5YY/iX2FF3Pu/Hj92PajEH
3uWZarfzRm4JdI0BnFmPJ471KjxQyG5y90Wrpyl/WjCqFj749mfBSm+8jNl6tBot
xasOfbF6jAFcJMd9tH9Ff50dgHb8BBJJSJiIxZFZGC/bO0TAYSJmrEqoj8CmJZG+
FUo033GXgUGn2GFjf6T730GL7mNFIQlShA6xW7KOzvuMxkqTngHwERV+lfxcmM7t
OqnKKFEOyjfs4tiduEwg5+Z35PknYAOaRjA6WXQZe8ONo6aIMeN/K1HVuQqFiWo2
Xi3DcBoG4YxHfMhjL0KOgMPxjfYaOVcTlpMnA1FnVkHuK8Iu7exjXJ4wFieGdylD
RmCymRNruPyuotcgXJXEgy99v3RcltBUyR/o8D5ZpfR7tKAOQnfbM2ye8jNMCFNZ
uP4NF/937/KC8jykAv5DFsmr0lDHtFUT4Yfbztwg5SmIwHnwKgaOvQe04KVgXYe8
YFIhQRKMOFvnlLTkNJAO2pltfFKeY3tsEhHHrYjyty4vDVajQ8+DmL/ZIPJ++CRP
N3gxLxpUxpFrXPNDizJCzmylRtu6Ie7EY6ELaD8eMSDWuJdrURyABlUu6OsaDPoj
XEqh3LJJdbenpi03HnoNVb3ccM1J2fCdaT698jypbTWsatr/sl58w9aFs7RwU/Tu
8CA8qeZ8fGDUaw24SlsRJH4BALH9X/rz7DY+oOHbGQMm1HQ+BqOISIXaqHJkgx2z
u/67dj1NeJWPPvWLaLHmllpng4IY4o8owzimsz+3mBySgsoguK6v5h6braFagih+
pZdF1JyRoInHOQpatZ/ivstZ6aq+UKG/ZpvEP5HZr9i1PiuoKGzHw0afPqPoYFTY
19rf5uNksw45m6NrFwYYVqwYq51Wfz08pP4+0IZRTEYgA95wQprMBCCv+OmS+KN1
FkBzHA3ffBy/qyUlEgKAQ78kz4vPn+Fth9mhHdbsDIEBOivN85uYT3500bpGYJCS
ZxtZxJrPLDwlNMEFktXmV6+Z3xk+2GkpchG97EnwBOirvuEo73K2kUHvRsmEks4Z
6XQBwtcZLu26VmNl+ZsPtbWTsY/JPSoeQqV9XoDPOpcazpiHeJMDFeUfUapA0ybM
E+Pmd/XkSqL0vLQK1HjDM6hIzTdCqW28+Gt1niRnqX+HbzEDSET3GVh1QOqEXGF0
jcPzapP8RpEy3uLl6ikjcHACk+p9P1xK4DfcnpZwb8mFxwLMLBVGGtuMF/YsJOjF
6sUKKduK3pHefkG4TU493GG/Dfn5cxHvY2ZK877nj0+nMHTdPhMd3lci6/Wz9zQm
cBYpK1IspPIeN8xbLuF4Ym8htWWuQOB2gzvWvIVDGDf73l/crJpURtvcAiqo/tPJ
PDO8BB1tGrl06d1C8GrXxGgpOcM4fOf7sYDUzUzxNUYdoncvRfCI/rJY7cein0vL
LmBgsqJ3xrSv5K6HiIqs8jcZJHEHpSL/jdos9msxg4FJk5KDxfPYfDLFblspuqvy
Wpc6A7p+umloEY8sOc/OEuT2HqPa4Oy9RJGfsV7PDKInRJpN6mqgLny/ypOcIUW1
ubSAfI3rAOETGDBzpRER2D+Nggd88a0mVg/HsVUTUHRd7sSrEQLn0KGYaLq9T2y2
gp6+yG9Bft6qvWF0IL+gG9XOXIYBznzGhbcVc887rA0WX+G9MWz3MLOpWos3e0QU
mg4O9aKYbgzNKB1NKi4d/0Fj9H34UPLevwgLbMI3DBHOjGqFJmSmHi5lBhHbDmWp
woU6XDFItdQy4AhutXe87ujs38drxTiZDV23oJFxVTkCvCqGOkPk7W0moDLQeqMi
vMOBSi9SlgreaEqjZVgWrNqILWny2eJTBh/6eX2K8c22M+1eNxyUQyD8Kkc/wY5e
JSFS6mAslPnM+RfJe4FRXdciY1sSmlG1LR0XuPgub0GkBOq4zgCN7hdVnt4YJiRT
kBNSFZkDv0GSZMa8/Hc7R7moW36MoHRdQuPVve4dXRewxzvI6YnjHHv3+GJjEAkN
1YM2tY4L/u48EVU7mSCpgjxXCIBQF+kZOCOGJIOEyxnQb8gXsy5Q3IfbCvuJWm0g
O7yyMxpTjPpXqTiObH/mVUGrMD4BHOT5lLdE13LYSQCo4RDLLFZm4n9WY5zFLxlQ
ow167sMzCqYob7gGI4dO1G5pKJ9OXxB9sE/3v0Vfms+AMPMn1ciES1klAf7vvxyH
x7viAl70OuW7gOsZY7DTtEAFJNZcj6lIcgPjznZIu8NsIC0uTLjRk5m7+IoaB+JS
vK1VhDY38hbI5mHn2Vn5a7yIlOsDQmnyq9OmKnmOc5mRQCQKx1kOQwW0+LzsKlF/
+yBXCYz3XBbO/yre9vlE0Iq50mscMCCHDIoKVmgJfwhayiLJ7QlAjpEthe/c7KI6
9bxNB/ib4NH+dXvOBn5Ky+cTTrYkMgIFrLG13YRCMvYWKZgmSTIh05XFft7n55f1
ljHHlLr3Z6p8g3gBAlWoGJVr9nMu1ntunXZZFlEDaPPN6a/K58cCId+JUtOW+4cN
zAX9o/Kg5qa+VxbA0z9eY1CxAJ2h5LM3KR+5D1Go8i7tNmalNHa/a70qFZ5g2++B
hyzKPlD9coaqePZ3DFSgCeSDKAlAylNB9X1E77Aca9ynlvs4hHDxJ1TulkyEm/pL
LdpUxseUiUZ4595VNjiUxrZI+65PQ5IscGOOXf0wmM5hTBfNPehULJpdqWhh2wNo
RCRy55s66iKLXVtYsOZQZjfKPeyH1LJi/0Qwsmad/YbVQUni/LZT0qbfru9DXlE5
1lAwceDHyyqorQuOJQAftF9R3tWfOcYY/IKd9gCOO/up628t6WemlE2anhtlObju
+27KftT09MKy5w5aaNGWO0ZW65L/z+32XCP1ceB65sCaSPBvzjsXmHtwMz9ytadW
pnAoeN2fEYZqG7LxbwD62JZ5GlbZCFdI/mZugkY4WJaXx/hSsqlWcFCKLA7O9p19
KVr0FZg5i1vu8zina1BEvQxO33jNFuvNzwN7/qWH2Vvdywt/l4BXukYEB/M3HYSP
OGNJsBnLqnnWzuTSpvH/neZhovUc9mXmOa+sMJs6f2ii84K9+LKnq9J9hJwplWu8
fJRKM8EhAKfn1lPzjWLWh1ZzZDMFcY1KKVqQ2uFn9t3eib6CwVeg3Qz+tEqkuq4T
FNAfog68tYIuJRzheubbtO1l+evxXVENRiYqHCs84E1Br62HzzvzB+SsYYZ9zrVo
F4aCP4TB4z024L9nwCMcQsYbzbL52bkw+Hood1uoAXtPhO9zGibDV/bdY5Mhg802
4mK4HMioWK2gj3nrIzvWNVv8DK+u1dpwXsFav+/xWDmuZwQOPxWdFwwc6VI4FfHV
j7jny8HvRux4jJM9uv4R/X/SNHYgiXx8BVvVg2C9k9RVebtZ6kt8ebPfpRkXdTLF
J2qC57NcS4H+3MzOaxCVcnNxe+mWj6wOM0kqRl2GiapcbA4X6wI7rxihDCF5cP1O
aANMIglnjDJw0IWKtJ7chuxT+N2Lv7njWGsL5aNxk5KQhPtzGqudZuHuCApTVbUF
ST3X3z+NI2eVhIssRPaMEDm8Oh8WW/wfauzmATl0y/tCATMtqqjtFtm54bAFiSj3
9/2mUc8zPwYSkmaQUQVZuCh1DfdU+c76um9g+HX4nSKRVVN8LLiC7DiD9U2Jka3T
JwyFd6SidiMnGS4DSfcAp/ZlchafNLU+Q9oAcJydkNl+jKomqHIzlRIPa83B5cef
p0cxBHQQDJAjRnY4brLp/VutLI041+Dc9Zqz/GsfVsqd1TDY4TpnezSUbDjCvmv/
YOaPaIXbsS0QdcDFM4KbtHwKpd7x5etLzgBKZZd8n6q1xI3MSAsxgTtHqW1VhrP+
OIuCsUKPYkjx3wEJTglLAM7wsfKTXEl93YS8/GL22QKkfX+BDMfAMBbRVqyF3J77
LyDzeYpCJLL1smcrFbrLmCoazNAUP+roOvK4CNsBPxAivn+hWXBb5lNav5rWeZuv
03mWdpXiU4CMykWldtLLiRm32rfGb+2WUni30t6snpufTdhp/0FOFp9fvF22wIsb
J/nI2jfiHgusrh/AwjkunSlW+rrazH8fGeEzHkvYNJBCrcnFZJl+p7qwz0QYURX9
rBK9QjPDaSQDSgXvOmid0a3KWzJQdEgnpiR88rGNrQCpsDxzjkFB/11LXoXOhCw2
+6D7q3PY3bay+KLZp/B4oAgKhToIXibCUmu63oCgVYwmrp2ztoueep4rul2ILm6y
JYrJpfnFlx4NxSW0ACrOGQczTny50/zdwXzhrDwhFsh5nGdkqQEtpEUoqvSIk7I8
ldMaMpTyiNaOy1aa+91Jwlw6ilMGwkf1pFuuD1wfmBDtSsvTlFzzx987HMTOXPbU
E5Kq2VuaiQmmj5+nvOyOXpiNJS/6B0aDb6+I+BcjN8dvzi0ICf63U9vOb0RV7gyo
NPfW0akUHli60PZ00/Qt2Q8i4iOCNgYd2s3BID/Xn/6UDMhqAWzWDfFlYuLyk3Im
9dmC62H9rk57VuKqUvAAlgEqNnwO7ErM2liskFqS5YpIp2eGvBp32xgHRhJQ1WNB
5kJfsfR+1lk4hbyAcIZ1kdZfoO9dgPWlAQmcCp3CJhy2GLTUubNOho9IlgE1tzM3
C+S49IDftowNdGv38KFo0gU7IbL1sJWfHjYRhLoGeG06noPxjS/Wjp8AFyq0irCE
MehRyrgTWcw16xMHDBa5hxDioEa8JbHYLQGZ8SFIvKWe+Gs9kObLkuKfNJAw1bBj
XQ5VCgCSaxBJcQJmE8A31GX4jQTTVa3Od3MVlM/OEJ7+5ca6juLiXon1nhHjueqT
1TjZmcZB84v+GsEWFegX/pXdyxJvdGUtKQpe1FL6NMEgJ3IpdnC4T0MeOpavYpNo
/O5Ztv9xyohi0z/AkPoqUfqTFnwj5bj1RMY4M17u08gg+hiy7AdqjpvEvHr2gbi4
//lQ97CVOc8WLL3PWCxJr7yqDkfo1h1fw/OYgHr8yEGpVdwmqpd+E9bc9hM1pAYM
Eqaf4mONJCXtSG1uC9PG5iaLP+s/Iz1BFg5K+coSysfGm28LasUmT2QAgqBpUqKW
KFCJ6ksFNuDzEPRzVvy3GS/9jHKKvsA+s/bL+a495sU975qxbwQ3Y9SFqaynBlrL
4EBXyyhLs5KI7ccrfmk73R86bdQBE077ALabgKyGL1UZabga226Ws1pa47KY5cWW
dAdY0qtPJ6ejs7pA8CtyS4bpkbqag+bVjYlekDIjJ/vyz7uLCLYNsLeCi7Lbu8SC
3A/jPYQc1B+NBJt+ay6KhgFh8KrrPcCANArQIQPjA0O8s/ELn7Kk1JSZbqSpYgwg
Th1d0rOdCiAbt2q3s9VJRC42+kfswFr9nNot407h3Qge7rQ6Rbk1LJ4+nwX7noS8
VYHBMD5Ps/eFN4lZlznnm5he/pIRe22oYATqpaGBVaksYpoPnzFq5Pi9QtyqkYA6
rm/FKqstGnMk7/UoCsePi/DyQ/B53SsOdoV9vFE6LQl5tedAZu19zmc2kcWGTSuH
3jz62yU0eJOIiNb/xB5Q81UeXLZorILHyDRxp8a8mwVore45pvbV0TfI6SXOskbY
5fuLUCQ9FGor6gR1zb3tTLUH82zFbwdgJiVrcNCiSy1v1tl53SXYMyiroeZUyPmU
VVyLbmgVjlypDvkTm4FYZtF0XGbOtYUqHV2MNmaxKVeTVfj1+Z1NHHFbvRVVd9kY
Y7THJP3u1L8YMI5nR+L9iDI5pcDUENhzba2PUln98GTcIIRimNlRS4K/YaSRK+r1
Q4XyBm7yzCIqZuyfYGFRRNjFdu3CZd4QVQOMjUYk9AO6x50j3qtXfXCgWfdDIrsd
UVlu6Ga9gFTPZIdKyrLh5czO9fqi7mSGvwV016O7eXQh3Oyv0xfbZ9tpr0nP8Eo4
CSZceUzEdS62G2r9oy5fyQiRPgRuzNZVPAFMzIon1h2YLQLbIAueGr62NrxG0fxw
jZVTzaP96BakwmTr1tm3ER4p8Vozr3fwhEHq+M2lSNeCJwCTAMust89uEbEbWI0Q
+k7ZL38kGyn0+hPs9c20/Wc8iaJ3N8yxUl3a/DkUV7i4iHZZqTykVdGI3Iv0Y2WQ
dxid/cjmKGCnJT/zpFPm6BH8kPKHM7+ZiEC8q6OFaU+AjS0xIZKDhTJLicSNTi7U
h/7bptcUHcAQKSKubL5cuyJVYPnO2K1mhgzV6nsW5F8boFeBP0xx6p7fW8sANhlp
6LrexxTo8joy1JdFwgm/tIaqXpnzEb2PK/S6G03eiUq3/j0xdZDKodN0qKVuDxmS
uHFCjSCTUL1hr4OWEwAS1dLJDNW4voArsJi4POJee8Zj507vLDPBCT5+3oZXxy+4
BvDIMNqMD4SWCor5ampUTxPtXG3kPMgrWhBLwgeivS+wuHdIijiGx2Vx0uYkAyMJ
9D3o86YC9vrev2mrBcK9YBO+xJ2Fgpvb3Fn918HwO5ESJWzxNMJQyjcferjWD6ag
F8b+r660c48SG8Cz/PibjGDKg32U1wZk7f0uiTc7zsJb/mxULqSI0liI6AgZ0wUT
NQbhGK77R9A6zNkxuGs1EHbsk/k/V8DzwKCyBa9jk3wCHmxOlD3VJjyB0HM7OMTS
LlW+0JGW9ugWU4jaTYyV82cLIae5UZwfdN1yJbJaYLi0rEUmxxV1HkbLSVY4H9Id
57vSQQyLN9HCT8+16Z36Bv7oqnaAn2+8O/OSZfKYLF3xubPOjNi7Me2rEZrA2Pyw
OGiW2N/4NR9o1UkN5SKgdVRWBBd7qvy6gtWNFFPYx3Y+No4sIBpZoF87FC76VmTE
QWThUJkXJrGE2D+S1UAYRWfqF69m4iUQuUPWdIOUv0D2Fk0wJbjT0jR5T/XlhNtn
yMS7bD+MrS0bSG6H+BUlOQd9/LvvMCdY/3XGP5Os2AUzGKvsVfJY5WreBm4C6xBw
96NDNcs4SxaaBOHy+nTNQ6XoO7xZPdTDGy9EzfylEkIHjUlSzEeuACOpKq2ZIzZ0
xIVfzMUc67R13A7A49oZ9P9wu5BdWKu4hiGFEEWQKs26+F+I7Fx27t8oyHnhzOL+
Q4mncaBLIA+fHHOEkH6qRX4lfRbMHOsH5CmPM56Koo5sxidiISQW82dDI/PoNipf
Dy6WnYPeFIWRgCpylsyfNsZ4/KNW4gC+q60CMaXsQVCeRoLhT8pgHDAG2A34isdV
0lBvu+PCc2rGqPd9Hc7vBMTk9cWmn5DXsPd063+s91eDofWueEt41ZTw5lVGiPN2
JgMtGdjMGjJfjz/OXBHGVMMS1FyZPqy/Wr3FEYh1tP0MQMN3sVbQ+gl/A5GpsfA3
hcO5NP7ofcVTNPoCfViHBv6/L8T8wCTl1gK1EM+qsZb7TE/KLT9Tfome+zVaZSGU
qJAveQHFxqHY46Zy2e5C1hGlJx3k24BJmMrQxRW8+/hTJPfb5g2S1poR9bFFctqY
IhN8hXD2csLZbifKd+nKbFdEjzhVSdBqnNi9XlisDyoWauAdbULppwRtRDQgaUxY
n87NRTrbrJObNODvg2FbBEXcv9GqN2m9Cv7TyvdtMMZw+xu8cjdCjkC304JMpSCa
/PQJjvAA406HVWlwnAw6AL+i0a/McqlTI14+3IrabZcAh6crrtoHPL90ARTcEpXi
Ag/wqHPnM1nasepXOgMv1Ztnm3/Fl0bNItVz2EdrQ//CRN7RaHxRh2w4sQdcc6mK
QSa2wLrQnkRcwLmIrJcRwgXn2636k4Iu9PNmJpHnjU22D/xiOIiomjaSoSNdUg6w
1/rAwXfMSAMUKvFPpedFTEu5Yo6AHImFLM1jVBorFpvDEZ/dNMdT26FwZiEF52bA
LrOqd0DoBRSlEpBtce2Uwxh6iJ7inrhLOdl90G37CT3SUi9ZnIxrBv0AC2XHj80n
Fpo+tSgpHLp19AlSgG/NlPvKZay/IFT0qZULm7zHAHnHGeDQDOQmGy/1hgOMquSr
M7WfXbjGYavZ8JKfIWezAXJIJOJSaO8KwaaF3+Rg0GPVuUYfslJScXEFXpbk0RYO
peHwNFjmu5rc4CO1omOJLJx3xESgeFpGDy+L7EdzNz7vmi1HLzMGsaowZSE+pFWe
P/VXTp22NqPBV5Ux48KsmGlLSYxniH6173Lj8GCTPElKw356i7UY2lmAWl1nZD8s
VFqworT32hLgwC5rXQGd8E4GvVx/xHytbadg8FM1ErsFQzY90fpD84JLOHQ9H5Pv
w5LmR0KDXpJok2mjvWB0OxWhwxrnC957xhXH53B93E0Ryz7xvALTnKCUv5/h/Byp
3dy6wLkQNTd7PHKLL7VHomFcVklY6sUhNGxhuEvBg1Cn4eVjb1lvf/TpslyQK1+O
X+ifufBGUnIrFk5BdSiDTMb9uCrePb2PeoYIy3HQ4w6C6Ioq4Twk+sWlVT0oMHhK
44nAmJ0wHxRgNqo9SSDYJMCJUQ3djJ3MYcebBmxr9nHmJoqTkCeJi5pDCBsiSpCU
mFuF7BR5Ei3m85a7v7VGOQ8cwuRUlSJyBpbHRynVpyiCO+AKgKLOaQht+7KKIFHJ
doEK6J0WyMG9jUJQAd0sXTNSu4cB4EN/MwTuQ3p96F64Z3JFcYQ9+TnXL9mYtFZP
cTnaQog++TQv2gO4Pcko1asbPVtJ85AE2IdJ1c45x8VgbzIiVUr8Ldj/MCjPlaCg
4yP0Bf8UxgKFKswfblyjoqLMfg4+8QQhgJIHpYOtpbvMn1wczlfl2E8/Pijit7lx
h1jFktoh0Ki9D41mlnGpSr3Bvp7C9+YQbzzECLmak23Lhj6wLxQ78YFT4reWICbh
dhvDnOYElhsR2ZvR3Tc6ubuwlfdhjqyRNKQaZh25YTsVw88hX7iSe2Q8JXUWkt0P
ZaZeA/NTw7iafF8zrTWRmaujLxwN5PcxgA59Lp26mzEXaP6iHbqUKS0PhaAz1TRI
VV2KzLdAmL2WMFd59/BRTHlDf92qNVwmBbDq9KA2Gw1fKf9eLeDPYLgpDjkRP3du
W2PyqyDsZribrfHWU7sea9hmbNVxUIq0WMfG6V2rHgqEF82I5ujOh95rf4J0Zi0e
3EFqp1Kq0Bu8DriCDC3ZWKFC01Yp6+VZV9dGrVSaY5vOFpMoH3xtiJkYdw87bRUQ
KivRG0FNgfYkNrvyx7L/t9Rb7x6GONvNDVfLuEATdSRtlc4t4pnCLWDs+N2AnwZY
0UKJShBuSc+4vYMfbURGsjua3lbCxPhOLKZLbNH3BzD+mEVGi1G3j8o8VYdrCQ+O
z2AMSBxXSAQrb2hLXqquBzp2aFA+Pt1j2pvZ69BBxsSUWyqV27vtFO+i8DpUg/Zd
hcJ04u2v/889Q2DB15htXhYxEQdrlfZ8psYD2tB31DmdwXFR3fE5jWITT9lHvxzu
n0St+7uOQhrecXuBsOrQme64L2f6WZBsY95+wzy7vTtem+Ho7rQHuwc5BoYiTIRE
OZn9FX7cRc3zIqXMy6Fifd7GvN76G3AUEisv5F+vdLlZU+8zGd1qOUqtJg7///WF
90C83nj4puNkOO8rrO6xxnvAguxUDmZLkmtm9c/jeiHPsZL609/r3Nhz7GPqMIrl
ySFkPNqVsqffuMRBt6CCNDBwEX4fyRZVEnN9mz5FR++1ukiqR+B78HHYKpf04OWx
h+dMK/bTlOv2mBTXtTXgZYpZPTO+6weVUj1Qtyf8Y0R8QQbCz9xvyVK7QpvWRRSI
eTnNR4ZPU2Uu6gMSmAAwgVKUzR4u8CAZ+5MGo1TNf9joe1SuwNs04LnWqs/5/uEL
4gx8lTH+VGp5sK/aB1R2adPg67NYhWdXfui6lnwGVPTy5FgJ99w6r3TmyLJI+laK
ya7RAMNe3wSOyUVedVLqYfaSKN5Dj81q+/8HWnPOK7RtUYwptbUO8rX1ao/apup4
oOG3iCNDgAg5g+ffTcx1BSvxdKtnigHUxDFUhnSnefyNW9L2lLIGSpyFgh3qWHWf
uuXIKoJjq4VjPYb52UcqIoiNzOdi1oXzCNycEfYxGUc6ZcFdrsd/jXcDWK3tt1cd
UB1XoM/5m0v93vqV0cwPC05JdhZieF4NlAUef/vT3qTP+ZsyhnegOqeL4SlNKhDl
iJvoc6U7n8VGdw2DGcz2VfoRz/q4e4FtPFergyYuXmYLnoYyzN6Z22izpsAVE2em
qrS28vsdXYv2LcRgxlk5ySrOOAMzqW53NYvJpSk5EWBPIpWEWZ06ruY0qw/ZA07M
r4JS1pmMYj2rRJE9wOjNgdysHJZiQ7gbPGAnuT/vBU4j8Fb4l9vRUbNL7WVnYOSF
GtF/Q8CqyeUKFXku2OfbRGsKxtB5U36lhvAMeckxCwDFCSpOQ/yXM2VW5YjKemD2
4eCpFNY+UBIu5KCAg/BjA70euKwom5E+7x11/iEtAdQk2p8aMwUMi+mr2zfWglJh
QH1sLsaqDs5AwzO5H7zQ7dRY1PCEr2MSTYYQYO0elz8bPwRSxvSYwa4onSCIsrSx
9QpfIBUY7w9HSzRQ4mvo+MvJRG82DftQTu6hKJw+WVg8v2zrtCDGyr7CWXF+PJCo
Mf2vF35Fzr6FR0yLrWH7g4cxlNlRQuUPg45eH1CPGgJwgS+u6osDWRdRpNb0QdSp
SEV4YJWZSbEs3ChHmjEY5WvB2ZSWVKBphB+YCkz5NjB0T3g6cqzp3PBO7hXewgCw
PzgzNUcyqmwhaAmLM9WNTPMjTxHBgX29l+szMiUCv9xfWToEDb79q2Im8is/w30G
52SKx6ThpHrKlNNjMkH90JoPRcVnxTkzaKyYjza2Zs+srC0jdF2TH8G4LtTHBWbD
z8vQzjMr7uJ2katO7sFlcri82h6lFrVFZ4TBQx6PdMhVu0vCRqnwdivhoForGLdc
gnFN/+U+RCdVG0YC7q8FQfIaembTeAE2WNUjPNuN1LLt3xIMSJgRz3Or9BRHEIh9
IJwlhO2GcD66bPgrbizLQcLfVHG98Kwt6ytFYgcSOlewknXilv8wAXokHX+iAM7n
Rf0zMcngqY8N77CCKvnV0jawPm1V3lJi+6bRAqimqmEFjOVQABMNhlvt6Gd4U/7r
j8/ATp0O7euMm+lYa7/Jav77bEyy+E2K+8NdJ9pHZwyUeOkFW2qolq8fyVJnN16N
8fJDuZQvZ7lpuY5f4dd8Iu8PWX7rRWjTKXXHUy3zCg9e8XJJmUgnDz8vI3O7mcru
G2Z6G3BB2QVq+oUiGi8tMDl7k6D/P4ZUNhn7M2FvUhtSywV+Kh343j8GYsgh+h9F
`protect END_PROTECTED

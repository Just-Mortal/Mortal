`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RgWWKH6qGN74/exq+iPaZdNA4F/EacAimoUVLe6nK48gLhqbbSW22P6Qio933e2
4NgxNI1UT71zuCnrWURxMcAsCz0VGukcLxE7nJllzLpU1K49yMUa4nCJVAJagLpY
ZaaQFlLaZW4XNyxQhGFTzWST98mRmkj/LKm1zUJ9+7g/O1bvW0F2vLDVG6Y/MH9p
Y3Z3Z75BeuJY7WkLHxaDEsQgHDQ+M2k8plj8eqtr3g516YYhTAALBYHGMktQJETO
zwYHmc6Sfqnb9E/PQXSgZ750MVh1FZ/ZUyiM9WNTfnD7bZxKiLxhhMvX59VaE22n
hYqNsjK/ML4vTZDYqUhJ5KRMpjDoXKJdPW5z2crFhsWLL0agPwNMOORXgVrhxnIC
7aw332aqaf6LY5mJajie++ceXzp4tcdzUJR9BJ9YimYkcnUBuzky99r0+l7xPlvl
eNA/IIWZil6wOWSDOuKy9mjmXuSRyX6YfI3XpnjNzPvmUqLMlHE9e8kcpI7LgsKy
hCW3iOmJworeSD8u70YfcgqwWTrFI6VmF5AIdA50g04nfNSovKytMsdOYiWVb1TX
SMaGav4vA2ZWwzVIt/UKauwgRAzuon49+s2hDxwzfQ5OkbFAq57QhDATEGLc1jFz
S9fr6PxTmfERIOGTz9+QPkKiZWTI8lcPsz7SFFGpjSZmq84yZrNR/9ew5usw6+hj
IfrTVQFh5ue9q0UAbBDBImGwUD3CPPaillxqNSJhQtjdYJmxFva7dVQ4YIiaKzF9
yaxaFPfRcED7jvTZJljTVrPoxVUP1Fhzc9olb8zQBG06QGXiMYmiV7iF3HyeaBlL
TYwAKc/SYhepwfadDpQd9yR2PQYSYPi+OUubIEI/8TdxvCAdo76wTUDZtqqgOu79
O5MCyjqpciZR1tbPYCNEQvB6eUK9+M2z7P77eTKJcCDB0Fw4a2CLbuNCWYHeTQbE
urWSFuZB21OD5zED3KFwrDZozehPH2BHWjEQGmgABm52oGWouZGLBYNZn71p3LpK
nAUbs9EAMMHL1BEcD3flDAcTKsjK7d9NbgjncgoOGdS+ZLhDmU/mx1VGqxmRulC9
VANusAZNfEi565qWegpOZYbnk2YWxFo78ot+0npfQorLFp1ePqv4p3QrF5VbN2gV
ZcnY41S7Mg58QEpw1XLEEnT1f0NjxVLQC8sKG6SED6UkUcJSpA+jzwZg/Pj662GZ
DYjespDINDV/See484fWGsGqn9xNHCYDeS8OJn/+SoHLBKCgXCjzUP8FEYh3j5Pu
UPBpiYNXCCXpD2tte9jD7B9NY+z3+y3RaYB1dFjPi6D76L0oF8/Ch5n7uYYlxnp3
BR+6cYmHZ4rRtBZcweUzoN7ehxXzC+9PzwfpfAyZ58Wg5/tyh7zGVuHpgdYlYwCE
DYCz4z4GjtJKPZ/H0Sz0jMV2E9cFxg/o9BpiNObyZlFZ16PylZSLDRPE1YVhc+EU
tcb6Mut5hekdPL9Sz/cMQ0lwEs0+yikKs0Zw/2sKDpeRfF4XSZmIbnh/RKKozHF3
1/doyRSBUbLOvR54CACPwne69gVhkN0oc6g/R+mw6ROk/cHwvtYNCJDHcJPspHQV
gPGcUlxK51jUpufANzYW9GGKDr6am3JChth2HhUDCp04lJ126AGjeAFbXkSPeQFs
hzPJK5r1Hnfs9hSy0EKiBgwnaTPZaT5tZbiE/9uXY3jRFbTMnSjO9jr7A8VXGjgv
YUSsYuMnbQVKbJ/98hlI2xhF35vOzsRvoMq/JLGnBpp3eI3vY8CZXf4fRsNp8O+x
34B+kem+me20rcxC1VOqZeG2udvvDsgzD3Eg/hEMxNvfDt5S+yOd5FqnmCmgEI5D
yQS++1R77vgzYz85CzmsUtJtfg6c7WiicDQlnlKNatB7s25mnDK3+NAsMlSFojQd
TiSu6lp9fSeS00IgDVFgj+Y824SBtaIWNI4eHn8fdHm28fiaR1O/VYUVk27myaHV
zmQ5p8RVs2H8R7gpgMAe3wjMq1+a/HasFqAIUmjOub1mps4xX2vUp20Ig+qjA/2P
0Ko5adbNnTGFnRMcUw312HMjOdJlKx3SI4g58K/hLKgljAFrgQhZR/ka8V1LdW3u
jAtDacgYLaAnnxKulWSc+2D1bnHtIIJps6esoH1HwHS7SywK4YnPtpQRBhNGwZVF
g6+BgsEKfCidjYnIxTGimDUf56oe+yjSIGGj8pR2slYZy3mKuJljwjKfJwqhIDIQ
OzaD8YOPhB6DenIIoitaxUV1ETHGKQFDDfwB5ti6GGk7vzLZx0iDPmcPZdD1fpjf
LwBnDxn0wUwHgDw3ryf93fftJCg83r/G3N1qzJsiye5vR1REzrLjPD4/QHR/JdbK
A7M9GAZsBdGQJRQczqIFbJUxNWWM3pzMkAtjKKwhry2l7f6dOXr8Z47GQh5FMlqj
MEs8ZMSrtYF5FKsTHgyP6moqO28Xr8sp5SYqLVHvXpD/ZDGRIKzn9yi5QQP3KICQ
ocMDTANKZMgBzhezSKiq/0J9TFvqUBwm5Jk7rJwiJn2xxvJzWudscjG1kTmnDwvs
hNy8dwrVjX5Q9xAEhlvOC8Y+gkvfMOvd2y9ijrCIakKb118CtWa7JwuZNM2KuZAA
SWhjbwh9AdmXcbGjXG7Xzsdzwcc/Bnmfrfkx22HP9slIF5FIhaJosKQJhIACCHcZ
vAjgBAQXocBDS0fTQxXkF7+fQdVhaC9x6y+eIF7DwIfOPgzlMyzOxQ9nnM9ct95e
WzuVArJPhHlgys/sIW2KFZePaz86XG0zMxPo3yBsDta/x3P7a1DuGeQN0hgQOEbh
eJFBup2JKqX8jozsaj5O5kZ3yKZPzlpzPazQNVI8cXcAWTH1GU6Tp8CcQiLshhhb
mpjLUufjNpu2J895H8DaOPXI1YdHqhk0UsQ4dKMOi3qhCb+vT6zsMgne3aTud4Pz
Z2h6CHMoxlAvPF/3TKM6/W4EzlMy8OqB0UUZErLudvz2nRSrs+GRkO5kOSp/2n44
eLDaUg500SjyZi1/gqjLcwvXQvADEA0T2reaICWVS4RU7n+pvUHTwOEkGSfXy40s
TX48W49K2PkhA4VMG/b9t4AZZVc/YA8TzTjAKPsJWygyr4cnY6uLw7dpFfFEzh1R
aAkmDLbFJgyE/xRDEMhcKzu95uYhfQU2B+CL+zueoU/fECii2JUgB1P/+jeHqWTj
+FlthnxHZ0nkg77JnE4+r1To1V8iDZNfl4hHZcp3h/wkuaWSs2I2W19EsAg4tTvj
9W5panBksuLVwFIragGoy+9NY4bPOxOQFFKUH2ytWDMXrVjkVUfJVBpjJ6kN/JeE
CZC9B5R4arNLToulL7Z8Eea6BaEUlJ12A89IQa5u2DVF1Vc4wRcsB3F+VVgLhVYM
+LvAFHnrOdMqAucopUhwskrEgQjitq5DeWws2lAk+1x4iGWDcw0TdW7NBRM7eZpH
Tflw5ZW6ECVfIub1Apgz+dYuBpSrNSd25aAcpiN7eTAoNOauo9ZDoappPxQc4jb5
evlPDvLXRZfja6Nqg5YmrDH3Nr/Mu9O/PwoKP2W0GdetE/4RIH0mLdluGf1buxg5
GP2c3K6unBSjlFskZI+wxTMvGCOrJLjBBVqZEOjGzHnBfNxyGt/7WhiDvjABGHcH
likPqaKYSJFDGPApRN4+kNdKDAa/vdRiTkDdNoRdk0hGYFfyRNnpeXP0ghfBV9A9
5w4qpyKt6aC6kri9kwyYq4P9sw/fd2Hc6QAvdWg3olRukhm3CR6j7wKzaO4h3Tk/
cGHv1qbVzP9L+MRQldZiB4eMEryaOeo64NHSGFAp/n9HV8JtgV+6Hk+DKnxvuDCI
IL8LYejlOg+VC0AZ3PWHuwQIIsQf7IHNyFaGthGnfWiAKGh7krVFCnIXTPGp14EL
poq7D4cfPCsdsCHOOAZhq9tx/OHsVutKjjGUkBOiKYKYr4LEvn0tneYKZQ1mPXj6
9wN6T+ZpDswD7NA/bAdGehiLptaHwRjQbs/H81b/pU9wyNE7r9CEtENspODQELRc
sWpgNcXQzc73fXf1xOSD9nonCRmLlmtqwSfda3CBunQxNnSfASwJC0u9uPL/cIfV
FeGxGSitDGj0XZit+I8YScsRf/1jd8MJzjCTFbSgKU6orb97whuJFTEWCAfCuhfq
sHIADv1bFXTIAUjZKLIx2s8rLs86zGqkjlp1Pr7oLWm376RKvEKU2UxYKEE3AejU
MPVuu/Neq2eD3ERNesvVNohPkl10x5F+3SAyZfC5ni/OnRo3XyWKQwI2hyMp2MTe
a2zWbIDr1JV6IgjT3qCkJUZ2fITGESBoLJZ8IK7hLJ9GckbGfnAPOVl+5trB87mr
zv/IWlR21qkVUGp2ByAddxfDZ03IJJJoNvZAKD5m93+qGtzpHzxus2fdSpjq0Kq4
j/24JS6xoAXJWbxt5GQreKYT5Fw++IU3wR1JQEKWXjHXjj59aOqPXRsxVa0FhMII
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/C+/QCaxlkg+lVL/LEwmAdeoGqduqa/uE+7k/1X+YSsH2YpD7LwWB4HSL0mc+MHJ
4KaJe48rwrzU8S9OvmHe6F+12Q2jUxc4IBuPGS/6ryf47J9NzfTNfgcedgVTrkhA
4GhjhCwNLDeiRKx66SIHTyrEKPz0K09pDrFTm2RC3eOP0sfapVrNbyZNa8koCCnx
XdN8+Al9t+14JqmTB4z5AT1SjJVFP4QgmW2+fVn12b/eP/ECb206BGyn7+JY852y
BNH9MJgcOvciCFAO17LPhdcdlczGkwMyECTdWJzeXNE13V5u5ou3AKnK2QiLLBTW
G+pOiRuO9Hmg0iW/xmdUgpfb2bXZ9XxWdvNY8vks4nToz3EOm1C6/GXz8yfYgTI6
MWKHjLZ+Qvc6FsIyfMTsXF+hsorpQkFn6ZE7Pp9KmzkWuY0lZcIpvVMrSio7cRkO
Dv4L1uog6BFGPIo54aMd+EwkejQlVgKbHjBUyolrQ8TQyh0SvUQmdpM10aX4Gabx
D2TeWzIdGhcMKDNmXktO0Zpw+yaYWUyx6dYb2hL5C/BJREXL780xY+dcy9nbw0IN
KF+naLVhecEfoFWpKMYBYC46uBoaagZTxmU5bxhHGgkRbpiZo9sKYAwWGmq/1kc+
rJ58UFoXvT4vvuBgQbRlksKZwayXy8LvTA5/5gPQQuVLVmp/cVZJVhctdzGey+49
ED1g8y7BjCTzha3GKbDcz8tehUYcyEseQ/lsg2ChyerhsS3RebbI4ogMm9xtsrW8
8utE4N0rwx+47CdIIc+Ew0UVjS0A9apXZqM4u+EIvTYMXTlxGrRH/8V7XjCUK97v
cQjq+pShgIbaX4ftAfZ6gKJ4hv5Xy33PBAPG4SvAnAyrMkZYE59SbZ5ggTRznZDn
qFXK20R8RQUOwGhEKHlQe4jHUkjX3lLo/D5Vt2uKc0OSGK8x+h2HF0AzXfPcI8+n
vsaD5DLjfW++0SFJbUfNyPeZF+o+x6KUE/URAu0/q+GY506hCh7Gxt0zIb9lU//c
AaIB7iri+s2yeJEV7trCKj5t6KHLjydWbvvx56ro1zy88FmuD2ULG+0V51Iu0ZCW
OoHtaCPYxPvWqHzrFLkRgDc6KutpMLGh9d+I4ZGWtugNpdenIDDcBvK/Bv2OhPUr
NhjwQyi1IMH3MobW69+DwU59TQevM7ACpmfU7Caj08/DvwCWHuA8Vreai31wZDfo
UNLr9t5XXkxLk1s5AyEVCy5avv4yInWvfts0MEa1WE0k8dsVfXyrr/thozDKlxD/
XQRgH0vextGCZrno3cxB7d7YP6G7bH4TKaiq/nNA4tONcWgtYpgJQli0rOeLD6XL
PIyDHSwviXZ6wEK8rjgHfz9Hd5/iMMAEA4ZGh5GNz4KeXszyA/sO3EVWGBxasu17
WvMjtrzGz8hBHmAx950k7jp7ucGxYwaxkqb4KbPTl3cTqXrPwu7ww1OYXjLA5RZ/
KQxWv3OoDvqrsiEctRuQhCQQtGc3Seu3mdqBikBynbRBl0p9erwVAy2a+er+5rYx
kaVizwqHiQLJg/NMmzFimIJXKOmyf0qCzp9uXlFZ4ptbmlnafdKK0COf0k9Mtzgt
e9CKzCQDtya1kPZJT2wPTVvGnLhbBtizlblUKUoPIO3acpwfOmbBTOBfkKsczfAs
PrM5fIRdLfFaOZs/RqIfSOKK4TMGvb8gpIsd0zSViFcg8GasD+87CQn5m+aSuLD9
0+ED5ucUhhgx6ta2z1pAqE+LFlwGqxXftPJPWlIGmDJGFJeZPNl/aEva8d+Th7Zv
FaEWsc+EE+znOYBEynWlOgrPeeQL6WIEuNMxD7UogCUJR3fAjj+oWXhG+VTmdSVO
DNz/psGThcqMH79+8Xk00YK01EgE4vk/EFLSbcuAB/PRUS72VyyAmxk+X9p/C+RA
7tM+9eYpGKxrMfX7YgTVc9tQnvATlcxsuRJdes7ckdiz9DvevxBwMp0zFGnJ/nEm
aLLfIAqT0Z58bIrGhU44CJE8bXZzr+OhOpubNjciehO9U3eiw4PJ9Dab+CeK4jk9
0+9BKpiLQU+e4zAHOQBTDkKs02RfTxfcU9oS9epr5M+Grlt9gjQ5xAbzROudlVof
oxjTsk0xjczxq8F1pgq963m0ImniB23poTfCfJMaOcZDHmzzeh6cgrz2RYm8asj3
m+zsmecPd8Cq7zw+ZqFJ3vGN7RcCXZgkpOfqlF4ks+9nMwCkKGt7eI9a3rAiy2rW
YbeNwX6/TdLMIupcIQHp69UKKQU9IvQ1rWoVdUogkSDJZwBGVdGCfioVRbmbhFI1
ks9QiSIybzTI9ZzjQFCJi2+aB6wZEbUl85TkFREkydCPqa78GN0hl0RDZ8nj65ke
btEmls/MgzcXJWC4tz9Ya3EW+KjnOd1TmTDA4jg6QuNeTfkcbjR1tuRjjghQh/az
/mPJDa21w1pnegjt3Za1/YPDWPv/qQH9/hOOdGuZlL8C8l1AV2DaozsAHUozOzCN
tekoY0TbS5/Hof7LruuFeE6hHXtYLPqRFSyno0q2MS7fvLQ9MlO5OiZj6R4KMf75
rbyyIJNBt76JimVFSEDhJzKEUmZNu+pRMKWpbjz1UAFfX5QMUPoPznO0mC0qW2Kj
Msf49METJIvsffh+mkebbqntNubTgI6q9KDtmi+XpuWrQpZZVWE2V6/tF9bPV/61
OjCyiUEWNwYVCbAwYC0dBls4dzmtnuwmKd/IUKIFI1lT+lt0ZzHGw5wN/8ic4Zlo
D6SgNpfsRUs4FF0/VldwcBfenKIE8kwk+3GFr7IKx+aVz58k91f9auh0mtIzVKjp
oxFcuXxsstWI7e5Ag4HVamxU/n5euSOYATrW5RFYzNcQzk66llvcaEoXKGp5i1LH
HAoPnCrxgG3B5AlnO6nyiOFOGtQuW68AE0HpEFonMmXt6AKyc2fHsOFbdCnItbxe
OHvhgnO6Hpv3Oi9MqC39KLusEuLE8NAW12A3RRbKjgGLqF2gWeP/2hBV17YCl6s8
p2zgEZvnQS3F8ZC9/MX9r0Rh/ZTPJ5Hmlk4bfBJMaSRA27MRezCnbA+S2BkIidki
V4zXdkOiZsMfxyPla9SO0nsntdZxY51X/IK2I5E1vurT6ROTtnFTvJLqydHZpQTb
I8cv5ADqThxMhubCaA7AKbmoUq71vKGizidN3Kof8FByYK7Y75t8xAl1cGRlee8T
1Ka+VZEq/AodxPqJyOkuIZtm2SGSb90QfOhExihhbd5cb5tWqIP/5ADKGvfAQWTH
VVCXKHXfnqlhnJVoAMueNCFb/dColhmJuJQRTEp/UXykAIa222kr5KJraT61mvtU
4eQWMVJhvcqm2lEKJEtB2pLbWIWNFTVmf/GwgBfI2IAn+rxaWSX8dsb95RfbI9N1
tmX+yhWjBl1gMv4/3cyC24nGWFzEIMW9CE3QBy59nHMTKxBzhoUnE3TP3G/RG0n7
y8sWOrrxm9y87ut4S8ajwUAx2HRJL59RbZ6W80ZOa4uI6j4f2kIHzqoW547OlVej
`protect END_PROTECTED

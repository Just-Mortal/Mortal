`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3TbZOYlzg9pRezjsxoZtYz7mvqu4A33WopaoqB7OoUd4zdWoXBxWnQL0k7g3YgO
I0Slyku+Y+9e+prCaZu1rr5fiXGLWQUK8g3dC/oouNFvgv3B069/wL/GQbkH4mN0
OT+FtZ2tC0XmHTO2ewHyj9Fy58GYjguw4Cmt5gAA/VnQKyuQI4GR1VPvHVBlomEg
QT55ALOhtjaw9CaEIQxojTNU1QqIpSP2MoQkC3Sv+Bzf3NS+60mJzQpFrVwvw//u
iJiFLaAdwqIrx8PuRFrz0BibhP8t80JlOBo+Phpl74DNNR/6kGj6xEZBS7OEV33F
kTc9EHxXzT1Fu/fs1QH64Q6YX0Nvl0MyHUXvxtFKkCM4CIUppOPJRQl58pLs5GSu
MMvoMDcH/7ZjARFSM4RfmLsau4mwBUsvFtnLCJyfcpIcSBn4myvlu50h08ewjVNA
WpFpPWOn7dt4RM6O01xSuiWC9tksxIE3p96fNPMopM39ZKvVWi5Gp5trTzgQCixp
cjm1/xSRS+L+1vFeEgQ/qv8R304U1ttLg27SdtR/YD0Ob6QXrMM3dr55vWzLmPtc
jf4b/zbzzyWq7y1x4jwiTDUs2h5pAGlEOUZkhicC07SnaQAR5ghSJKIKRqnJWP+/
8NUbCNR/JoGI99mQyfc2QXFum0jr5+XwS++V7sei55OaidL+ehbrpPiE3zNX5GnS
7yElrz+y5ZzKoun6oiU7/pkk4Bhjb7iubGsZ6U7otOwSJzzln1gbUbokzctlzlCm
4e2pZzOUuv8zi1tThBU3NAfHo2d61nqWsgZMZcEQ08QwCg3WnGBVCFfHBBr3/nRP
Qb7A0687A6D38u4Id9+NYVf6CdBoO6KIvzzbjrbSZvB3iLZ/12zrXp+vsEzHyjb3
FZsBZgQ+MhJPqZpv1Xj/eRjvL6Yy0KnOYULFgHCM4ZbHmPLFx7cCVd6sw3Ym4d0M
XthC5+VJOIB284QleiJZYzAFuleR8RdkTrC0cJ6bfWUo9dYnU6hljndUl2oJj1Gu
zgFcYLiH43tofJxSD0ma5JiBj+xgGx2Heo+gNDQqZ5TYdDn1ACbr2YQ8VaNysl9/
MNQRGmhwHa/OoiDVmy2Rd7WiVsCJiLQWbpxXJu+9vVTkW2XoVzyPBJY8lZPufI1U
hRtrQlpxCgJZ04EgPEHQD4ZIsvhasDy//TI2clCOOWWP7JaHIS46rJU1O/1oTrPM
1Aokj6+2Wjxf5/ZZRV/28byCgoXInxlN1vw6n/lqacAMQer0s7X+tmroWC3aNuTZ
RuwV+D8p9p9BmWFDy58FUfSxs6bhn9YXEmjgM+d1RL7QRVLhBQnqcecsmsWNWp4/
7u9E09S6VnV/Px8PSxCDLyIafKNnrLdWZZSCSXMvSKQfkeSPzO9ZkzbihXi+Vx2P
be1UmF4TjvXJC/zDikPu/QXF8zerR/CWV3O2lvJkieeJ/C/LVW8ssPJFjOP8hF59
lLYRJ1UiLdHElFIKOaFa04icBT+ioT4KgpW9reJ0SJgoXkMV5WWwG65tfZw47BgO
lcYrU1i7sh5kze+WU7PrjiWjcNF59NCYIWS+EkuJ8g7wf3W+w2gS8t+Iax+99LB0
7PRVhpXAKCzYoiKe0r8f1eij0z1kVxOlrA83X61YJzKUAKq9gAEB8v9wPQW5Ba4r
p55HMp6AqYbcFrzSXi677juyq/iOiXnxF7YqxgXA40yTfkwSU6pc8jAWJZwKiBhn
tzaxsoYL69744faLwLBgCmVNi6wKeqtaJPMblY8TLEfn8lfBG/bQvlW4yd6m8nY3
112Gulq9T8aPoQDmKa0/h+LjX0BY12P+JRbMzW8gzC6SuZ5uWGBegk642Pj93I4S
nxL8t4BuJEHURzH5pMJU+28EcTMtH952oL+HIoRYHWMaAF9/6WmgWppYtlxq+WA4
o2yeRkDjR73A810nBREzspCazyn7ksmaHlI1wNV8HyS2wEIUz4krqQXpDQIH0UAt
DnXxoGW9/Wl858DQLRZr1feEeyzhepgLhZMcQ49OkZsI3gsZfubZMJjgJIBuTIXI
FzwWC/bsene109rdzEoXP45SaTaBbDLtEFzScEpQgAoERAQfcJboF1h2vqMcOoF3
xzonc0CxkMoXgDI7Quss9GEvn9iyuqdan+kk5m7OOhCglluNzzFhcXPZHTbpeH3Z
KBU+6nrGR9k1691bxXpEIU3+uefl3oXcOa+GJncWfykDjZIpXWDoFbQwf2F1Q72y
0NXkE7WblROpWTe++twFZUvlwCwIvFBe/U65MgUqa6JslsEh9x6aKVs6kOE9WU/8
lfRdIF/0iWmtJw4uX/RzWuzOp1Gq6EXk4eSGUZKzhAYT/a5t28Lgh+qNAMG56H1G
yRAHWGf/rT5P9b/PyvyEszVbasnIxeRnh9iBFlN7SE+rAcqdhiL+35fAnbq0+LX/
7ZqdGUV2nAVYblCKgD5nvl2ePBSF5i//1u1wPktf3Yh6z5x3YrWgq38K6/qouVl/
cYUaJcPwyQxf0IHeBTLlVleaJauG9uFc4RtUTn97qyJmI/bpjZN3ATpuP6/F0cKH
k35dxD31r0v6HJaYyGEwblP/6FFDyDytNhYuxpsArUfiaJnAgR3r93jcSxF/o1xj
eOKPZ0jYK3e+mFlQy51Y08Phwo4I8S/sywdv+WBdGqSWr5Ne17ngTcUZLhwnPgf1
CWlSM6rZ1RpiIcrZpoqPPF6Bml6SD7JduEWUKLoH5YGzb5vVOh4cF7bHRQF5MKAH
+VmK6Xjr+O08LoKDfCQCa4IRsMZRsmnx17vKaASeX76A2TZC7TWz6NYomE9OyC/g
88qxTGXEy2BbUrln0vAjpV2hcNfdFmzaqP1NCjkF7QLBKG3Iv913suwGeu+I8AIZ
o7YsfpoukALOeCOjjpIBdm7E/0BOVaL8J3iOQwUxC+Qrjvj70aqAMCptsXJ1ps5b
W+PaQbdCnzRijfGlgj+fLom5NBuhGLdd/QGxwiCm48T5x2TGa8d5CnUfveKgCcg+
NCrXIRdb3pKjRIOCcfkEBb5mIVeKbQh+rewAT2x7trAf4f2ZON9Jrqcfm2oVo8i0
8iGlyqbfhuCdYBZYR5MN0sqS+o5L+MdwI/P59JMAh20BhKIVIxlC+K2KQqq2UjML
Zn54/zvp114f9pwOjOhTeFs3OTweFvITuP5efCpWYN7/MIxE1y25Y1R3/msDaTUB
tRv6Ej7Jwn1LKjvnqCELg8IHCBL1BjM544Y4cvN1/3jbozKC5qYck1lgE7Y+tFVc
jd7mF6XN6ZJOfPGUFAGJXygpHz3+jKsz3ZuyvOkrV7kmm6m+Ro3Le81wkeIc9653
VwhnDqQ8ym6YZr/Dy2+1lff7W5i39Pj5KlBOXF46obzY3kNx96XLRv5sA9Jy5RVv
jM/P0HEmDL9+wP9LG3JjW9asJU8fLP9ZOAmduHEo7ewIOiISNsP/mA7rTR3NgmCJ
uzkTMNZ+UJlz0UW5/YSUAiheBAKV+QTalHFUtZZ8/DOnGowb7tZ/AD2aIWyUqo4/
UYLD/zUWq+VTZNrIGt7zFOZ/yaUAFBntz6IDjt58K+lbd3dgXaR5/r1ymXkkqyLn
L6VXZjUsy6IMEXzKC6cJ2P7TVzwNDxwolybknKTdB3Tyg7qoUBca9kvMUjH2YzPe
EzO6JE0CTNjKGRPUmaiWT5XKw2pHl9WBjhSlQwH6RACiHqoQ1e9FDSrMCEXJbheP
xQesQk+NkmuTyZIb6YfYnMlmXXGY3J4PjFrA/6wtY0F2974JVWBdUTXZEaU7k6Pa
0CkL0NTvJCSzTi7o2v+fncXwxxk57rcsHUFczWO0z7rB/MxQm3mrs1Gk2a3OWED/
57WHC7dnAyO4k6/Yaf8Mp+Ty/XixjU+Iw1VLEDHzNv5IElTJGcLXI5CgzgnrkP2s
5OJ5UYtqoJNmIhWO/f/vYMh7FVyi3ZeFWMsA8+shqn6rqJ5y0wB3MMJNkTebcKb5
UtubW8VL7LdcKAHI7BU3N76Wo0OaTm6/sS/KtbNDgJuE8BkpHZ7mivHFSaeSvPNx
HqQjw35ALm5KTQCOMab+tHBJOQu1caRiJBKZAE/qVcH8xqMthp7irzDmQn1HIK4s
EOiEsu9NujNy+UNOq1dP4RlAnLKp/6xaGnSp2XbumN3lz1cHKKxhFhWiQAUgGAW8
la2XBxZ1pNKP9in0Ia1GrYVDwQdWizaGmECDFpQzFwdoEMPVviQzxRGz3JSMlhCk
jEApC9zs28J3oamkl1fBzHxhUp/34OSo7KnU6Pel4azT0r48MldY1iHhC3RJi1Jb
AZRIIviLYblFAgC+h6SaNu9+qDxG3dPPyjx/mzExBTXlE0u0Jhk9SX1jta8pud73
GnfbsHbztwvC8xAjklAByD26OTmQXl3/zJ1bfEpIhXD+ZzkrnQ0ADM0ha1+bk6VS
YjPyvR21KxZR+yVV36aZ3a00AJFdOr1BVXxsylL2wcepghNj5CB7G6E+Ki3P/e/G
brqhTG1B9gmbSL2yMWoG4b7U/qu1VhHUHj7wBSbKRodcC+hUzO5x9B22Y/E6YrQ8
p+L2xseJTFaGMqv2tc+n9lrwrhcg76iuKI5VWuF8+e1xI+4yZkEzE9kE0SQlXnzp
BCWNmc79OFTnjnVkmgXWP8ceEsAtH9NMiVW9PWg8P+hG1gsWPCMjZKG0KiaWxI5v
xrgQKXg9cWoUj1mHiAx1naz5SEs+Q4w7gq/g+5a1d0hV+2pLQLEp1aj/m1xe04iE
ObqcbZ/XLMuZSuA+3TtrOSbMFdQ2rapM5Ngaq1Q3fKfDKk2YJImn6qZQ5c9QW4F9
Jzl7FV/somKrm8K5zUrOdH6qFjyacZSeTQ8Jymow5f++xFSi1IgJDqeeRdV41hXj
G2Jp9iNB0VO0YnDfbw2ieoYHF600l/5LGVWBF/gVW6Z4gSvdlldfFhE/5FVlLf+c
d9WPnGzPoLBG35geTVUDrVF51eDzJpKYtAiLuqZ4R6oiugfMVItga2YHXr8waEDJ
FWI41HCS7LlDusc9eP7DbsT+yVhVvuQskq6Jk3fHoc9R0o01L1DovnEgufDmBB/M
bbdKvPDZ0QRKLhi5vKURcK6Y14bTr6ftWHqNvrSISl5Ks83L+Gs2rUXvP7HZUYqR
a5432lYrCLVJvX6SIHZUs0GNSW6aspUxBwpMUU8iR8724Du9mbWUBxpUwWXk46dL
GgivFstwlZ9fgVoD7k9tTvDqtHDDdHAGfKt9SR+iLzDXXLE8QfZj1G5/6+HMEQSG
+jWH5k8L5RkpyI082XoV8g1nln1SjhNrRhFfnobUxHfUhs4XvQgyqKt3B2aNkLo7
9r3WekBW4QvnXXFoC4FZur1KoWMxik6BhR5gGBfI1KxQj3yt5sjU1AqoFp8gOQ0o
jOnpihK4boO3WGHnEVt115k8SqbfxWJDuF7OfwpfYIbCEzJiFqEFclv4GRWdr9Ey
IWZbjahQxwNGP3PBj1HaXw==
`protect END_PROTECTED

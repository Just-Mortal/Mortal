`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMIZ1TQZ1PIT7J0oMCXe2GwVx761NMQAhokenAhiEQND0vw+o85vqxM7twdrWR/L
xS6IO+KKQ4ju4bZ1mMi8ws566FjY0lPA/q/O8ybW6SqFqtVaBRG2Wxr/iEl+2wpL
gDWPG4U8a3vQ0hZLaJIn4UQ90WtbbPoP03FTgRzM3D4otwei4Ci9Q7Y1yvs2pK8W
jYHIYWNkS///BI4ZU/LF6s8Q81nekKOOhXlDfB1omcRfA/I0k78A2AksggIG4h5d
LkBOopGJCBBfdvUiunV3GMyGGcLcS5QrLSV3/fL936GalAOu2A8Z9KezdDglCI4G
hFmPVhKvdMFEtbXBni4GnfjX3yXRgbBr5Pt79vC06DNy6osi4AFQ1fkfigPAG1x8
WEPX5JoXWrtQSDwDYDu46reTN+rHGRTVD7qannp8aijMmTptK2SLSlOvXVSsFZu+
QxirfFKHkAS7+FY9Pc/hvzu9e2pTpuD5nvq88MEXun/wZv33v5FKCum9LDcxOzZT
bLR5vpLESfa9PS8oSfREgyzl3iGvBcdXrgqxeIWBhFi3Gnsfq8MHr2q5YWZv33WO
PKzsLb0prQ5lEqW6TjeYQyn7OaigXN8661QRh4vkMzsqLT5X7lfNyI7+3hU19neC
R+0HFZl+mYkirYJSWpfL227E1iWccXDp9ev+U4TvNEQcyceE/9FeWve6Ww2WO9/4
u55ZuupUH8+w9HrikKl1VoccedzzDdPVsxQv99v+F9LPm91Irb6ScMQjy8d0Ojj2
4v4c6gUfBgOR3DFGrvihH641lXmwT97SA9q4w4sV1DD9GCsw0yxJcHkvuRiOQZ5M
tys+PnAoCt2zAsPEXPeyDL+Ff8Ppsk7HyYA9FawCyUrYuT6rpPXHEFcsrMaCWDOi
m7M1xNk91jH7D1za5grFvB6IO3Y8lutSFMzTOwYLL0S6MUh69QmqEmODzTmC9Wqw
z/a5XX4jr9PUiNzymvPUOOylzyAsKbXzAAb1fPGwqShtFQPgxtru1aukzroZemx5
ONxsU1KXVGF14wg5QnBZHQXblEupe1J/YgKMt+OVpQOIoxWnkz+78FzsO2p4dGcV
LF/wYFvCiSaNL5lB5AY+pdiM5+4dKvspbncbMkY5uS4i4/0EFWkxnlshjl6cT17r
O/+xxrSBqWN7u+brEHFOOybh7RaJ8QgxEg6kTHMOaFjJiFvmn+SKO/+cRHrSOhRL
bUWsBt30EnAaqoRnFDMRA7ckYt0NwQgbpXArBzz8DU5bCNszpjmtwm9V1rZwR65U
DekfZSAewh9cd2Uz4atgRxkSM6AmDzy43G7C6pb0mS7CAFomZ3xUFjVU7mjtBjZ3
9OWJMqcCGn2UigYfY4tvOVTZcH3iL4orRG9ZQFy2+AwsZ3O79//oLngxtE36K0lh
EI5gP/Sy30oBSp2vVdFOtGwxcNxQnbnLcjz8DOA/bS6E7ij3xQUpSDV9h+GaBN47
NXZF0OxkFqWAgcnpjU81mLqjNlpY0ah1S/m06CSU5LLM4GMQb42PTgQQJ7jVUP5L
vU3f6Oka1KWQc1baX5g4gWgjpjOXoeEB7Qu2ZSlMjNCpHzi7+9x5LoaR3DrbPw+B
V2nVFXgR+Uben1z9nmqzqi7kfZc+2YMyZukhdMBBiL/fTi1eqEukgZjoBCdP4Fey
OvzlUiYCB0w3seHNjuByXgvxautUj6kXfKWQzCKi6v1FOK3pP1C8p4sQZi0No68o
VeTg2edfL96TigBPraZgUTgf3uiUqgZnuL6cwT+oECGRrH9/LciMsxznPCqG7az5
IVevyuuTdAkMaOlkGVJcWqozOYVzAq+xmLFcQ6sd6772RsbUCcUr0Q80yU/c0fQW
RBYAwGwa9936tfD7J0bhdjjPzzTeU6qN0ZiZEbnC4gg1T+6p6ujV1R6gm6gMtqkz
FUKDAHMpJqIWxd7Mg0CENI/Qqh/TypiXbu1appTRgoDpCGsus4TFowXg+7UfIwEF
mnSv25zfajlS8/tzujz4AUY4kS18jp2BVqb0BIq7rm2aWxkryanmLciZZaQEQMEK
JmdTm7IT57RXZz2F5Xu2khQz09nKVvjs6mDlI3PweRGUm6Y4WnPtkRKv4mtXeZDv
Vc5RGXQwsA+ukweOBgeDsX0N4CbfmyMJ5+XXT1yzRMYAih0RgOlmMBf3N6pu8/SW
qeXouLO6rOsmEic3+xLMbDzkR6xR1G89s+Y+4pkM2DuIdWfiwFB0JNunnY0rFKfp
+/cAcQ6MERYroLHGAzgpJFMWFLeDU1rpWfuM0S9QexjePPrFa4NN27bQi/BBgjCs
xDwVX6SKuz6WSCkmY8QPjsuHjRe1ZfQurm9zrsbBlqoNIGB+km9Q1fmxNOYngdxM
grJTp1VK2QKwynxNtKSa3ORhtrvLR7sYIQVOe8X6+Uyi0tq5J1PnmpnlMPUs0kw/
TkGrbt5wPQC/zgTPxPlfLTHdtXjDY/jGKShTwo9PeKjEAYeMSA6h3R52BulG81vj
h+aIzQZQm90YcegNmzu9zLMHi8KoYPzQr9fFLPYXHR2TFvqmQwKCGBQSr3X8LYXW
th1jyDdB0VYAHtHYaB1xP11STM7RyT9AyvVtveNnYzEFVyhiqA3MtKoYiC7eMyN/
IuZmXX6OqhzVraugPenBGDMEyY4VZ/QuXpjrqyOKpYImUND6LZZJy+G7yPEw078z
JY6KUmjDZUVa0PjL4v1BUH0+Xf1esgbQ6a7fJL4lKwdkqCVah1ilsuJkNYXqKrJ7
6V4HcKr4c2NPhTIjskh5Kn8DBPELJd+mYKvLDpqJnvGWLn9Bjwr646JH51yh1ru/
Kgp1XylSZY71uM8EGpzr65/QINdHC+QuwxBp2ATxoLAsqaoIpgVeRJHlm3BcVflg
vjDAPkYkG5yaf69Z+SEEmJI4H+7zyeuFMj6qEOWrsDbjE/CGIYqwnenvYIzXKdR8
DaVg8k0n9NuST5tABuWM9pJEfkjCRpW4PCTYv/LjLV71JCwIydr0O7l9poeTHXX6
neyeI/sWsEQdGUhNeFluRWrax1Jmzb3kVihAQrwxAhtTcn7U0xJRBT8wgwH2YPPj
0B2i/wcV+Vb5g2n+4DB7vR6xEfImowuJORKOWDnPr1HvUy7ZnbSpQ+/K3KCGDZFI
szoqWbpeUMbwMEFHXpJGMXDJC4mK2aFqnJ0AWikqerMiqjH34GxTj1zce9pCNQJB
Va6CtNX+nEfx/2dzVD2/QYEibHaXL6q8nHmrkSVEPDcuCv15a1Wq5OsiQ6ajIHLT
b9sH2WWvATfeHNoeLgV0xNNUdlJzscvGimp9vG+EdzywSPPknbNWQylP1Ed76c/C
U7X9vh8ggAtOXoksVDE5pjFwFsa1/lL3hRUTieFkz8Tdbxlxy7w8YKK40JfcfP0b
wWJD2TL608EXVd6FCiMvndMsVxWZfw/kf9ARjSQ38xMvXf9wQl2ri4HRcj2EtNbb
sjBPd0WdRz7NPeTllsmdd6CBqDu0p+8s93AEGpzFoYoCqBhnzU9sSf7ldI3Tn1GQ
uP1Mri2ptpkphy+L+U/+df2iXLkQMsI4GLNwSN/+yPjh9jJcujnjdDdQEVk3UN2g
dawZxOu2e3eTG4n33VFfunj86IFZrJFZ4ObVk6Ex4G8hkOZyXdTaNlLDFjlp7xV0
Yyf2vus3H0QWFPy/c+hws6Z3Gb6b14yaubdYzbYdMR935XDIG9TgP6DurJ6i0UWJ
/WVGtz2jt0zMP81CL4fSKK7khG1qFocWuSvqXaP2hehAcKHOn8HTytpmhWIrhn7G
tkhxHIQZB0Rq86RJABl7jq0Rv7foSmZ9HpeGjKu56MdMnuqqpdgwf+xyko5I2cjW
yJXd2fSS5MQuvFjKX1Gg6F4QTQckN4WnvDkpyIZUKAZ21R94yVpHDqRqkY8i30hR
ZOqfycnIq7iwZThwBXUjbwGyiZT2v00XpfCKZWq9WAJXnffGyAInaqdFtm/JWsg5
mP3b0/XKWpkwz72YHmceAfDAPpJoP780izNKuu4Medj57Cbe/6ksTxD3FGBolS/8
9OQBBYcxjWy9GF6lfWhb87W39I9lLFny1FbIKLZd85aNLVGmKOb5Vw+Q4buKqU+J
RmlJFwiXipZHlzBDSHfc9glPc48gSZXo7Nbs17D5bmUgFC+h9nX7J/O+7udmEVCz
HBMs4J9ubC8Yn8fVHQ5DlIo6I5w3AUgv8vRlNdaouqgB10SPTLti2AuC5ZwnyszF
gIiNtCR8v1wDXT8dYNCP+lk9s64GnBRkHVpUZqsqG9G5vZL8w0Pa/mnJ3PdXMW3d
hRHwYB8rRVBiEpYcjiXa52jNe2I/3l2vRUMYrth0hsqGVLuHu70qzLiFo+Cuh7Ir
0cdFwNg3NZXXlj0g+2ish1Kb0eyOqB74DK+Bpdu4J2qOldHSEkXEKhj+Gg76hTo0
kXVQDpO3imkw+T0XjdIo6Sjitb8bEBeygSFX84VfWN+sH0S33CrT5AAiOXywtEHu
FtdHetsx1VQT8dBjaCWZ01vQ5sq+iIg59ZDfaHHhVKIUcnIRFOGjbCXgOHwFLICR
rPZcAqc/ojkkweTqrtN7L/7z0h0Vy/WwKofZRCOmHaMk36dmLU75IcUtkag5qft7
LisSAtFkxSKKlIjze+AI43jo2x0b5OP3tq6tcVzrY+mdbplWDUzCTeRYfNhI4HPU
XN3Mz5MOXVyjGq7xJ6ULVuVo1IIsYmIPmPcphRaXX61Mj1SXPXrYYm34FKtyqllU
Uw77qcwBiMk4HPPUfc/jax7bGUGf9AhPx+2DJ7xdiMw/sZU7rt3U4renGV4hFWiF
v2wC8CrW2pAmPnPAWdIJ74RzXmhRTU/0eUZ3qynFPPLYXbdUnC3WyUzB28kTlYeo
UOef9NziLpF09yr3sG9sGn7012mLUkGs8YuunbMcb0Ja0s8c6/f4utFo6nah5nVK
ej/9j03aiJQpw7NTf5ZwWppeVijnzwvOg+/M8neBi+FoyYRJlMjwyX9vxE5FXl2U
8PYD82WY853EV6T0W03ixPiFcEax67MaW0mf48QiQ+ck3QRolzZFB+w1arQaZ4ko
NYbJQlqn2uZBAVXFJdMmqvZpM7vG6vxHJmfwuFEUVMfaPanwzSoLZKgQLFvHNzEn
bfyGqZZFXVS8yXRfPL+1FU3EUspX2oYNiZPDprgcOAdjb2UVu4DeaY5Aocl/IEch
+s2ZQUEnPJBznqNfgAUrYspqtgJ6Fx7z7yqoOC/lUNZIURKWuI1JjwznPVi6Migk
cBuf+zddHBoVEyYWrQT/zPzwnvNCJLs8D+yHuliJLEP+iIuGXQnuZDPyvQKwma+q
XQpLFprDRZL5E8edpm5rLiYskGnVYB3pRNq+GvTgjEIxidnLu5oOwF/FeYeRyFHS
OogNMpqG0WjKh2zhkPzG7Y0YFCLE7+YdQDnFryGlnhMiaraFy0YtT1dUyyveqNX5
SicR9JrktipyAun29isZLc+NM/++z+Ej0xKgcF9j+vv+buCzosqdYqGJ4PwJM08E
QDBZSJyBEBa+qknZCNXGzxLNKH5ShGtJh8ENyerpHjFa223DcmAcEOZTnX7pUmY/
VbacjAyBFwUeZ/Z2Y14NdoOQlifdYQMPfKysLiufla+1O6B8QoX466gYIpWsmJlr
cBgAdwTyeq9EsLGJB37nhgZXCnC+/7EvmieJMeI7WOB1fGxI0d9cyqfN29qzYURz
jcFAeFoS9erRWIGnNskZOSbEpaaDmLwR+6eRA1io3hDL5enNnfHKBlvtSQpElBLX
sFbOulmMFcEZ1cd8ARrP7nBq4H5JYHNGmogaGAS8ntFofxbFP1pkbEzfP1kgeZpn
/1T4LSHFqskJds896gD+edWSlsut9tCscw3SUtN53Fb341ZsqclfEvgUbfFhA2T4
onbN7w3DktPBwfeVR2D5a92ixbrcf9br+HuLZ7Gyl0WR7YeDh9X1AX89YOW7PKth
hYJ11jRKmLIiGJeAIAJtiWPwf8YXxmTEVjvr+rtfWAvI2k2bxgO5Mf8deSh870XR
V47HVM6gpCYoUAaKvayFI1dVGPH0qCnzZIJNpORet66xeek8PExTmoU1NBAcjbxU
rOALoKcXeh+A89s+o11Ziers09Sj4g5n6uFB5bSqXw334q7U/EwBq4RexP1OOjez
d4EMdka13//Moriu1TLZfBG/vrtsF/Eyc2JL1en0wIZoyUk4vp3iP8WBlUcRu4W6
3sfVXUHxOb3wM90dVqHtQBDXoQ9FDCgnI41IcVJrayLb1UZTS7NegBDTymQsoKhA
hjZMGOnGpYmGiNMh65sNrqhDJ5nNF4gCssOu7QWctr/KW1ruD5SpmUuTHAfFU05m
KGgumgn2OHRsay8ziRWM0P62tDNZNDpiHGlQHFqNVxYPQZ3SigMJKDY2YhxmvLhR
RZh6M+YCGbVlNrKzsEWWA1tb875ilVHdteEw2kN6o9baykpC/WRyPVHTuC2mxygp
v/whkBs6obmyYKe9ohiU/eSMMO5Fo6MgIYZWvDlyg8cNCmGws+IgppVGpPmpomPJ
GBTzMcUc4bG0HaHSzcUp/xqWnmMn+BhAqxkNDPhqBQJeMq04AxNfQJ/R6EzDIkpL
vxcYkvSL/JunxFWtFcOHz3gVLKfCfMx4dPKEeVnvqrRUHURm0U3PXz5O7Ig6BJgF
i9lClRNhIH0sGuxpBpwaboSvEahdnVJF24bZD1KrfC0BIScs2FTMQOO/htOSerzZ
2wEgDg6ceqBV0Rty6O8SXL3ErkzCaKZl23ac5YjUXXpbD3U+TmUAf3ch2q753GI5
8HQalfNQdUuUt3GsJ2OOqlRBW7wFUIjAWHttxjszZ8Mx6M9jQlxd1Vw6d+T6v4Ce
ydPt2QKDX6QIxErBH6BJCMbcgdw2TgFj1nzaGhDXsGE1NCeiZsSSL5MHG5fBRNbA
s9l7ni7egapKA4a/0sPqtWPlFmAn9qQY6/Xyyf8AllLpKSuf2a6owclAmFzsCjSo
iZeQsotXP7X4FMo6l4r12i6iJwf3uhaWYGaBvBok+5TrKncjEPPAMeobDCT0sFSd
UhjSNowf6RURYbYw+/VT9AKnFmomQqFssLHG2vuP56rqF0I5HoVd4Qk4EQvaxFsO
baeffwqb+zie2Birt/IU3L5iyIH5SQa7S8jH/YULFWPRGIm3uGuFabfd/1oyegty
+StPl8mszC7MjxolyBEScfVRe+dYTU+iJWPkgjfzcb6WMZF9MJQPE1bjHOVf+LX4
Esl/AJHFDIvqimX/7xE6HpTcRmrkyJm/81XHSpxju6Ed0obtAUlBZFRl/4HOxh/S
xBd02Zam7++iZaYglpBLg8IsE2SbNw+8QjIKFv/JxsvGKNGK+m0Acd0zJLMk5Ta5
43MTt6bhnJZ0IWu6CNAmzM+5iL+e6SpwRtOMrcxx9GFkkeKG4UNfpzP+D0smWQ2d
GgheCvmJEYIQpc//E6o2pOacM5iGZVhOMKn1bg4B+6sy7e0QxJVxzQTxAlHDc+5M
aFJkSgvcbznsHkClXzeAUKys353tWAm6CxxgOHzw5xeSdRmEHTICMn7pl4t6Iw7Q
+TZ+Zd7JkfP9oK5/3e2V55s0sy9FGqOkXEcBOTwFrkxE7Hqofvz70u8EsbDkiLcK
1bG+ucTCHfHVwLVXp/HNKTcep/4fcbPp7PTp4D0FBW8iP1Qpaxg1XDSu5BEYXb3F
U1sHmNLH5k16sjbaIGpleKtFhitPez6oCqQWodLOPXP2qgSgOCOY5vxU5AqBchip
pyVNn32MqOMKCdvIl9cTqvD024e4y9JfIflzaTbgEyoiCtcuDu06TkO6GA4WInNW
Wwzsmo+GM1kIbKwfE8V5kXZ21+8/r6r7cpqoDdUfIfZXIyX9Thhe4xNy4HeNc9gn
DTKSbnT2bAvg/p8JJq9opdO+XpGl2VO2zBM3fc89CplnyLQljAmfkKdUJRTImUh+
hLAJieYorX1uONBK1lFyuvXRoFgwh4Bb6ocyGOdp2CtEtaD3P71jg995B7kDpIzc
L74IUVatcNxSXn5qfFejrBpUOeqAg3Iqcuzy6iNGPvUCJCi+TZtcbA/F/Hlotz0E
oS562ibcEkmJyUt1K+peQLWjaSK7vwnG7Qa7ET+BqZYj/rMdV47J+hph/POTZmxO
xly38O78PUmcBgfMFxTVcIDv/o239MNHGfeutZsabJQmOcjnNRi2nQZgAJjRAc7b
PaESK44h2WnRibgBxl8IzQ3M0pj9AoroPVSD5HF++0Ttq1l6PWJsACjYOH9IdJzZ
dLwxupiUnDOneU5YUy2iPtyEizmTUkvkFFsZQNEhwXkD7snpOPobOk2QNE69CQhH
l7/EOqnY1PoYUa9fec3mmCocOS3Se22T7bCdrmDsKkypH/Scxi2PqDooS+LDXGDW
/mZpQ/sQ85iWKDUtHHsULuyKerI2BhIjyJa30g5FSMWmys4udd7QnHMn10hVUFtE
ptEr1jc6LRqTOtyLamQzrOKMO/HRyoZUOr1XkjsI9Dt1tF0MYh19S8SXHMyArKZ/
Sd+EzCrgRn1qK8Qu5Iw5RSXdWy65X1diBuFp6P/izCmBvmjUAKi+Ab/5afE3OuHE
5dX41V8JRVWh0D3JNRsr92D4RsyLW2rcQ28qRkHDPUp2I5BphnC9R6Z+ZFjNSYhF
43je5RucI+76y1rXTgzDACnzHvD+sQah5SkYHs0A4+HOsFFMbMR4gUIzXKQeSReh
GhJOywl0ToC/9gsD1gT8NRRQBNJHnBDbkOrFyXdSXOeiROL0P9LJikVmXaQj5tzL
dnBpDuYctTMgE0natUbwAxqc5LnEfK6FWB5h2Zv/UZpWNMbLB09g2ezh+8OmWFNk
iM9LKkcS2v30lMsTleL72FeOWWfppqQLMqqmHeVmbJw=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jIu3I+XItkw1UJb+l4CfFAlKFzNRiSy0SXGYcb+mxMzZuR6JpZPOm4A2kS2UTdag
blFjKWEcgAoaA/Uva/utAqN8u1dxP4oE1XEzj5Bcc/zGNTf9z2c1SJky4pbIYxU9
xGEqEEwgPwkOsIyxwCSVOJ1emjFr4ZGfQaHs+UZ/hERgkSt4Zqxu57HLhV8da9WX
Sjj78mrV6jD7ic7sv+uqSXe5mGUAFRCiMgN++kvxu3Syf2tkN40QvoFIbEaIxXlm
6RYPNvrZ3nNBuVq7dlbOEnvxYH3UM8W9Qmw10/JmLLqcVDq9ZOqLIRFsjerwkGtA
NvJAe1Xg/MzfAtMJgZTlymTYgw/yS/Y9sNPhIhB1TW0r1Axcsn2qVUXlAa/inHpL
NLfj9pr+wroZSDDk2lXJdZaoTYO/sf90vj23ACbNiHX/PpWrLwIsB8At6zaWrtgo
apc5sYzgnLc8b6tn2trXmkC3QZQDvmMk5tw7uK/0yRpndOOLb82KQswstsLi+MFy
DiaFl1rmUfFQNAfYOVt/bTsFOcIocTsTm8r/LgBADdHj595AAJD5+gLu4M7oFngJ
3iB7tt23Ln1UjvEWpm9sMqImduVdKyX90KyYd/0lQYumCw7utjgsq/ROqnHAo6Du
HyUnqDFaO9tV3iyy8i/RXH0D7Dx+eu0eEEgmh+KqHI58HdiNnraZ6rrcQQ56Js/t
gZUF0VolcKNgS/JMCzhmadXkCV3QkcP/R02710Dk46SSq4qsAfK/namFDjJ7Y1Tx
E9t3W5q3Tzw3y6YHRo0rEohvBCCCpr5XE+DBWGcv0OSzmUEAmXuOupgtxnb7weI1
W7X5aaeTScC4s/S8RO6FsLqmG1eG7i08+0SSMVgoJapOT2TQHkxs0u55D4IXJnSi
ZvdYV738OUMq4dtsPACaiUFsG7ou9qvucjXXpsOocaTqWR5O0HFa8XWFOatKyd2Y
PI0l2V8/wRn7giBUQWWHTHUBwMiSWD/XcUQgwvn/ei9hO9ib4IiXoS2Gnuq+NJkH
LEcyj4xBdXBH+PwmBLNqCYUmbUc/TJhDx3yocMxbXwpEeg+fu0b+AD9d7KTcCz7C
0Z6a2XYM3M/intMmdOBxjAlYs0Saw3qJ6zv20C91UpprWIJoyzD9T5NcOcheqJQL
afyts+bjVL9n0RhzxkDxQfm0mFQt8CiW7rS1DuPj2CISKDBXhSAx5J2wIQadKXE0
WyJoW4nP6UtvyPvoCgVTMHFjYr1YvWLCN9jo2eOqn9w60pJSuMMMm8Ce6w6irgcY
LEtDSub0YEB/lqCAyxpu9bzAF3lPi9+17ox6rxaIMamx+R/bMysmxdUcwCVYBRh+
bkEiM7+6fngkXNdIqO8D1/V2FJx/CwdgKBW7Kmjb948xKHUjVY62z1hs+sJmvMw4
f0dN/BcxE3+lNAp/4j9NJ95s10zIyi4rwkar7d551ljdztw07lvRw5H8HXi11kin
t4q5wSdjDzyOtYwWcHkUybo668Xiz7rkYYJGlG0FdXCRorN/MDEkTnPhOp7BuX07
By8+lyeLgV/iOccLq/NNBZcAvOLzsrLKk/o6twY6m+y/Tr1e/ZlCzeUp5/o7MqB7
1ZiEcyQWNOSIh88dA1pDxiUeWu885OLvygNQ8d49ZMbikw/jVE5J8XibCFNu8ZwB
74xr2ZceEC1xMaOCm15JS1Ixe3KW/vSBD9HCQ2XVRG9C9bGqCUB/r2RCzu+QO+cv
KtL1MDpajMmqYp7r7MKUKBlHI8CysWlnkfJpsQr1Y1dO2z8720QltBuFXwcukEL3
+IybogIxQTnhuVdKBfrtdut0gT986hpkEwe7Khp4Mxpn0Q4NpbJqRKfkdQqSjYvo
Kqv5al7jSibajGRufSu12HyrSAwm8LmU/y2VcJS5Fa3NJfWRRsUk0AHJyqtM/hmy
dciTxdbvoXY1mQxqyiCvJmnyGsJhj1iDTOj6b5dXhuwu+K1RidoeMeq3h6j2XMyy
RnQUPzw1TSN3VFTL6d2tkCLsRd7jg0NNy7vTIpOZX8MD64YKp1iu4M7mBjgGzTVw
zcAIW9uhEo4aCqOQgGPjw8RqA6VFXG2hH1dMeSiEl35ruLXLusmdnBPNG+VjVnIW
DUqtY53P25NLcdH/EFvoH3zDubJcOJ72rhRiyNWPu3mAOSfNH1wB21ONCHkmisXH
00VxiYbTnHuDC6AkBXPJLPiVmcBOU0f05ea7SDza8PqlXoOps/IyduByNlbP1cy5
H7so4y/aI45syP6yNqa/M+pqquDln2oolaTGVWahD56djF3wp7pIJkqLIycYKvIg
wZUGeu6hO8DVv7m+8uMQ9fioi189KT27o9deS+gNqUKsqpgD4AE/owVgAHMGucT5
Zgge2XTY2exG1CFa9F2gXvZe+6WfsivB9hygzPQfywjFKjQ4cqp9qRpLhA8ahU8C
G/HDowq+gCtE9dWaMaAdPNwF4HCt9+dA976pc32ux7ud1yP+upKmfQvjGSpITmSJ
22PCIjuZDmAwX5eyXSultKvRqpSMWWytF4cFEXxumK9ijxYUI1dH3aNTZp0cxuvz
VtnoQ/4O0YatgnG0OsnP4CEsd6zJoY5f4DcX/1FpeUfdnU6ZO41E4osyVROlrxic
MOiyXdZA1WxU+KI3Kmf7ytSUlXZfyodB1qmU9RGlPmCzfk8w2Jpk/a7ehhJznqre
g0EpzN3tKZhBwetjpe25n+NEdgklhW3zAhqe+7sxUiPvr0wRSe5RaJUjUZhu/vZ6
fC+OxdnopDcZm4YKTtdREum0w3rLDqVbH0TywL8qGBAg3KKYxQRsfiuP9suT9vLh
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46J2KV3CVuAiBWKBBTB6tOnKGlusl6MWeveuK2uTM73w9DPgbpshhmdrR8MuQV6+
PfjMOAbntdQZ8cVUYaZ9+GC95sE+nQEVOTycCZ0+bKm+mQW5huSBa9W0YtiYtzEx
w7KOQ0zeH1srNcW4qKDs1J90nI40TEWsl/hj5Tkz4oo8s+QTnFPqpsHYxBKTS7VN
NVnB1T+/ywrTuX22zQY9Si7A7xXaPbEFOj2uUFY3K9sIajAAowgjIuFX5IslimA1
kzaKAdKYW2FGsg9W1c4lmWnHewvB425JJAKBmh+vP1aAmJK6zlPRSVaoqOO/LttE
Z0PRdx8rtbxOiZzf8TW8rpgrvaruRWxafJ9W2ObCENu9JgxGyjBnx8tMtMtJVEPU
/PtI5hmxcqpTsFJQ4rO+nd1S4UBYBSSpCu4U8N9NzXK4HZTjg8U5lWJ2xW06tsxl
Fsf1oolBWLq5y25dD8VJyQTCIclA+AXUDPbp54Ct9uRqvV3njMI7xR5tFvf7h6uT
InRcpZT6WOyCj8QsKEK9EODJTp89mCgeoic463BA7mumOmBd90JCyhEBn3QBZRUB
uQ/igXc4nZwH7R2xbueiWlzxRtMxxZKm8H00V7snryPI9ZW7UZchvkCFGvF6ZDHM
cM4btIXR5/6zqGRyw5D/lcNS9jX9reuRurtQu9+vYcaB02CWXebZ4a/+VnbFP0yo
OXY9qhOd7wYASu+DNnHMu7tbn3PszcaOtdTNKEJ1N6ICkY8bcbqrxKlhk49Bf0+R
HuVTtyk5ufYU3tSeVCvuN0zPFKt+J8LMqMytNuYYaPo=
`protect END_PROTECTED

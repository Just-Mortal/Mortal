`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Og7WTknejldELZEZKXjv5bSFpx+UpBYMOxR1NzTZ3mIbu5gqReRe584r0S/aX6EF
PmAlG/mxGvLp1ti56u7u/K6mZRO4PPOgOGHiSYafwLpxvJEqcyPDXAUfCZr4ccYS
FOHb+chZA9FOYrTqZ+bITdNkYiHIY+bsao4cA8hai6hBDS0iTLAxuY7y2WYzIRDc
+gxNR/pE953hGvD4ljZBHMg47TfLlMVqDeyKoRmEXpSCx4GXIreCwi1ugCjcD93X
QDm5MmPKr5cwkuEZ2062AioE5DmTvJ8T3H4W45N8XobF8qGE+6pI5ODxb6Z/7G8M
5q/yEZGRj2CeTgu25kYbNXNdCoGp0jjv3pgxZ0SCrMNOtc2pFEQ6hO30d89LFpqE
7mdYgn2CEBT2W0+FUx+FiqbHP+H5qsbe6g2Zkaf1RuRTmOPhFcqm+F9NxhPVAkUh
mirx02yEJpsnEH0lDJVBBNbhiscLttFrN6fk0WJM7KqyVrZSkhjDduLiDQp7yijt
mPsTyJ+s0B6chJ4UAezAKroYekdKvKAefYt5Unwi/DOKuPzj+atdJqrPCjR54wlz
ZmbEpItIa/6zzLBPUhooySLk6z0GAwYWT4eCHAxuyQLa4jryk4Zz1cX57+3gPpNH
S/pzM2k7NHUGBWXZA7+g9Z4MTiUoRGSziXeyJtFcR+dzTueWwb+jBS1eMdJ6hto4
UehF8MBFgUd9Rybklj5agrrUbPOXklK4AcICx9y99prHOXRcUkA2i9o0gQCnZAEb
/Ekpd/PM+W6EDfvmDrGVz5tNVq8BwsvpSTobF55kGwt7nHl7vdzRvrrfr6rhS6k+
kT6SVzNi4fBSIkcJerbpxoM2fPuMpX7Xm01qg+OvQfGafT+88c9B8JjsX+RKWnV4
R183xxc6f+phUf2O+a5sv2EVm3tqBAAdNiVhktPrYlNUeQz4eEl9gcQYZ+tkb3j4
gmTIXPZJSDMw8yI8V0up5xjJJa2ML+HeEOvKiuuFMBasYWshS9rAyUIceouimSxp
cLnG7KuAm7aBec3pEcPRYqO18GV8cVORoEdahyjJOfHWWngWgx4Pf91uxWXpqxDm
BLV21sv9GZS6Ty8EnAsVTliy4t8W12bk7+DRx5BXM/UlI5XZ6jJUGgF5kwNipBJu
v3EUfHMBG04oxPOnipGQhSTCPvWF818pcb/wpq15AaXNai6CGXxTNUBsd+5Nlhvz
z92SSZudHrWxe6QNGvT+IXqXAnpoolMtVE5iXoJSwZCABI3aazhBgqZvLhzWL8DA
npKpLGNYyDqgOZvXwImAzy03lXIbERcFVjAqDR15z5RlCZdBRO8BL83eGkZmL+Fo
000+pwDvHkVyWsML3oIHxWSdAWnmas/tz57F6tfkbN/skRKdRhJGT4G2F1AtwcR7
+qnPJD+eXSBJgiRRCcZdb5hMiNu9J7pRn7GtlPgQNrkKtThCxQ8KXl2+3qEbmbB8
/JKkuWKMWyLBrUb07rWOIz25t3WhUw2LcHkIQjEhOj6RaSwz4+12hIRS2fEheimL
nfQ7O+apK45dkiUiipp96Lz7EB/baWHdu0NZrE7kZxxhdAKi6uRBiH0vpanEGH+B
uKsQk7sIuoIQi4n1fVV9+WsQl7kxuHRTCAB64uX/gpYDYZtYTACyVAYGgC6HWv1p
b7z7bAu2g3InFflLMwvctPmzkLVTRZX4s9mmUNv7rTGoxcvdiD+LMLBH86lJZ15y
mkA3oz992q5aj4Tts0zJ2ZRqTrMc+BPVltQ4WV5yPAX6DjYIxG8oDEhWO+Bu6MJv
G7WxPUE94dQeVZClUaFvOcg49r42X0fFz9eR29v5+zTMYHiqhleZwSUtqgRZD73X
aN4G91zchueDjeCTOAVjkzo9PifMJT7tJug0SdftICagQBYcWiwk+QGAP4qfq3J/
1KZqSoxYN7S+fqAXXVYEjudckiYyUF42fKZSlNKESbKNPhOBCTDDxL4+WTgD5vxT
rEaEjRsRskKmJsK0iwTtaaoyNMrvQgRXKVsF6pKUVleMzJHmV0YIQZQpLWFdEBB1
xrc/g16fNk3L1BxTpa9AR7v3CovrgxD5/uQiZkMi4MPgLupLuIj263J3Qa71kfqZ
jHupPfFpOuJbrdoxt/vZlh6ZgxUGSlNnGTFYWA0nQViARbNNIy+EyghjUZ0F1c4o
9lNHN+jrNRm5jpYP5SWnYUQYqKDCZjbVDs0mxbRziXc3muaH/MiZxmo+r1VHf5+7
vusl3OyMLi69W1UJfHW5Hk6I0OR0C9aahP1N/ixKH3oDE+5TUFgRX0TRyNpooUH0
9lUR/gzJd8kJL/pVTtpSTTrCubqOUk4n1hq4ALjgPbN1V9l9r90bOGy1m6lRwBHq
9TDdJs2emEFbM4XnpL4bLsiXc93b8HKmy9URVJv4JYxKMKGDSYgPJOMaMFnO/t3s
HtBSIbi7sNidMBfZEFYEdLPLwuya9mf1juVZqlc4PIp3hC1AVgk2j/Q9z1BQuzdn
vX9u903lpM9Cuw+9ei6h/Tt5wSc6McSTv8YLC3xbj5KGZC5K2bHlZK2WL5G4QYur
KLei1lO0I9m76oC4gqRyPBdXVWANeTu2XG0x+ntD25GvyLcpTLYJw6CrQRQiiNNc
GM8TzBa23ehG0ASOxupz6U3XWjeFPjkH5R7OG8eCjDDvPOzu0M3LXOLYHd9n/77W
Tq8z1f7WwfkzkQK07wi/hA7WeN/2VtVkxolMSZ2T1Ihzd7XyQI8MXR253+9tuLrf
diRhulGJNncMdixoNM9Rm2JJqQWe/v9oy9M1AXEdEl2hEu5w60n0b54rLOiVERLh
QsmOZPqyeMSSyPvRPFK5/ZMlZyDj5XIjp7pNl8v9d0iK01gCwxlFVJ6iluDFuOYw
ap3ngzZi8xlecfyP6tYOElfCgmNWyaUlpuClGNE/sGCca8ENXY9LqWZB4Dx2yb/P
HxsNxAiAz9Wk09e7fxCu/efzj9MmiPQTUagH/9zOcJ5yRK5wtxyDm6om59QE9J5o
ptTXq2EJ6wqkoHvZxAc+vFhOWgG3JNCnQlsw+stKODTQVvlYC5vrtd23HdLmOf3i
e7kIAcsnu/SmZBFVvtYMiu1FO7rrOpXO7rmonOhoM+aKDmZb2/xzpdNIYZSBW3iC
mT/RBVMw8fe6KsS4fyxL1deIYYwOzUAmgIBYJZ5bM2RxroumHwDzlmUJAS+7Urzn
+v7aD3TpJHHSnoV+4pHLlGKtcAQ8XfPzxebVS7o2hF/xoodfOjhr9i3EkTnva2dJ
jDjb8OBixLkIKQNI9yzzaGFTMkFv8qicRlX3dB6DsUXzelltkC8zj7iZcIFqSVut
SvzPSMgzfl8vP/io5P+QloMPAkIrrfuRGNACfnBsJVS4mdVi+GH092eNXFtivFH7
RNtBhDnPSJUxsAfc6mC2AjRuoLCBbb7YQS9OBzTmjST4M0WR/zBt+RLt8W3xSoOt
wTp0VEY9c0lZFVawPvsF4DD59MTYgF2+HXWSbYM0ryl6xlXzgL5tOHI9zsbmyo3i
h8POVxUzaS6/VUwUkn900jf10mjIN8ufdiQAEs+ARROSdsRy4ZsGqBHdwtmyZ9Q9
uVF/FuMhQrOBE/j2CWzpLfNQyXCgyoCqtK5sXLm1cF7uuaOQXotjRnAAVGITWi7g
FJMKJLTJsmhVB1+KTi2SiK5bXv5gHo/01VhJDa9DEtEPoCPts1GgFnYU0xQ1y4K1
Zo6jpPPJSmiM+/h5/nYmSwG3j5x1ExBMtDpSO3gPN0S2VqzRh1QaPU7nejH+9Py3
bvRzEWBOYFoiMMlVdJaZ76UGOpt2Fw9seB6p6IS8MDF/4EukoCn9M01NptuBjNBd
rWz2nyD7hCcCN/JcJhTuGY4Sv5brEEnAS92m3MQurGionsQnR9uvmkRsZKyJm1ok
srqDFC83PBrXxeKjDKQWj8KmRIc8+nUN2jw9AWexhVN+gvmmD/+To3f68rDr7ZlH
MbZE6JjQwEQUOLdvooQKvhABxg37MMndnfGm3hdm1HIYrhXyBO+CbHN0Me1rNx4e
p4ophmRlJbftcSgPCggIPY1/B+MOUt2eTXcQ1LxEuxwzk8LN4zvq/jGcqGRD6dr7
g5fggXGWUjXdDYPG5CtDIHnajXvuYTwMk3OxGhZfaB6cHFvMp9OySdyMgZosGeLN
IqM9TXnFJMbn+zmlZdc2FhoMQD7xTkawYlYBQzUsB9AG+FC8mdqm44a00NKmFTD2
3S3HWLUWTtbVeLFwRk0wG4XH1QjyY5fwCtwvHeSKdFt3bowK1vFUzyrTxDzI1zWG
rQlGTSJjMPCdC7y+1r/A7ndax2FXG+X2a1Bdo7LlndbFxqz7sdxVFYBPHKEEyjyT
NAiSZN+MzD2jq3m4NGs+cwOvJhcHisf7CnLfS0uTqA89R2qz+Xy8y8JgKdDr8o87
ddsSjhUQHTkY4Qn59/5DcdI7LU2X1q7+xk1+OL/5Ob+O9tu2QiCpNhLSw8aExJ31
2NrFehHDpuTD2DyhQZ3x3G66R57g8GE4CQkx8iNHGjjQMSof3WxcwGnH+aGYdylm
lfL8C5tpoRx/Em60f67flRTfrDg80r4bBPWurq1QuTq/nbrgUeyYExoS0XBdiEpC
fuAwFpcCsZY0+wM3RqogsL8VLjz8VbptisnC36Xa8NIwxRY2Fx1oElxi3Pyk4QQL
6q8kBk1Ok9iPpUuFkcYqX9q1iWBbCRo9Xp/m7T2HyRY=
`protect END_PROTECTED

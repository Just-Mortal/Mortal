`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lzt4BA2Xh/afV0iVE9bX3VyamCCnYdyiIUSTajtAXQj8eQd4rW7UAqhR17Zroyx1
AsnnYXAlzw9Gsj7AqDPW3UMOO6MOhL061cUnqDc/Ro40QzJD4iIeJwdnfq6LyTkJ
Sr45jSirlfCjWP4ne565FHQAgoQ1JppYnS6qbNoGo3VSjQTuEXsFhkTZIy4CXV8c
4fHA4WH8Q0YsdVkYLRPiowPjigM5+RTY84FNXnpyjyrI/Yk0ETdJxvezxwyrKgzg
t0yz3bIZvTb7g3vB2Ya7elOFX/t9DfrD7TgDGE/445pVqNsw6V/g0Y5qp5cuteLP
y2BZ1/RHlj8DUjjPlhF+390qa9NZI9yRElKpMEjoLb8UY5SDUKskT+R1H6hWpTRn
ktB+wjHsUGGBf0Y/dYfB5Z2DeV3VtsgJY28D38NXbVJLHttSyM3jSD4KE4OGtxYp
F3n3a8AaqvHxD9Rwzyf2i8OwrI+Nb+FesciR4zWSpMyGXZB6Gd7+4dvlVuku5CZc
qJIOSEXiyrpcEWP6Q3bt3ebvCGSbqcxOg/EEN7EuTZaijG1ppzHhhj6PcYnWwRfy
RSv/y5W++CT8FMMvDnB9rwOh202WbqbM3q96MRjFxEdptjd+/ZRiNrqoc8ukUsWr
N2Jk/FREiW0RJi4nk3zGO59Y93ZTszmoTkM1ab6brVk8kWASAlCpJjiiYJozFpGK
ekqks2oWgAB7agoP5yQRzuc4x3VPRq1Me14077t02PxwAXmGjOdNN2fCdkn7Shsc
imCODZUvQ4FdWHzeuk6Rlu3lqJUocvLryeC7VOFtORCRecqNeL+LrYlhnt5lkQax
+0PuenHTi+XDsPb8tbT00Ik4unda+HZsVwPjzJPlzf9pf9l2E03a6wlABk/NTqm4
eZ1PxJVpRLqA/8jBRN0gjceGXtRmk7jEbUEYc6DWa7ACEsDY+b+KoN818WGDrStF
DUXw9gwMT4q08ExlOVIgn4G+h1efN9RGMW9JFHhwrhOo/J6DHUI3SWtflfu7ILmV
bDk4DPDwBHxiZ8qvN74HW01G+e373GIpsOLKn0QZLoY11ryCc3LXVwDqKm4yHgkJ
kcjk421p/9BSPGD69voBuk2Me8G+UK04+OKX3feO0YVXp583drwfr8pjl3w8H1Gs
MeXRX6XAJ7zl15epIG7XC/3Brz7gjIp08j64CscPFb0bAzOC3OtLOkRPpgpA33w4
tvUBgUcVi6e4nvlU2kG9FzoCy1P1yRkSE/e1gPgd/70=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Q4tCQx1obPDPXGpzAZMOOafjQIBWBgJzSGwrZu8ucCnFrvpFwBpjBsqVl5LPFPS
GsAdh/bTJJ9zuS3udp2awoYMSy0las6Cir7sgGz2GurbprmKLdBSNg+t4Bm8gDG9
vhx2W+RZBxMAIXc8C7fgQ4VdeOFUdyInGGjW0rfCiXO4xz5EotJeL1WrzN73wnCm
6sk15NlmA7oHq1YsyBYlzKTwmGhtz/uNpT4ViyWLzFTIsZgp8A4mCshbQUsSGZSq
HkIISaw6mWb01hPUzfiYlImWv8u3fkOG+gbpLxO4nrbU06MXLT0BlKvSzpsXz24e
6btgFRrfVsRrhTVrKdHt8YvgB3DcUAecdMm3m5ZQTtsWYzDsF9mjyaABZVIkv9LU
ehnFX0MymYomotXmi3hgUTW7F8cF4eQ3/if0M4mbPHriJQ2tzCAqvik09exmwQjv
iAtP4j8fwA29BEFSy5g9WQV7Y/tdD8bvXOjqfYBdN9HNqKlmvf+Vz2/GnL4WNpWb
HpwmJa3rD14qhUgT182LNENHZRtwJNYkAwEmkYvgs6oHjQbm8sWz6ilgQ28ar/Bc
anWmUwjU1HO1UU3h9/bgtyIb9CLOJjAaGkp4x7W1DBbo4My/J6lXEiiTXy0C+Qac
yUy4XJ3hwAIzqS8VoQIH89iRr6Be3me/6HPRCEsP7wPP8qrnEtVXXUQewESbQwqk
JYONAoScY03qzWs7VxRu9gPt1l/Qo97VQyMkBgAhw9hMuonMMi1REU5PHTbLR3my
m9Jdw6YhxZmOTAvWDZn708H7qsq0Qu8e/nP4At1ce18kq+S6u7l4EpPU2RcDYfs8
XzSi2Clgw6xMElHfW1pE3HHZnZo7pvdWu1kbTeV7ATcUwJgTmv7v7N8THsdq2wbA
zcUyZQiG5Zx3vbG0w7HWfTTVtjCD887kCeY5/N8txAjCTy6MyTWblhDDwI6sTSKK
nrWEVek9+8lIqOLLp2VBoW8JClsuwqDTXpVsVYfPny8yqE59QriDhPJ4OwELxczz
ivJR+WUu/YDdOAB5A6Gmtku6Fk/fEixdyUL0F0nuZnjAMm7oLkQTBgIhYLqUhxzQ
VUJ9OmHIw7Sc2i7gZkK/qarTIPgfBYn4AwOuBAtRoFI5sR9Hby9s2O4hm/BQc6JR
s1wmB3McTJ2buwDK8ixjSZbZtfzQiOktWlJBDMdGnV9e+ZvkUbHzuMYC/Eg7G/F3
oHJWfdM/oDydydtJd3xpuP+XII7pdLHiFlQ0bDQDaNH81LkijK9vAeDSdj12vuow
Hcq9vfXqpoGtXNvp0/8Za83m3GFz9YS7mKSJ8GMNbpqTbV9j1GAV6nkYgFC5ATxS
koTKrgB4IylrNYETYPJ6bvu/rZWUhYh3DMJqzE7oYN614KJSX4gijqzi/AD3OsLW
U0SNnZoO4O7jZfUn7KjYIgiKlc4q0ncToI/CyVh93LS7FxnIeIMIYS3Y920+ropr
HqZKXRxrWxxyIgHFlqmMBm40H2PbjLoYwQMVnriQSd3Hxx/BivaAkgy5HYRRYq0n
`protect END_PROTECTED

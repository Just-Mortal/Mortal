`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtL5xw09EnsW//6AGa7gdSf0H6QVu+G1ToBx2zskTUgvvJCqmPcfVoBdJTT9Sc79
OQvsev961HT1AAw58SXs72dCbuuhppszaD5FVBmsBZxj9nwggWWWaIaArV5rimeB
gLqkasRvpCuAJ9o9MUakVbBGI6lAnY+4MAQiL60FX7RUOtZ8OGWM3c24jUjNxaws
KE94DCX639GhIv+oAifNBtR2CZts8taO3QwDX1NOp7UMdCCV1BPqMUmAx94y/oZL
hwwLZNGBTHNy2XCCUFYyQBVvM2st1YHl5avygB7jfzDtgRg7GY//6+XmYgddPBLO
8LjR98i+h4ov+GQjZSBxRxHMzLKiDO93a8ZfLgAPLFilDIPNfkBZUknhFT8ukQuo
e3WOlQrl4GA4Iq4jZoKuQCcjbUH/jeLw8ADC+SCJwRCihJ/PodeYpkUoevzauI/c
gIpV9Ps0nVRX+bepcPmXS12qjjwLDD4FV3ri2lgekL42+vsR5JJgw9Hq7BOQODpB
S4mnAHyNqbMA61YH028S6m+vn2PxxgQcL/OhYLvMTtCmnXrnebvsXapa9QIu65Zv
3LkzV3+7c75I9jzsmuWOod+8kBAb8A96VUQdRRJvrsJ56lsQOn4x0z5AD9+8DB30
Mgc0b8Zq7PYWA2umdGOLTycNLKsKwP7dpiOHugQRBlGaJ3DOFa0ThVUGmHeqfx8l
ep2SM2nAdaBgbND4Mz0MOt3/ysVux3rdIXVkFEJw2Zfxs8Di7pXYeZR3m8ksyX20
CIg+9+ZTYoxHq+Yn/hDMPl4EMvmbTWx8ieZU93oBkx4T3gOrEvYO7Ezwc2FkjFKR
mmGO0zU5Gas7QDS4hMG9LJ5XBw/k1JO7ztgIIQz/QolUFOSuxY37ZXJYt9MGS+nJ
T0naG7uQFUxkC7A9d6bvmQ==
`protect END_PROTECTED

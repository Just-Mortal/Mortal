`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vchKaEiuBKVKW/BrGkw/fHVaUW+b9DL7GO+kr0nVbHDx9SAiynd9fP1RYORxy/e1
ktZHbkGFYbbPQuS/iOJ2Mzi7rV5BnfbQmgwneOZI2rBKeK5rz+R/Dgtb/XAVraMC
vcRyPg5Cf5oMXYQpzj/mqOw+bKsD60ImZRI3mW/jn6m3bnXT+T8iY944A1yiBH0o
GawqT4f9bzM5lSy7uSYrwjUNfQWHJnPpH261EiinQbUCydYcI6tqXaYoRwBTnoHi
6Sh3f4RfyPuAav/gJb6unjvlmoFOD8lhQ1yxnUPec6r1RJstl5Q42idbSUrqojhr
w+w0xgVhflkqAE6fxQQ9lSqbEfwtRgAoqnVOcjAG5ml3sVO8y7SJfAWH5qYHGjDW
bI4w7UqcK47pcxuB0hPIvIu6fzDiNpEEHhHaP6BE/UeUXMFPV2c5NdgQ23x9ewR3
MvhtYa/HO4bAkfLCzVHD3wo4JltSsjQcrq0SzjC1AqwIsFJTlohHWs2st6S//HXO
cGw8CEPmU/7N2DEarYBi+ystveco3CiAXe49zzze5CQw93Sp3ZdSFBsgYnwilJjq
vVLeDnXEb9BF+755rTGzwE6Mw17FBAPr0QWRC4W9B0U8PchAeH3IBSdb4LsnE6Fw
VVohJ4n5sP55eagNRsM4XnmEoOOEufJjgkzp7xlx6Q/bPEplM55fGLiZM7BNb4U3
JCrkdw6LNoQzxieFQtjnHvLre3xgzrwWWlfdk9OfhCJPfOmV733WWJ2gy+HhiVh+
TdmoYlwYbiLf9+FG8A8SR2g0qcGaEHXcMuLqS0zUsB0WNTFuc+BwkamCctGyzkLb
M12HRmbPyoy4iF1DfMaovWOB+e60H5Ugtc+bIDUBFPHxEIoXxczGzt8affFaV1Q3
SQaFlm6LM5vahFLnj5GIeA==
`protect END_PROTECTED

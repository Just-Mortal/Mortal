`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXyZBqo+Zxsa9pDrOd4BJbrCjx6JSN3fSUb4T7dm2Mye3KPbqnTFBE4JHAOykfYS
b8cmjt+VP2bkg9gH2NLTKPfpV1RciqWL9MnHEAAoXyHiRazzfLKhTym6yxqBAZUu
SwMTRcSGDHgeAFImMicY9HE2DN9JQFIWHe1au5UCEw1zJLkpI3sr+1CW9ao/hrhU
u1opRvU3S/uBO5nE27U7QqfhRXspl11ciwqlqP1vTGJdTzoSbJQcNLzvX/dUzNhJ
+q+MszsQwfx9l1slpkhAQnKYdNWd9i91+wItPeHn1H/G8ddXlRYEaPqc+giVP0tr
8ca6EW+NbfCl6nj+Yl1slCFwU60sRPOHwEpBOMqx6oDhhG7i6kS2q3riv7fbq7Mv
6aOyyHblBtKOHomSYm2xjLE2SG4bBpKlL1eL5YcdhSFtfuUFEAcdaUQUfBiLkP0X
R6lX4u0hbCkeVYnswUrvIYf1nu/Gcfn2FHnMXd2BxRMva77OO9pj+PQXKoNlLf3k
vkF1fOM1l0SyHD25iRf/e1XlX6NonjxSWZ41u98d5ab84NEqhZJbDUaB+0rBNIDE
K/0DJx//c3MS/AD7nZlXRLmE0iF4hGqAf9UOAwqWQj4sBz4u+Py5FoIHayINR2ec
ZjUfjGUeUKa8mK+UdMMdyr3kObIEDpWr5PyUgkm/sjnJ08Ob1daOQ3EyfwWf2n7J
ntUThLrlO2s9LzhpGcMFcLCIVNsmJ6+Zg5ReRtBBt4kKIqsT1e1hUhY6sjuUB8JZ
vg28XpMVNDjLDtuleFY+E3vpDjEbYFNnKQtR1MAQR44ew6fVhQU60hQcOhJegsNB
jtzKPxCoz7TQNnIh0422Ep+zAwdQJr/PzwduPuip920QBIPwnq2lj6+XThv7bpo4
KHaJUUs9epp0Rgx2Kz//1u5JFVcmr/ek+qcZfGTY8SfPOGTkdCfinh4NXogC29s8
gxiL2if/2x9PN/iYnabfP/2WRuP5m9Q5JagFeNdFO5FdKNwn3msyYWBaGwPzzoca
y86HP5Nt/RJflAGNAwtki92hMeiskYa6FlofjSPoRPrHU88Rejgb0MW0OEALSl2t
61LowM7eHLhw5XyJvZR/2sGt7ITvpKRoRi3KJVcpZ3CUBmg9X4KXhnV6WHvO6tpL
ar74PkIo0xn8Ts+UaQDWqviWGfnzH9QXxOt8nJDfPWAsnZQ1xpS7yWnSpHUeRIny
IAeVAwST1okjUfQ6OzD/F2FZTA2qsP0r1EJ76MELZ9iPwcLAiTYTg66dgNQLhhNZ
vd+AgtKfztYkg7A6BHVgrlTKGKNmy37R0walrJZeeEF3bWBZVYcE5dXAhvbSvxwO
RASXw9j+YvXZgeGjHuSXx6KDVPdGMloW31FIun9ULJDLgRbNpy6WQr/0VFYhhRGO
zMyzRtz6jFT0ob1Rq0kpPZvoqs2G+tAeN6o1c7p4ke+o5iRqLIFytVe7yjntZ2Et
1ltp7lCP2bmcRFe55zBMNniAozYhsS3gFc9+wtUlhxNwDL1++7gTK8151s3hMjDg
q2tO/hY65ngO6ubMGv3BTwfDHjQviz9Njyka59yvaxyxod3quH4EpcQAkDB76WLa
fQmBWtgdQlDgelyFKcNmdDoeQilYeLeRyzYU8PMOu3sobEzS5jprJU3hPpgmdFlE
vPxB2bTH7SrGmTcpx0ZQb68a56gl8eM4AL4zQwaYq3njA8XaveGJAmtxATDJ6ykq
MqIEz/oN9+YLh4onhKO1WaexHmGgR95/TqWNDWZcTZGtFDvoe5uKT80PdYSAj4nn
oKgJXP5+QrYnAUR8jJtsGOAbJwel71Vka49uvZ/2ju72r5rQg8fGnk9rHD7Z6/yt
ypVyEk2Qj60sKT0Q32ZvRkNW/EH1tdaUqcsleiwAttiOJRGLtRI4oZQ5rOPbim7t
IMnTga3z6YbQoquwwgeUzDZJrVgRi134Hxm0b+l3mInj56Lh8PFptTJ4MoH89JfH
bexf42p9kRsxZKdWUrTZNmHEPIqBraU8sMqIj+TVpAg9xhQJmqD8tAq4GwKFECLf
mAnPFzBACoQfrQbClUpxHwmcJYXbj0vzhOb4HH0rR7BDw2tzAemeYU2bHJDiz9B5
l/9soCH5DLT9gcbKC7Dwrs2WWWwO+4eRp9jDP+1+cHmitCO8K87M4s5xn6RyXHZO
u0cf4rA/Pj0Y3eLMVLc6D7DVwf0pL3/36exVKtD8TYMWdxECiQuS+WL530nyBNXK
7D/NZqLUCGh86kzQdR+/jAXv1U/isS5OIAHWmNaaY8JPceCacr/3sUUtheOxLohl
tCD8jRYED+e+wtkV9uwV1784HErKWAhuXXnyhvY7UZ7dSFCsebXXljZdIW/6HSPp
Y6hRpN7AYKtiHp88v3G+mhxlpxHN5yLjUZYMP3oUCXI7oaGfT3V2Cnt5cvYjL9i1
UWcVjOeD+4KNSk+MPen8+dt3yqsgGLeo0eYFqmvHG8fK9txX/8eRIFtpYVnzy1jr
J06R6RAZgUOOyPCBXA3u1oP70ix/qXU4pid9ZVk9/p6R2f5ec3rWhR1spQEgo+bS
UI9swtumZWfryxC8fzaX+2fTd96m9p9x3OPrcMzaSaFY8nQLNir1QMa6GNpzC0nD
mwcrQ52bPX4HAjHMI9I8z9Ec5kIiln/Znml9l79Zxz2y9/gdufV/ByRPm9G8bZ2c
tGTj34bRW4H/zQd1D4bLOkJVvz5ellHeRI+wy3nAwqxKzho+KS0BJKd1/MXBz0nr
PfGmZrzlZCMik+KjGjsZjTUdL9PiXqsibF5jgXwiIOm5ai+ZHo+2S7Uszk4VdYWb
FAALObtcjEsw8A5sBj7VdBlYcWVW9OROVV/HaHER2jsuUja7j+DAEUcTaqH/hDnn
E1m6S5myGf+jTsgUuGiqp4VwPHBUu2N5jrU1tS3vjN5DJ9Jh6tA/fCGM8jkPIO9B
H6M9C+Z6F9IxBFISMyXpS1l1Y1S62FC72aH8tqjsXx2wb7BcCmQmrvBFqyvb/ko0
9q1pd/boq/ltjGoJxztJEk8IEvsouBbSMsIhoDANUF0HKnybkqLY6j5ESHCLVAlN
dPQdz93bxWezin6IJXXVqA9n69ZdsO7H6ILTuxPcCWzpaBwI0/2JtG1AVSNMJo4k
0y3zbzc618hOjmlJGidV1KpKp8gTKQDt5ovA0Mylw2ib1678aq8RZ7C45G7Ge1/Q
lE/A8ta2dG+83lebiqZqMRJq+vqn6ZIhmNUaaXCBPWIwFKNIP/tAmueogno42DXq
PqozzSHDYdRkENwiHdopedcwyg2oDcn+Lp9UhPkopueff/KNA0by2SXdaNwBfsrV
d4Pyyg8mKJ81PbvdintGjUX+Xyo3I8Set3hbqUKNFjS0SgjV8rL/n7lKHjQF/NQ1
KXUOdOwiIDE0obsNg22c5/w4rFh7aw17OyJw+uwLzhL5so03QEaVK67lgq7rPdc0
qAEeC+o4ytRtM+Er4UFMX4tIGZTnEoAbQ9eUiPfAE8t7x59rBaGPj4hCKcBwRmv3
rxgqOiMjsWTu3oWEWk9Q9A3CZG/NaXQmEinz5mSiWp+jPrJ5lCF3VEsjXjkDAEco
4a/CkCodNnY+gMOw9A6x3bRhDZlTp9me/YBz3m6QBXgQ+s48sr1Fq9FzS6WOZGuS
hxE4nOlCXmISnj/XtG5cStatPV6a3t0LaLhMksOQ93RtQJVO2MarrTIFz+kDY5u5
hbQnPFfCv6ILcHcKv1meC3pt1ThnGZoZy1QIzMymig5pjkUKVC5W6QkYDtN/Ok8X
cTG0SLR2asY5DWlVRu4mrsiXB4nZ1x8jCkTvGkhBcrYZRAB2E1AR4/RtjrE1hYRJ
rbu4lbInN9pV0yMRAu7fyDrFfTmW1mQ6rQIHPjZ1PmlOjUq/aoB3A4lYIMYZgyFh
fyPHcQBVqDBsxxxfzbsusKj+bAWVsjLAOtdoNgETJG7K6+t6oi54pzaYF+87Q8Bj
bCikK6bqEbDzDf3FXTxaLxPy9JFFQqsBupeUYxZag3XW7lTHnVdBxsFKrunoA0se
2iM7+c/AJ/zn8mNH6mQZNfBk/hgzszhhwB/6qlGysrZMbcpByuM8jsq6ace7vbaU
807BCLi1Y8P1zqADcoTg0bInvjCoOWNAwq7HgSbvSLvks8LXPYiSxHUuyzy1nJl6
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QmBxMDnKnlDAaA7+ovsywh3f53jAXiGE/7jxpRFO36Fk6CiOr1bQaHsuW3cdbdh2
e9lSHfD5m4mZ/ytd00D47vx6hxlhV/Rk/UGprESL3ag5faKzjZDL8ZdDJnRveVFc
Bftwo4c9OUtukejbjm/jdQOYoM7bdcoJnTJcQaxC7YbjkFcU/k6441xN9bPPN0DQ
G5GGq4jvaK6pG7tMGX5AnTRJfOthIUEQWQx4KGW0afb5h1T8Hj5sMh5GPFOsC67d
EQFOM3raepSomKkBKTwG2Nn/KBHnZFD15oy/H8m4TmrCvD/h3OZ8yx4muZmLKbBl
KCpvJLo1Xj/D2qd017t2z5I3GDETG3ROoWsocKzelOCydcroK90f6qc6J/6SKl3j
1MU82TVTy733RDBvzjAm+IfKs/uVuiE4EGxHamZ5oPxw9te9t0xm+LTIWweZufei
KmCJFivvDRv7CDyVitrYTNoUbtswA9S4Cb4DDmuJ6dfBWUvVIv20LI79Gw0bKhvc
samcgn/bJDxGDX1vfKKg3fnujaEZVGYi5XhgPSpHmBGz29GAPdURVyu7OmbkC7KB
L/FDm5LRUv1M0cqLxIXouqAGfMjBPd+PmJW3AnNZ16YQ/LHXSCEITBr+oVO9wNFH
PGwz85G/Z+iOt4ed5ffadf4FuULcQlAPhDbGTcQPZu5PjkEmCdBYJ63mkjtnTEO3
UjVLkRfjBvIxK8kNFAst9SZNqt0bo1FI4n2u/lVzOWKlKe2chdkdh5yE2l45fj4I
n9eANYXuqZtlRVN5pu4cWXDE+vYeWl8HxHVGKEf2QiVoKY8sUbETQChSqehdcQRI
Jv94MsoRKjNvnAEbBwMkK8XuWcdnPcTka/iPzyePfNsilTKqeRVqYExX4vD2nTIr
GACsgCl1n0xCHZrLGlNgusDyqQaE21FQ3Wy3yK7LkRE641k42yTLRiYRUsL3odqt
rRwXJBZEX3cP+UWleA/Zfvr9vgIc6ceeUTbAC+vgD8jgVHyvuRutVigoPT77kVMz
kBo3cF4GFiEk+/5p7PRBZDWPvZAF9jrvsTaDFoN5uX8vYqbw+l3A4Fpd/uqqU09T
iSHLolnzvVFbsP7pWM43H2y8yDlHfzCamkn/juVl1XKPh3ULMgPO2lUcyzzxYhL4
ihe/Cl9S597K5JYiV2F1huO5Xmqz1fCCpMGb182Hze4AgCPfP1W55HANrUCP+X40
y+HsQe2fTrcLwMS6g2RXNI74mnJlhPJdkvpSyht7SSK4sbvClbt0Cdo0+xBpt136
Y22ljm6O+CSebvMgvJutZHf17zHSNqpsp3Lex3W8/bx3YaKNFdS8ejBJ+wccGUZn
C5rknjfpUOUUja4M+dZY+UrutJgM+4ssFEOkiSJUzchm/OeclODxaLMbKK8Luvww
9mQNmtuD3ZGxU1XuDcs/DHihvzzp7f5xsd9/2xIvYlfdL38sEv7nY+tCyvY0VgW2
qFcJzzxbczZoNj5pEYJ3bg5QKdGxkFMFQ/DEMthox4WOyiMKHyxZKpVjlz3IMFY5
VCU7MM8biEEe/JurNTSgvMDd59/xlK/KSP43LNK9vAaxKmA0DNeUK81tdLKJVk1f
knztSJrEm/NoC9FabxegWqLP8/qAAX7nUsKi1+ekJu5zJH9eOZT95ydHrKhlVeB1
oNDUuNsax7KJ8wUsx09J5eTED+wzOsN1+8ywXNzUzfjY0mGMwrXQoQiGC+Ukfq7f
xBY8CPH6iz01TFVsa+MjMjeVdV5xfOrovJPEJZiT9osk+i9MXIYm6aYQTjJmnfqC
qs7WEVAhBbvVMfFMlpL6h3LuWzl1NUPNYDDrcigifb5xHiv9AXVNx69LamQyFlh5
JRg1Q1PUyilbqwV9QS15EwGPM/Bg8/FKqbmuOo7yN5NI5DdVTJmh1eYdfRpNOcgY
aik9WplkY7VrSU/yRF1vSmLyYSTIDbIpfdC4akHZqqVjy4z5mVJxaKChmHNPTSDC
sa0jNLNYoBA1MWQNiy78BanXAQHGR41fVXMh25CC5P9Ce6lCInrZinqm2Z848ZcQ
DTmnm/Sf0Qb7sHY/dRj10nqhjjnauPICWtZ2Q9s6UCcuzEWgIyfvBWgiijxV4wwD
NC/u1XjVLA2wYGp35CnE4JgKvnpV96BzHOqyvo65M0wzm3ZKYO/VP0euyFM0yJwy
V3cbaXuMyEybsGCIryjHaMKvV/fdBZtRwLmfuD3AFZ0ndprdTXhh1OVpyzzKG380
pzZF+IqnepTzgHHUNQRVfqUuI0PciNuqWTvIX1iCdwZTA22AWLV3iWRu9E0n6eqr
lzwDM1RQ8fm1MKKYi/oxXYDRKrec/L/SqL5zyYUxZZLhb8Qur7l3zJ1+XxsQvPBo
t6kaFwJbJkfda7K4wFAWCzZjKXDxmiM7iEOLrVr9C5IHMuzI9Dv5ZUufzcRKM2UX
D/nEv//DOJYJS9ugBnKtHZP3nvCMM3Co0I94Ia34w949XOGsyA98jWt4BhAj+Oh0
69G7K2ab7e/aKbTa+HeAkrrZwMfb0bdWSaqYI/y+xRlgKppjHZBlOmsDpj7k/PmF
0xmhilRWm5EfRFc1PgABYpV6rRlJRFeNSS8j60Wvjd8CYt6hzFJ4l19ioTYUao50
sZ2z7dH5xepvmuEIXYWO39lHL3kVlFCngqBcybmA6xg50Kp5RSGLWN9LjnLendd7
L2UVOKMYheqAiHXd2E3rD3WjVZYUnUFnG3ieGJckixtLQfd/P2cSA/dnlYNfs5eJ
DF5nEiiGzqHlG8t+G07uQFSB0o8Ijk1onPl8g85N1qR0o3MKaPAhXXpdaasCaUkH
76VSw2wbP4Y7qlkFVEu1qP/xBJvDA/+V+pmLKYS+2Diw3eSGHIzapO7wLqK4ZE76
H14LnVAU9IHxCwC9GcMGCigSCzFhdJosGBqSwncAIf/3o9Yh5DF5mosci49fOeLx
c2bieeFaGCt/fRymFa7l5lhgie+tFJZ6k9+9APnly3sIoWJPklXlrhMePDUJn2GX
RT4W4FR4Uimzxk6cSx1IEs4ahjRUr0AogveoxBPeS58vO/8MVOsAJgh9KEi/yjos
xvzM5s4NxdSrtAR40dnOrOhqFt916Q4gdL137I0B5XsGSBQCa0K2RoYSgbRkKuvW
T9P6dE0wUZuukE0yCED0+QUi6X3wnoVqbWJAm4giC65vSXxheup0jsSuuUynpB/0
0wSQeLq0srXe/LA599u/LcxMTlTylsu9IdUG1aDp6yseumEpB5ZQI6JHoBLFZdmw
TPdv1+pbLwiaThfXSiWDWIbJpGvBBb12g15bD61/2c5vvFBpt2YCSD6ydzjB1U3d
yl/FMj7t+trietS9zw4z4wVwyimDa/s/mK7HdGj0nI8UBs3/DI/oaqCSc9cXNnG8
/eL3TztBRHnJDvqqyNfTvRRukFhBPEv/7dAvE0zE0r5C1CYTfaWIawL+MO+p6ocI
Tqw7eHy8tRHfD6Xe9hcHuXFAZVJcWdNlq4yUEsHxq4K3vKpTps3CZgNboJUO5mEa
V9ZPwbYfap+2dfZaP7oTt8zuRcprMr3xzCMQDis5zDDn8bYHGlKIBXbvS1/m46e6
UJjEgonkLV8IX+enKcr6nvtMFVKtu+MQunvU+LCgQw6/AJyqm2SBZbn05GzhH6RB
JenTLJIPYUDO2Yswv6QOI1DVqPAD1xWE+mRHacbkYXyMzCl4wLa3hgIU93U4etKs
N1MehESTL9mXKFVbF/BItzR2PxiBHdaXmqL3Fw45tqCTmbpz7PId4faorm9yXIqO
Kh92YvZ+94EPjRbVjBQDX6Q7j8c/pCoSr77cVT7obkrzg033ofKkCyiqbWYUaniv
lg4anXnn35mUcHXV3qZ0Os3oirhGiAoiXBqXNXPt8yWBc/g4VI7Kt94V2RT2yzxY
ZL6doWvTshrBKDiOylL0h/U6vCnpqP29ShKnazsOkR8vVwdX87w7be+apdzNWCxF
U8+v/Lg2l3ss7Gvgqlx0tphLlbHymETxxk1fsI3FbkoDgzZUjY8p93p9cVpW5Agr
f/AwzUlk8v9+8fdikgFLmKurKBzaTY/+Cdf8vmekacJU9/ISvIj1E77uo6p+PTdC
pbGQv7DjtIPAz1klKR9x8Poi14qpZQySq/AV/QrFiZ/492jM2XRGo4z9+S3GDFL6
U38aqNGtrEfOFcAID4JwEgckfcz+FUmTpJhXUPHaGjVu40vxcEsE9oQqmVOT85hE
GVwhpOb+aPPpUdL6D8IhNFP9MK3y5CXgVGkkwugPNYKAExqFHHjGKYKhDws9/K06
Gnta5fk55QpMQE/bnepyAeZdNWaQ0l/cpy7bMSSCgc6m12uxyNxr/8SBxw/TSp7J
jW33oP1i8CrVnvh+5hOE3ujZwxqszIK41FyEUf3OnLM=
`protect END_PROTECTED

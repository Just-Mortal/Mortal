`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cfMYSDJj0TUqxbDReQLiUR9o+S31EP1SMHv0WtftVq9rYNro1Zg417kU23x0dwzy
2Omvul7QA1F34v3wM+LNK689UMi6j2jBzwhkWPPmxsZNDYkxLR1z1BSEwwo/04PY
td+trF3bvBaPZ6i8XXAo7saFYqeK5ZJRvwISH3756PfhiO7a597H2nZk710FPlpV
H6O08adOisg4n/gzJDxx89gkRHCA0OS2EQ5lXWTHfM2f5bvtKL3m3NH0XyiSsqG2
G5jhXqoSC2KGiFRoksWtsC/nthgseFmfnZUs+wjnxzbW+Im1fLWqcV7kAp1A37X5
auYHMAblBU0mGrMPXhB/LlW765HgRp/Z2HPevyB3tr0=
`protect END_PROTECTED

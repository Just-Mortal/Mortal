`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYzsxmBRDDUNKveVDzpKG4AMf1uaE/kJ/79+gR9yPsX6IDTzQxQ+AQVT/u2o7p9M
K/vOBtVQt+bM3AHz8WlwBCWWLjvxoCdWJqxlGF7t0zWvddO87+AWrGIuS9mHq6dT
Rv1xMcuoY9KByi/3dIzFILIKbvgTEyIHoo+rsrjQl0i+9PncrkCcMOLZYuuQ4L95
me+j5LjweHp+y/MqVh9qoyV1jnC6ag/nwPtPByvGEPdQx8PgkVwnKyUH4q2smCVA
FGEuBAiPDo9jsLlRD90TWF2ZfGiZ3tPaesco4uwBMIAwIQXw4ovY0hCrIJzcz2Gk
tFsfFseOg0S6E0jNhswCVE9t/RZd71kuSfETWrO4zedvIOpzD8dde7czF4vFTZVd
kuZZSku+4IIB6xczH4oXUV5kYV2w3sOmi+juNwpw5084SmoVdHf4RmFabYl1Ut1O
HSjRohbzn0h/37x5FlAYOHYsQIF4Pd/rcD3LRnN8wpzbm1M4wtynWOnATZMtINsu
b50Z+zzm0mPXv1veC0xK50GSPTAYxrgxfjGYBKg3URy4vYWwDwpqpDTWd/Rl0Cxk
nbifhfqNWJ34+FESA6ybHlg8eA/CagfRlGFU+cTcuF55Ugo5XOGfy+hXI2K1ePwg
jUs81jdztUxrQWZahdaNFa2RS9i8CqzhFAHHGNjlAsDBC8+hIUr1UUWvjUDnHXgV
Wt1bvuhG1k2bdqCYVXgxnsAT6Owif614s0zf9Q7y1eO3xraVL45PpUrILqwJOM0b
+djAS1VOt0Em0ipqHwOaIqWrQn1Et3RuRe7ds2F1HpyZGVO+j6LzfQKHdbuMtiRN
MjO7F7cY8hSQD4JvjHwB1Du+wOdV+2eYNjdYwbR29iZ3+XosuDL3f2PZl9SEJqX9
kYJh3xGGcNpDB8lhuuGsIpw3y5dJQyilNB3sKlMt8Pnmlj+08wbTCuaX/NjCD6uN
pd6X6lB/6qDuqOAYDOpAvwFi4OFLcM6pJcP+ok3QHQYnx6CVfaZJK9uFSZFxGbMZ
R71GbaaHVX4x9PIO8d0oQ+MQsKlU3ldC2vv8TKNWBnuDc4114ymPrhrFEEc8ajS5
/pXgOK/Tfj55HpMI6I09eFM4SNPHXBiecZogbIIG8jHXlLZW2hceeV9dHGOmf7uc
CWxc6LbWcOv5QQGzgIv3SsAB8SvpxOS9SKHYLSXa8kU87/GJVlJdXbC2SIGd3dnC
MFYX9JcLlgVAmxGDkhYIDlz3HNodQ2zWemqg6nmU2w/DF6AoJYUuqPDZSAwbxWED
hrmBEmrmUYzmtCLran+l9AHu4t+Z+p1Am30KhLS5IQNDsEBZi0gbvORFiy9gCBXX
wP7XeFkTU/WXM+PYdc7ndanvOk0ZntWzy/PLYl3NfOW+tKSFQWmyA26cOdst/hqO
J7Dk9TYONmnNDSCapIxz7GmbNo0w/zdl8ivpGS0cb08r4DvtwUoCb3lB4GUaM52G
ax8+SpIAeoDWqIseW2N9WldR2HWANl8JlCYxBMPr/+P2r5LIro0JnyMooH/dqi2E
FERJKfvPbfReksers8F3aDaBXUaSS8lk/Jzt+YpDXR6xsulNhgdOgJBzKdtwceX4
rjgeNP5+nQQJSsdhB05C7H93hpU8YxAI/dSsNIwrUkHqHZ0PxCbTOOtZNAJENiBG
B93b6FTK3Iq29sFW+yQ6Clddk7oQ5r4Mfd1grSqXH8i05S7tXqd6uXzDfC9o2j5v
YxfDDWdl7aTUHMTT+j15WYglPGsz8CMQkdguBKiKOYqm//V62onEfrIoG2pjea0s
kESstOEmsshEqnSufKF/rvb1HcQYLX9nhBHjOgPGXuELaDRpl9E/n07d+2wcJbBH
d27r6KRC29f/4bCe5qF9ttIha51mgo8pGIsT7KNuxSEJgJxWk/eQXDGC2yiN/rNY
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCYnyHbtUm9X8JpVSGWnzBkA5aMvqmfSJYtMBSkD9YN/oAsENiGJc/gaxx7tpRkH
n0p191PWwYqzvWRvMSivVLNBxelefuhXXmULi/f/boNOnIxzrxAkL9BzQN/ojHyY
26HeVTrA4rnN2D7MgDigQ0BxUnm/X1iu+ji26+xSDUwtSOxrt1+tbLAlzQppaYwl
pIyGeEfAnb+RLoNpB05Bry4FyoayNQMpD5Fd4bfh/T0EEAeqGtTnvoO2emyUGCEb
vyyXBDdsbcEM0QeTQzVA+LVhjLjpWPQx6k8JDEYAWBPWo9ARi2qlYswzMjL6+iwa
z9IIkeBIqd/esYp7tuJSppH6oKW0+diyeruxRR7AaPsswoh1VTM+I3UfW0oLUzM7
u0ox/eYPp1cxxdncqzYLjQ56XwK+mgblDa1cZ3IHvVJKHTAAgjpVSoh/SPEyTB80
5ALaMAsAgRi5DvF6VYkXLXDZlMv47U/28rmhE4FQ1h89qaFSxb/6EsJR5iubuuTO
F2U/uMj3y42Tm8QpAI39/9gVmFbMEKVjr6iXM4iYu8Vf+YyFdJtVdu43pCWLX0H9
Xr7B2rVczSwXKFn8XqzCNg==
`protect END_PROTECTED

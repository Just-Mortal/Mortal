`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
slLTieVOz3SEntTs52pfJZQtmxdGg/8mQ6sIrwdtGgRmBYgCqydVIMkBPHo2v5uC
DvPBAktjF0YiWsjXZxpbFoQ0x7AnytkVZ6nJfQyv90MimF4g2h24v+Bgz8SsaNa/
BmANi2nO6XBM6vFqLhRu1hnEz1QBEv8Q7tT5RMiFROCRnKdqYD54jUDYBX9PBT45
wvmFUp9eVnMDvoAwy20Q3A7Cx1lOCs2Kmk43QyVuTxPHjRtc1vad645xFnU+p/Vy
E145brHNrKILy+zzc/O+3L0idS46Wn2Er/ks2YoQaT8BROoS0yGbDp4sTsG9BgXM
ArrJfaD3bKW+P7Xg5UvCRvVUjaCHen9wDy1o3wHSfZAADevKBJsXdurl6x6RrY66
j53XP3/F+jZOHSLbkQ/fvq7hNePYHEmdet1J929c2MFucmIvhaNMtBbttObao0Pw
RKcLX3QfYHix9ScCnRRgVIahrt+Fmhalr6lHTqNqzwg4I4eaux/5r+qesdsOjtHc
lVunxCgP+zrWBWzz3yVOH07UjNqocFZzmeNWOBQD+QEaOoTyiLBsnEuYJCoLw9Tn
PAKQi77KE+Uz/fje8IRb/ZODDUfDeFu2vVXTkSseF6MyDeZTy8/cLiD9J97NHpko
2hvKrTegaDQslvudxmI/Qhq1Ma3gHjWDXkjjR4bU9V0u8z1GCkb6uY7vwOwFxRL1
Sn5tixK+3DYXgUecUGVru6fHgnZfNeHQQ+TTGLmBpMMbZyyV6o8LejfN4VLDDn+t
oKmMNypeWBQwrsCwY56gE1OHKrv1/mSHELq0HIbM3NHYwawwErTRKGy9sB76RcwP
+BQMx6nDWBxqqTVAde+n3SAWG90Iby5PDNqP4oLDIJRW8uEhkcjyyfmgY4adyrcl
M8qMBkLKmpJAbLvWC5s0I5aOmkBnPBoBrM/Hcv0KEzzCIZeuWCXlHnGOnHvEwlRx
W5XlaQxIfRPLPSbihKRoLMpTlCLzOFwxa3fk+8mOyfFQlSN8tnJNdR3NeyR2ICD9
Zca/J7/e9Mo8peeXIllxNBjJ3q+C0kIM/c+vTnStcn7ASRWJA5FC9CD7NAVnF7eY
LfotsjROd7tm4AGiPH7m4xcqjc4yI9jOWO6w8nMkb0OvTjx+qFUMyYy8b9xssndc
zZ7G3n/7PFV2cHty9Y8Q/fVF/l/bjwgbndkSYKm8qNky6zJAW/77vioJQPX5DwP2
L+S6lRFBHjQK59MI3bZs+h1EZPEzk7sQSKuFc+SjtamtOSYeDxQ3LFkYpOs7z7in
Ql6lXkubchqUOBzEgUzXsHwO7tDyc+sBZ4EBnAQQG8UiUugqhafs8Uz+qnKXza1l
2tBsspyS6qGNJ9Oy4vyByPyOEC46c1p/ayvEcivCi47Jf849i14yuMLClaTQnLLL
4wM+drSRIMuqJgV4eTAVDZkWJW8SLO18jgWOK0BoxQZAaq0t4yRhWIZ3j1FOdyzZ
a3G5v2+yOgpcYvNKzlEz1sg2glvwo36m9JPdIuCvGg3q9VtU12Wtyv1jJUMlAibX
I2ewV8NKXUa/M4jd2h1OyujFlx7X+OO06glbh7zTsePe2POb95Q08UKlmhbNhJTj
BT3MjZp2UKZrNNApBqe6hb/lHCm0ktanrGga4uxqRDTxrV9uF0VyVTRC0wefpR5X
qgBgMrLNWwEj++vjnIKQbir5/QWkbGLH/cngudhq3mDUMYYU0F0scFPsNE5SG6fo
rMZh6loWkATRQ+94bvyQQZCfDc7jQHII9PY45iLfLZPCJegYvoxt41M2sv1ET7hd
fs7fVoZgvG7dZTcxuRPvFqWU6I5tw48pkD8HoJiYzkwaOL+ny+s5VNvTmLxZncL9
qCON74UJFQ1Z2oHYlX2t0xAvMeIlwl566Y6tbJ75bH0QmG92lfM1UXd+T+jA0sr9
WK21oIdRUiKzFHSwgQfcUUyuOl5woMzaUIHGZQuy+dsnuCJo2vINxzqfilznqJYg
2ANGygWN2Iv2/sNsSNVYI4BbD2ScgdzbvyXaK79Na4pkAB0m/y02HA8DcFnufrRs
NPjWvkgKOzvKs2e8OgSalPltWo6AgzS702/wWiEcEUKUixu3SV7QEmlzsmdA2jVd
upVhL45r+nRlC9rBDkkTPNwWFBn5hk9+t0OYUWALxyaW/Tl1fBPh/YMoMVMdtc7u
rdnyeoGaw0t1iT6l/0xDZyuuOjwH4p6uI79r/XQ9OyQ2XQyaV8+g9NX8KjzMRtU8
K1mWb77AgsDS++H65YbmeMGckCZ22hNaeIlgTisMZwbp3XM8DzBKrychagR4pNjs
+6RODinekZQUXs5LgPtnE88iyrLuQnGHU2Kw6niU/6wBG4yVBuJY9IvTEhANH69G
P3uPIFPUDUPewpH54sby8S/DWLeDniMwU0MBrM6QETHWadLopJWP7wlQsJCFu1ND
8Eyw5lFZHq+mdlXOYD9PidsO3/oy2OSoWLH5NksyLar82x3w1ImDcM+xrn3ErQTR
tOitE0Ca66yNwG7vTJqmp4CxcJNj0WdOx9Fuw5fzG8IpfPw4RNWBnrzHEv0ACtp/
/vdWzBzsgmL28t2cgNKGUhfESn3lq9ivhCE0APWzaNs=
`protect END_PROTECTED

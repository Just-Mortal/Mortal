`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k2LQGVqbbzsDfT2oYcgHPIopv5lD7cPlEHwqIl3vyuUOKnX7Thoqmw/3ATSaEUpT
vc1b2xIJKHr/JIObU+EUyH2LuCf0hgRiam4cLAjy8DnI0HLVV2QCdBDI46IKQpQy
vy9kY9oMkCc5WSR5uHWNCNndkbtRX7PARSqM58KYcqlW+/2HSlz6vHu3G6PqLKsI
xjaojA5MsxWMBSN0tBuRWypcu+Sl/ehTtvxn2jS9unAp5mdaH8JiqWy/a/VgC/WR
P1ydhm+euQJRbhegaYR5x8hRC98ypu6ZjXrM8BPblid70qHsC6UsX4XIkZyp+Pma
2xNfwmXzlIVE73bwSTwIxMr2LZ0i84lxQ+P01FURFujRrJjZzOXvjF4kx35nS5H3
sUrsqY7GlooQqlWIdah0B50JyxGr9IgqxuBvI3/2BXWxbP/OaQ0XwQUVqDy4Xev0
6l0kMk0wQAh1xeif5n+nOFGGFnEqL5LBu1Dmw9v+BoefUH3W2RFfJG+ga3OFMza5
ZKOA2lx3FzRlU0U+3jqB6i3mlzgyjAIanpk66FE0i70nKEz1hS2Hbr6/ZSZQF+eW
gKKFenZwZ1vTJFr561wYY5jEM9bdp13rXq/OSM9S7uAQ9+TL+Venf653PLuRaIQG
STRIfj0IqqHIS6celAfPTfuDF63PLCdw0H71PV6gT1leHZtMFXgXu6iZoc5yedOd
Z48kQj3sMBpgE2uDey5QPCiVzPubdIcoZHyTptseb9AF1f5wcDzESRkJ4Aa1jRKG
vhafip7ntFQSYMmVeBul9VRWAhPhZBBIqEsQ/ElJrJsikKe0bR9jy6+1nb5F4iml
qnX0r9sdmqIL6ViVT0mQ6YRWFoN1KTVnX2RDWjYwfBtV78aVXmsUlemmaRXHwK2v
Ff8RBWbXzxJLIHkkEZTp04eaJjnvsls8Au75apm9rDRC4S5AEvoEyZcIS7Hd2FU9
VTvJyqJftLcnGXpMdQuubaC4J9BrTO0YTZwlz3SNcANFEkfo+HOYffS+lS2yy7cF
yLPBv9T8SyzocjuiuYIG4tXHPG8yqwmqz/+4E4gquwNnPY0kzvvoJ6xrc5ozq3PJ
PCZbXw/LKnubxSj9YpsmuZ8py7buicR5Lac/1RNcg48lx/XIim58jR1bKmkbKqVP
cqtH04prphgptA0YxQpuQ+9/uVKrRmMvkqsx0r2zIgKEt8FF2NBGTtSVWSz+zZSt
eLRd4vMnf6aX9XUxou48bXZCj7hUAFJN/4Vr49RiWbJYrLlX+doJrpvDa0bsS8vM
Ni1BUbc1Nvmpn5i/QguGlOlmi8YAP0trRkKoOQLfuDQkifLCR+m0LQmY6ixHAurJ
Xr0koI39AtHNQJMWMADZkLW+uNZduTOMxSNITRglC9ZEtHoT9YXbQlC3BxEnLVmJ
DedWuYAdR9FH3jiAWwTeEoeEAM9v3u1S5/6E4OBqqveapxlJL8CqiduKTbHZ8pXG
yuiHcEwNOOwNFuMK475lZgvoPzJryFV6jP35t5jOuB+/bbCbr8iFyejZLihlviFH
kPR4S38KjaenLIabVsbqts0014YOYiQjtqdt17FFeeCx77Nc+2Ni1Yu2Wgh6aiBq
/V+ZfNdmx97Kxq773Zk2eSjD/bxQzavdKeey+PrHGza09ab8ZOOtICw3jkl2PNHU
R9H404X/LXe2eEkhVMvbtjXMeLOyusy41Lwmisz2WdDKU/D+a5E6pEvLocuVlOxU
RVkr2kdCQ6Wz88Cj7QTzHC6pSyHNiHl42uaW8QgpWzgLwn5bZL0//5XSWU3Yhb2x
xTYmftSh/r0sVAh/BsMPMENc+Z4hwHk2723G53FtiFy4yEPHqe+Q/eF3RUtYMpF+
NcjIHh7AtIaqa783+ZGExslb9fv1CKIOi3y7iT1BGOzAhs05Gv8PvQxrLIoqkT4r
k3JeAILfojVKFm9TBDacBzX/I9J41moNpaCiUDySemsD/nf6zCzXv6sYo+U3zXp8
Y/RwHy1cl/Ank6zLbngyB1QBlqxsFRo5algd1g3tLh8ydzjnMTlfISNOvxs4ubhH
/N0tgXWddC/IsBsfAUC2f2qt1KOuf2qqZThDuYAphKwsJ7K9kGA1iSF+LsX7SVtF
w2j6u7h430/q/V3iJD/u3Pmd228zs+Om3oMyZnOO9LxvN34B2bS/kB4RvAUYiB7w
dVpwy9F0lnbG2i9lZIanUKfmRrsm6q1XLZ2R+/xn16HteUZEs3vhunHSlRx79yfn
XvZSzCdJTfXov2S+4HVNb7yl+RGXf+nnx/4Y1E4ewydLCI/AFo++kSX2hMSb3hdf
O7U9ih2S0yb/ugcvineJ2DJFr3rToS/dYUIOBcKjWCn9udcg6QgMrOkeGqssq8pJ
EuP99twy4YORMxZ3tuv6hf/hVx5uNMFGUGtulqU3vd9hm/WmpoeuF2W+29JPUl0J
I3K6IT4Ji7Pp+D5ctD0GVfkWYmslNcKvGFPnU3eNhemAApCtc2OgBpzeAOevG8IG
DspT+1oUK+1gYkfHXRqpxEwbkOlHGtCFt7rvaUr2OEKpgcRNmkos3SkP9wmDgWQd
urCZ9Uw3PXY0oTGaGloqg04YkCntiVuqNBOHG/+sCKSZKkPbEUTeuNbUU2W2cm+i
bEcwmTXlYZaL9ilL9XJQbv6ncopFoHp6AVn+sqBtFJI5aJK70kp8ivSPuYBBo7em
eer8GjPZP01+qRMFEBQdu1GLappxKY4QikA5a5I8Zx9BWHAKI8fF1J491aUlkMsF
pQeH6uW31OyZvzo8RAf15kgM0GvSLaPdhiQSTWB5gHamWSHojhSTfym+JuVmM0Bs
tmArE2JSn2xTMCMh+O8yxH2Ti8t8fWeEZgLaTXXc6P4s4JSJcksgtq5hX17w+6Dp
4lmOnQYIAWdFznnCZ1ShtQRAf6b0cuuHSnjW0w9pcb6VV/Exy5Dfsu930nhAtnwr
AwF1EJUUMaJhRbFx9iVf4ZmTWTUfZguSz/3FsBXon3pXz9hOqGfjN29dkAQaTZWg
sHSqZvKhoyljWWbRZq/ndN1Tj7tqDQNGHARBWUWVLZFgJkNn0NmkQK62ZF76gLX5
V3scoPFszPf10DWgLx5+bW62+TA9TMno15o2kCK1kuLYSs6j9/6DFaYaX3Szv8ym
VuXzTjOZL27FWfbH5CTr0V8S3JClsSjWkdKyhts537j5IJokmNEtBHQMyjUhW5iR
BAIi9sRjp8PKvb6gJ7WbOLspN6V7dOPek8qj1riFq7xlLXUi2CylFBH8JmQ6sULe
IeQfTi0gyv20i+lJ5U6zdKGMLB178WB9qvpTQ7NurehC+nbw3We1FJmuNWHxgwW+
Nrlc0rbgaMtYlLxw98llfjR60EQ7z1vOW4sEdi7IGPAeUT5IzbbHpEsIhJI8OMv/
2pdRtj/xDRRigxl1xk+O5FTNcWjX9lzR+VCQnRYGbsaBEB4LQsmgA+C+3RlF5x2n
o/Z05ROUcWjrQyl4Mic7tRZCYHy+oJnXWssbLCkDpksV9mjCfcE05irqGChRb/s1
d9PvfOl/PoRzP1YP56v/LLB/Hlo1PqcqAI4/A0kmf+6eMYuH6bprWUHCNAmTQlGZ
jJq7QIQapx2Kk2xZsbUERLAE/hT1nNi+uNt8gFh0aMqBor8y+W1yotxUqS0JSskL
o/VdFwX9QIegIkynfosPusaj5IYMDD/0SKn4nXB3G/8cFRWeq5qANmPeEivlHq4G
C0Hq33aDkZFTXYhvckUFhzNzDIKTrKolC2Z7Adc/jDDvsu+/8dqLKeYQqDFriy7G
5tNtrcrKcpImmGPQIDuHddctTvCSyGUJtA2JC4JkD9MhgX0X2G6b1GcZ2s985E0z
re82+GQZAypBjt5vsfs9BY6GgtK250bd1dClrjm6XaLMMB8OC8UGBqwOI+ETA8GT
pTNNoemY9MXR/aDv6nETYyzfiivq7t/HNs3eU87wH9Y+ugs/vhPyc0KPmOpc+7zE
l6xCHgRH9bdYy9XO7DaYMqtXB+fh+sO/1M6qDKEwnBg2wiEvj4eLY0xXGhsjNvOv
9xaTPAKv/9m/qTv7ogrzmQSUzqd3VanSnfTtrEEJpZ8TrVS4wXsld4ZtGGlSLQ3s
/jpbTMNKfiv6gBltb9wVpqJMlGxsQqAncsGsfIXk8X30RkVgEcDU6QU18UC8Os6/
e3QGFWggTuT5/o04OSZFqyHKwJUFZ9W2PSwEvxiLsoFJxpuEzdT5jK1impub/Rd2
LaA1yqauIbNbtoAk0UczRZ4n+gfrd0FZBgOSXy5uyuB782vHRxxXRQHCnpFke0UB
ldxMgxtzwM2vXoTo0SxV23pn+2wpz+2OBxO53aP39ztOS8EKYdXl0s16Q4/iSIgT
D+ofrxZAeZsc6JK9mkKtF7gBZSEtTYqZCrNHD3aRzZc=
`protect END_PROTECTED

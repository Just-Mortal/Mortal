`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
doK/b6yKLGAz+OctO5tyR53Smgnt02NzkYqEswLHeH6WG7H54vEwJhSKOS9KBKdx
7nykbNB8zboPa6svzsKxHHoTdXznbOSkNSnVo3MxSjxjzC5b5bpAc47MiRLHJA7q
vkuYv0qxarb/qaNSjuJy6QYkWzwqd5pYnmRSeeh0q5hYzNmqCH35gHmTPBfTskgf
FCvMgCARaZ3OS32dmw6TJQdEQe/WVtTFHfgQnwB+RVZPFIZTLRK2i/l83IbEpyYy
JJ7jGOR5nLGEWEfx8rUGLkfKDXxO+bYn/WXcL5L1z8kPZOaIcQHKsDbBi2z3/cMO
Ah00m/0+DxlxMII778alZVrpefO4V8iDI2CSgx62VYhhoj62SiLzjlwcukEFd1vV
Cpb7RKzVjdRhbwos47OfJgfRJT9QRwmrGBxAuw6Js5k7zeJtgerMlsETg14i5e6l
j1Dqe9Dbv/6S3p3IyMS2eAwrCiYVDBxLyuSPDOq8CP4zLV6HnYBz7O1LTip1fIPM
TvK4hn9Fd0JwlvB8fgdQqJ+0sNOiDbnykFvWmdIw77uWNYRwCWW+1FQKBMNBbYTA
cHPooEj77JaIhHYlPk8GsJXYm+YvVpRwPhyn6sO88tWiMUU52xO+0HI6YPo8Y2nG
ktBJrBHXus5zNP5F2hw3TQN9zq7hwxiTTnBKtTdsu7ZqMwkMa9Vzz53Hl4fzrMwP
eFipgwf0G2oyy5d7dK8CNh0m1jPbkc+mS4o1rqfdt6d3bvUowPUQ4sqbF6vbMMXw
iifuI1fihtVhqUY5WI5VnYVRL+AjeKppF1ucBGIHLosspGS3l3a6OcTiARswEilP
zvmuo4oIIsrhDExTEeO+nu5KYF16ivyVzaal32VbUS4oeKdJ+sDkRFrT94MfeH0W
j2lP3gGvsPJYfRr4oLOEoPXbeERgK4bnWhNHjIiV/yfywkh7dcQ/QcaDtOs0aQ+l
/CJopGwCPaba2UsCSpgj73XkDZmDsouYCkxf7dKZ/72ZKTa375H1rxg/y4wFOkgu
N+lzj/sfbNOr2NcVZ/uAFQlpkNHnEjGJFJ8v8PAgexN5rOkmKDs8JIzMquhXKW5Z
wwFJEr8HZ1YzezmtN8asKifpiupPOVD1y+2PXLdSFLHQqTkbGiokyoQRkRx/gXBi
G961rOPndFQ6JhQK0ebIr22QQi7SwdD74IxQkkPUo2FeHn6Joze9WqWLKkC2NM4H
545isFQd7y81Is+FwU/sclt+mV07WCEfurs+mqVXF494cFRycT8VNyMuMcBD2ynY
q3l/R/ynH/QFj8uFywdMURpLP2+V24ywPFFJTar518S/NteqdJTv5UwoAJVMEGT4
ivaTWOPwM60bKI3uoF0xC1zskl1spa/xtVe3QkJaOWAyJyt2T8uIfx5Fk8bJRlep
v0TraK90BiPgA9f7GSX9lIzxPfIVBzSGfHcmyla4iDm6eScTyIuHgr8a19T9AvFa
iaGGF001U6ZzFjAb9B4nnJ72tlO0kT2z1w2bSAp8Naf8jdcpiDLPWWkZayAs+83V
6FQV2n0E7Bv+jFyhkcUOEAYzMlMrNFad8TATDAaJ/1eYdLOswuR8bWdUBobx03oz
Zykd7Qu5oCbqTqqLZjaLw0omflWd2pCisKeCC0IkUNsB4Qg8g+0Hujy3oskGhm/q
fnLeyjfR9eorr1KL4fhjKOM1Y3Xbsm15MFtYC6ydla7LN3egFo2oQiwOAw3BgOk9
mpP3Z25Ib/x5OTte9+xzrfdO719s6lPPsLyk9gnisLEkl6PYL+NYItzVeZc5Asne
+FNovR1N/gA/2cYECw+eudy+KVncQKjn3PnUWiSRBt5gvRdaubeBQ0onRKflKk7n
lfFHJA7SooOOjYvziIbmqzrLl0jxG1FR7SPAESmegY3aPQrHUGu9DB39S1jAfkDP
MOouzfAyxgxAEuQHDQ4KEyKX+LrswsjEWMTAsKshEiyb8mbBmtL8p0yMgwPA0xmj
KCSkB6DcfdL1MvSisFyODHXRGMjTR2i8jwZSK4bddZbnoNbwvHj9jRPC+5QBQjj1
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqkVGuFXZ02muDC4xQ5ZxQl2r24iu4sPZHperLD8WPf6qNIlcScq2X+WLIEPhZWU
ItVB2vXIgpL3ojzFSXO0/aawXS0ifuBkjFV+5JGgqN8+1mQ1ddE6y2fB0yyTME9V
K0mPbwu170d/FP7dFoON53GgVqjZ/ORd9nIxRD20IxAM+/Yw4qV1OH8YCsf5T7ot
wx0VfZ6fdmiNbl6vvCki+zf4BNdX0CSGpjOsnjab4ZIqa8pncz0VS3EfhChl2H0A
d0fEYz0JmmL34VfjNZn1bPiHrSFPBoH9c4rI5bMpZVMjd8+XFjrkR45w+eZOSOXf
N1bakpjd7w377NpcEVNrr59zhcjWoPQjmibC16uRBkfmioECU8KgygX6DSRSC/gd
/0r6TFBMvIxQ1GQ8RMyMqdfivo/M9CILzCYr3rI0msDAuzS6mrNxJl6rFeBrcCGT
BqqfW5lIGoeKC64urdfhi+qMbveOf7dvi2whCYwIuCNnWmwXBFEV+oiDxhziIhPN
6SDKadr42ocMNgzDm4GgzNGlEJYQvD+dWqOmdZF+37RsHJGqvU5lPkOTRgpKgY6v
NjqOhASq8NENc4DQFUlKMwfQctzoDz/ea5EVzPwhO6ME1VNGl0m36cPmxy3p+fYH
YmLy7KRoVi3+chyZS6goRTovsRdAWxhGYf4FwSU1VWmBzHsUMe12CpOgF0RDbm5M
fZqbXpgtgvegEAKioTIfXae0METQ2XA+oI31OsTFtqr3jDH3PbLz8rhOFRQpqpD4
LUdZB8xDBAhWSstl1plZBwbU72sPE+MVr9c+PLX4rVrWnoR7nT90sHatZmvbTg7p
hv7/DII9siS+3dbqazr/8y3MIMhM6XEr7k2XqvD7ILlsuJu0KFvVl914WfTOJN1t
yFwqtdfhUbfASYzRf5RAFKGim2hQhYc1XUW/iEQcpRs/YV9+Ot73jQhnyfJgC/8R
gsVb1goVOxl3ZMIKhb38RmBWmdRIp5EQdpMlAXurveb/It/1kUkgQit9V58P+P7R
d4ec17u73eu7T3sR27nMkmaVGY8NWY7EYnV3KqQ4yzvqouFyYPdRMSMnctyqli/L
vrgLzMPibKrRkWpjuP9o6u1bjKKDl3lV3r0knix3S5m8vdbOKcJ8kxlMmW660cN6
kO7eRH7IUO/kRcSP3lhT647ajkiSKW59WvpzOfhwgNfYzw8U577ivxI8I9tbuV3w
quw3920F34hgxqwqzy5gHGizVzb1QPPIN8L3KzqNHHruXfvdjwuiRr/3xzncvjh8
Yvdo8Kn0kTGVIugBQpyeRqENc9gsmmB6aipH3VI9dQ6tyoglOQy1ZPRU3cQc6qf3
FVh2pb/XbMS47UH0W9KbKB5d/Agoj3wsm4bkksLfJ60BpkEUfhXEbBuiMt+rs9PO
yflY1dJjD4zBlyfQnXYXRr3z0gCTLc5Ssi5MyDTlGRkK4vzqxOFsDBt7iTOoslBt
9G5Ns0GQSEkWxfR/LdpRYpexQMXjxnXLdkbwT4sysrYC81Bxab/AHErEd8AEs27n
WIX2cDzt0aAJOkQFfvs8T1XGkQbQ9CFcWxfRNNPCikV1jT1IEVo6wplG5gUw1zi3
jEXVdscLVQsyfsJdHx5Y9ODtHTS1Evx8HJdgsBordXTgM6+3AmO7TokXIuXsJEY6
avSiJLBzjkRRA/cfXBqVlOq9nxa1hlGj9n0MRhOa+gVHDuFdzRuc1ilhjd7C2mlx
0YAYxqdYpEXvFJDQQKtiX+04I/5/Pe6pFPSMkxeJYoG8IVBoxKGkF57fs7D8vin6
tsyjUVrtcBRkg5N3bMYfJH3jz8ytJG2V4KFMALsiXbX913CmHtdCwTJh6XBRELQz
K0fVw5a74aS0KKS6BTKiN+NqG0ULNm4G4fK55RNvC1ZRCtJXz/PzMi0ajPK+BZ+y
kAHOWF8hWnelqwpG5RPS4M39O/XjOcwEDzSy5O8crigsmtXMHskP0xW0IZ/Z6nck
eahVGzW5RA3RG3YPmEQ13/Z4Bz3S7I2w9Ycqh4tncWc3HtDJujWG4NnN0CnROJVe
d+syOVm8PpGDzufsQEEV+vILXFo2tK2hW2Kf4ZaMbbqpyxIg44jGkSK7kfVEj3a6
4ZYnnO35ZPTFQf4AqDJZux6hqjOMo/2T5tIXfee24F4TAI4kq/JjwVSaV1IGjTrr
2+9oWEOy7liQ7WAcXCJVk6RRDJsTxL9pQGxpI3odnDc=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mnwDPSOdKcJHdyR5hSsKjBfVJQbK3JODq+rILFJCZjDx8L6xxTTTz+9iWhQOWo2v
agWtc8O6Q9OlEFOVIRQMLa9DN68n24PwAIIgDFZRgNy0GEcFhL+EvOb5OJ22aWqE
jHFc0fNUzFB5gz27tL4H/jtW1lUmac+tZb2xO8hEZR3nUsxHsHPqUijIFdohUjks
pWZXvpiM+v+ioCI45KLxXO9pbUFsZofto4KWdHUCuKCIic1CmZDNds7AfVsBE3/m
niYKD6a/Te1lDf4TM0+nNj0YOOSbhmfX+36nI/rZUOhyWn1h1I4I01TGpOtzwOB8
S7tz7SmiRrMkdgALVYDwM2I4NKVTEg2V3k6jLT/+Fa4TAnm1zOVFHe9gV1kmlMXy
v6K9LbFlLCZCSd8M63nQsQiBRPHNDqCnKGjzbIT07gU92Eivq1acg2cjp2/u5qa4
2ji64pxFpvGu1PfoMqU9hPxREawQJ2jI/Ym0iUIqpQU85bqikox3Bv529rIMyb+O
/Uz4k+ITvnWYO0H1sqIS254uzf+d/qNN4eDiJV2stvRmEXbpZl1tHvT2HqmM3LNs
RR5DN9rN3/TcKfJ3nGENhaDCS3baHYPkgErSfaZHhCc9g3enxZUEEpXbvMUrjs95
kXkZ4ppYfCLbDSFSmzjht50WktK5WPJWVyBPmuGteIn9n/gvX1WOQTTHThFbUR64
zz78BWJnccjgKx8bkyWraksKE0xZ53xFdzHC9ahaA84zsQGvT2GMwwGSCrfTWZEo
Bgr7ehqAiSpZPmvlc3kA0rqL9UAI5cBCiDLQg5GrS4EUX54et69Evw71r7FEcMxe
FTnTNE0sUmipnUtANl3lvM0nRonXSsueL50Ze/WVdhz/KyhR+HcItplNIJLbtnpz
At+PYt2uzU1Awr8Wk5rLhS9IsfE+eDaQ8jT5rdxoqxPPwUJGg6r4c1P8SuKaWlHy
Vvw69jMbgGQR/QMn2IVQRywEa5w28rTTUamxAYveRKlIJwrVCxbjOmsHkkv3Xmm4
It+X8x4sVXzs/aA1J2YbKo+VVn9nmwiLR82W1gQNMH96MNkGUNmZXVQj+nfRhDSD
pST903z+ufIljkO1I9TUN/g74L5aNcy0nyqb1CeLXztCK2LwJHmfTJ8MzMOBFfGK
pbvHIt7xgDWDwq9YHwpGv8IV6WJ8GfzUH4+dm6rJhiuFdxMsVi78U4wVOXSDl5iQ
LWk0+wx2/Zwuda0Rh7lWvZMVfbpSBpuA+OhZaQGWQmN6zf2ShDJkkSEREP+FypMQ
8QXCXDgqQYjEam/GIRwXwv6/nwFgtStNiMjLfGQmlvD6Wr6LP2Wd/YKPzBzLfabE
Vun2pn7On1coPVVnxcFY991GJEbT46AasvqASQ2u8qbJzWTZp9WrMpKJ/V89gPsm
bggQawQNLuXF+aI2nySqmYDrlkIGI/uA7ZeQsPjFMABYvF0d1UwsbFSd1wgzdw7G
ARph2A291j4e6kPhoYTS1CjojTrSlBb6jsmDM7KnKfpxxamhYh+ja6S8R1rW/FaV
0l8TKtUXaAF5WewjNzpOljoCFnzP9d4xPTCfW9OiZaYREK4h+X12Ex6KiYNkMV4Z
DTFbg6Jq8MiX/agsJNZesN9w4SdUQ1OSB7lqvP33TdxF39aFaP9TQ1hQ30NrAdlO
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eLp8mcao7N/zf0fymq4Wl9GAdq6hWwDVWJd28VpVtgVPd4/FxcmhvQjPHZJ3WWDc
vl8AWdoca+eOEXXMtRgg9skgspOmTmNN0tQe/ptYP9XCBl5q7eY8tL+KSdz7ZsuI
U8BRsSFJEZaamRlG4QB9tMz0jBNJ7deD45m7IECflDdC8tI4LpDn2A+7WfQUP1ae
JKFg/6060iBKoCqVuVUv6aRnfWD+9LudQ+q88JGSSl+7k4gCTetUF2R7qOkaXTpJ
KiePoLq8hZp2E6c3QIS+ptz4CKz0BTOKGMSxbNk65BY8z+lrQasr2n4X/fUzyS7I
2fAC6WJOXr8CjFDyMBMNviheXyk/G6+6M6JmscFij37xgmozhTEDnay9spnfsJbQ
03kp5Y44RAcP2cZ5C7d8lDv9zp9ZEZ4UbEAN2xEGYgnoUzKEaC/n6Cg7q+blx8vC
KnLsbwsxi5uPEzLuq7CGzZIWkqQ/J4C8SoiCEhv8m7oWrStXNzASzLAdyoOqAEN3
7ftLGxJ9GaoI+cAd2UzbOT734YewyuDWeKKdoVqIMLWjosYLCjGuW/J5VCj2Y/MX
u3SajLEyYcx+hQCTiH4hF5DbggDyQ0YGJ62sIn2h3s1/ik6vvcioax6MVuaNLYO4
b4ETNwEADs7XZModPMICrczOwFLHl0SZSKFh0GgHMyFNdPtxoHUWpY44lL5Ienwn
q/xhSHrFVvAp6aYmLZyGAlxQbprmKrd7aXHWyeULqOsIy2bvbMH7zR0xOhHNn7D3
uH/bbZVCVfB1dhWSlTLYRX/+9oZjToxHYzM7jDmJYy+B2jvrxp4gTueJW1aRHZ1e
8FQfxa0Jl+k65acD8KEcMxi7m9pSWwodT7aslKKSBS2yVogFfWOFTggtI/GDnT/x
ZqxFA9FyPixsU/UK0L6B2p1FoZ9R796qf491/PPsshElOFsWD2MD2/JcOIEZftAk
KkXuDh75T2qZTI784Y4zWgwM/YcDkEEpREaoRfXpniSMj6zqgpTE5hsPQqctTvb+
YdxPyE5qG6p3qggmBI2d1NKjnNledh2luab7fVCof8C2pXH9W1e5VSo8LBmELP0s
7bPcYmO96K1ay8RISE+kJClCW1U0/VL2eJWtivtSUznifN1WTIC5nxQr4rV49G6m
piraGASl5z20RIKqZMhC6bwHG8wYj6mk8UExkrYUHa89GrtHlTsZ781vVaWuLtst
ZzrHP79h7PlMSoQsJDdjQ9VzZVKkr4ViAsEdO2KvzyNyT3QE5zYYeWPSj0oCFrGX
CLI9L3t6N9ERi9AS5m1tTB6/UFi3moocc2IBwoNCAxrsDobf7vvxy0LQNMigTtG5
3Aq9pbp6Gnmm5vQEPjkoNU9w/zesbozS05P6j+cK83mQsi83T5xupN0Lxek0Hwmz
8mI8XD+722UavhjKC6Mx+va6g+2RUFtDmO7HiBwLnogA8HBpEW18yw/YiZOEZ+Qj
3wtd1jiAuQvOQkJrp1CntqdSx7zMaaZb/OxoXxrWiJA3SRV0nJRJmUM5F7Mq4h4/
BMM9cPdzlklJsuzSgwKCmGbg9LhzO9mnBNh7Ot/f0yXXRnHY0bIMwOy292Es9pG0
FGGO98Ng+N9bBIWyjUsZQkv5QyYgVuv+5ZSfAhU/EAFZY2VH8Tz+n/NCNXWEW9C8
9USLcPyx/TgqWJJGU4jVOWLmSQETsXcRAv7S2vN1Nbg=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHqs9Q8kRSLm8shA7hiTfh5Sl0dJkfGuFAm4JDygvesbJAIZMbDdXXLKlSV5HnXj
WBtDhX8ZRdb5LA5NHZNCZy7+kmDBQqNoM1QlzieYqSpdK8VC+xzSgkhjZ8p8VU83
MHhT11bcag/nWZF4xcr8rGfkD7pixzb1Y6M5TmA0XqPelFGHLyyrxqKMl4XlzcuD
Pfp2Im40VrYfmklMkGd80rDHM+wlFWxLLh6Vcxy7ABIuq8nijSRM/aTem6yyfpuX
5LSO0lu8iCDPKXe7FKFiP7Gp9gAP3f8bQde3W9dakmLOgflbOfxoYabG2pM4qsqc
zzV0v3LkZiZU+yVm0IHI/NbWrBqPDMqogS2YdULyFzlKmSP986/bucpR2/yMBlwH
jkE4cq69bommHZesEZBHqmPXLWs/Z4ke9SpueMluCzfRt9gpK1ya+g7RsXKqY6VM
aTIlHVfoyuyfqASMrFEHJWCHD38dYu0Magppwa9ST7tzeVsAJAJgI5qP6lXWT4JT
KoKOffXvnztOsT4YxsRP/522NL2N/b9WXa8v5+2psHAbv1VT1mvQ8qijPwW51niD
wk2YUqVAxp4dCQGHl0AW75PhRO91nvod1wp6KB06Omb9LDefYHXqM3X2I1+4xlaT
IOWxUzknAlYp133ZhpcRaSN+UreivjqxRhJPC5XHhE4zuL+boMkcbZ40WcRhX6n7
9g7G7gEbo06caBf2rFzz28oWAiisQ/b1otPwfjTcEVSJzLzozR0QWVO7zI7j5TEs
Ilo55W42MwW0+k/tjl0uc2RU7HmrQTrhJp/9L2Pnal9BczNCjUtxZYkvN8LRrYVa
j6oD9QO1/P3vfzNH3jwvXUVIQ4rbApQVu8nKutAjL5FpvY6JSf0l7yIyWVWjuVkg
0bSUD/vJjbzEsqvhtP7pmPPBg8P4+Ri0fqa80s2ZRRnTVs4sbloMr1oG9OKN/9Y5
ceDFUszcrxaeD4Ee/l7rK3SqW7MMHD3pWso2HIVtn9haUVWDISE9RB8LN4H/YEFW
4bJr2ywL+4+M0HWTig0YBorcniP68ryz37f8gCbtBtgwfYIpfjEjdlw0fbAmHMT4
4W1GP4bPpFCwD6LeQZ9HiPngQq1rTVqNEzY/+qcUIcM17dpd4zVUHvCPCmD3n8Ja
+DzgefgC3C9BJ2r+R+C1poYb4RensT55UhoBSNzdhCP5XCtYFNI/yaKo0ndQb0P6
SCSAkP89RNsj6AOt5xigppE3FCRobp3urtb2aoKL7nVtksuq/ap+n2sxLoMjZMsb
tzdA43Yp23PXClYYI8gIRKEe8if76V0EatTJ0Sx4IxJ89C9j5pIM9HNgQbK9T0Y4
qM1qwhxli8RRt5rT+yWuPRPPlnUqeDxrSOSlnzDmcgfppD7e90iyB+9oxo4Jf28i
KaUpriUEFehBxDeD6huDuYlqurWHVnn82SKW8REpw7BzG3rEg3U9YAhZtE8lw7Cv
4pYRzZZTu6CMHZcQx6+WXV5/isFw5HgyUum4Q6FyMAivUy8wSl7qvm+M+qC6lcXv
3u2b3a0j7O/4/K03Ug7fp9iPb3nVn+2pY8CtOwqDxJAF1P0+dBb4yUdZIydHObbT
/TBeRtdJgNakjapdjLoszb7CdCVPu8/wLmECvz0v+ySIotJf2ioBl9kguwokSc2T
1GsrslwBD94azQrrvw0o+vpFIrzdxmoyPY9H510X/dGCKkuS0Y9jvDqfgph3blA5
HDGvnbIbfxsdOeV0r71TszhmJWQw37hgIyTOKqKX32bUcFGjnttucZDFzyDpge0B
i1XydbGkCDs0slWY3APOO2LNdkEkeJR0EKB2JvH+QmVUOIxFf7kXNF4BCmicvlvb
WmDg7+18WVrhuYM6rlSjT6xKMwZnDKyhfSyGbxvyEz9U+1auM+pucP+w3mfp7B4v
+iCjBcaow47tT6vnG6og0tNq5j7VcijU6pAfHAUfwq+MWZCJv6tlx5sx7mITNH64
o7hkJwg2/OBTFbCWRfQwla9x2mMhiDADx3wGXHdnT+0quxjBgr6CJrG5Hc0/lauE
GN8206cloHo6kBZiv/ie51Fs+/5qVSeIi7a06A7aOhOtyMddD6WFgz3gdd9R7pYM
AELN7XJebqSyQU/TuQaKHKlnZkjTxKU8PORTyhQX2JTA0vnMhTJfTw+i+Xy/G/Fq
AAFyMpdm7PsJVNH90PrCh1r4cY841C078tVLeB9fpxZELOrcmWXktnpnQ2nb15Fe
ibOyy7bJOvbos3qsVnqAtQH4jrAFKm2dMQ5NYqRSuTuguY4jcWz7j2vED5h5TpKI
9FuoU2izdwPG35irWkVTvKoBZf0kQT7fdv5JNtQTo+yBUn36Y8S7ivimuFb3r/Uh
ToAhWafBcnVbV08SI9eaPx/fR4RlH1FbY4x68/vnGFj4WLJn+2LVU6rIESjQXHNJ
MyrQfyRVWDZ1iFKrftn5wBil69poVLzejCkE5Lk5rmvSTGpRC1D/goRiYae0GQy9
JshQGkLb3PjX1UUd2Xqbxf64hnezf8yJ3ZA8kxiQbntHPim8YhyzVvcCp7E297xy
cB988v1yfoB79raQrKXXXUIUUoblRetnuMUc6yjHf1g+m3R2gBdzMxQKWJS4Gw8u
nNPC4+RcVPURhJFCxCQnSSdfgM8YugBaRINlZLtcaNS2twgGNXqDEswpfm0jS1Hq
BFA1tbuOSTGe8w560vQTsLEF2d2l+uDhiheAJJQYGdbJTU/KI+N+7qk2EZNgfQuF
1oxifURTLPIPB8YTRPqUrrKBY2o27v6u4D9+eEj77uvIGX4934ENoPmTvkIOTtCi
FNC5gy5sgCFf24JY27XI9F2KFHjgOWR9Fk6wcEqkZPV+ibTw73SY+pFbCwHpi5mW
T/R2mdfTpp+Zx/B+skG29ZLvSGwrvOMGF9H1B4Rhqw0VNZdcgpZyJAAqSAN9uVCm
g6UjTBovMM4AAL7TR6IavNXex1qwT9Xwfbz1bHzR2AzdXebaqvPZPORCMMF7ea0p
tTvteqVEevbJY26BJzAaUciYQgngf7FbfF5egU5yn9DnqagfJCIP0LRhCTnzMUcr
8B9Ua4YXpwm5S/VmVVZtaaPsXoN2l2tuHkpamoIDxBZdpVwgx5V6TsAnolpH+uvb
5IvMIDlPPwkCSrRVMk72pDcTdFiyOHw55m675AHiRJVKkEt+SElZ15tuWRoSeqw9
W4FkLx2rekkepvjofdch7DddBMY+k0qYsVoa2CS1OG37elCAnq1NbizOJx4AguEC
SqzIpVkGS0HySQ4o4kAK+UErSccseJPvGpBaiYPh26Rirlq7LJlHXHw3+QbZhrMP
KWO6Nl9P83jpropkx5P5yT3pzjjKuGNDBxjfJwjnFDU8LULCNpMIQ/3WflM2wfBf
BAQiBV0MvQ1pE44ogkf+NdWE1Bij7hqbzD4o0EfHTLB8VXCgc/FKkghpK7leHfYW
qhFEJ/xdElXf106ehGHn6o1pyWMBw72RDIrmu1tyjnH3icZk4ueEnEhIGhe28VOi
LguKs12eCWRKrlUfYLTBqM/h6PE4hoLycoAIhFixOz/Gjh+HZWXjlkEhUVn29ddj
932RknsgK9A+iuBa0XBzvSfca/SCG/S9rFzGcO9oFlCY2X28i/Md3MhoRWpYl+s2
okS4RbSby/9pnC1NpaJWk+pju2Y9hPACTDSWh3kiCITwUJS2iixwbUApdq2eT+nD
o29bo6rMs+WHntGLZ/785lv+pRoMCmDNSW4wbi6UTMu5dAko+Ct/Ka7U4V7pRzMe
tzQ/vfHEjFoxmICflWteJS8bJ+/eZjqVbJetq8b9H8jFONlLjflkWfuR/ZcLRvjf
BFA4vYtddb1FIWZgi+tQ6cQbyPhY3FH79tDQQX+XIHjzaJEX03+Xm7JEsBoJPGUr
CiDvi33Gh7Ei5wta4PhLrlDaI370Pls+ljk+4nQ1oFm1/h6LeH/p4gUjbsZjVZkx
3b4wV62ShtP3PBj7aAFT7LsQdpO4+DEbNos6NoNaAZBD3AjYGWry6mVScBpip8Zb
Ce9WIhUk8uL5L30Mca4zkb3e4oh8GiC/iKeCxAvsVCjfsgYPL7YPkvjwxapQrTpu
eh2ZdzJOJhuyzfC8F4AUqTXyxHZxNsEjYLTpShLe3hfXkMoNX3EN4cl8v9oqyL4y
SH9afCds2J/FHo7RQd8X+2zeMp3uadl7vqPNxUKy60b4tonm79SW8y2t6hcPw6LI
zR1VTcWRaIVXV1lDczCiSESX0sqUmsrsScJ9VanVbEuTggaP+FlkcdponoA0aBY+
qHogl1JysW1SFBxtSgtEbcUKYiVGC+1cUUovuiK/e2S2vtbNiF4Z7vekOjQfLmrT
qBujDm7pKzlTHXqE7PCf2yvPpC1GCALkbK0f25gjEoUOvxW3pkXNbmQeY7HXO38R
OJytgSDjPg9RRyc1q+i1nwHIies0jeyOaCNh8T/ft+Am82s7qtb6XY4WRKu1yDPj
M1S906jjUnBSs1s8LMvsQqW51b+SKxY/ngKZ4yiNpytdMp7MO6NkI6G8KE634Yp/
k1WtMBJWTz5KHSTbApkHzW/9Bi5+QVktcoqTZO52tPrzgJAeQRMIKOY/0n4yNr6n
jbdm2/igg4OE1ve15T3OprsZ+JKsrUagZ+DdCFdBsc6AeqR4lpibsr26Z23q+fPb
aQC7EyO/zZbe3FXZwCq5ZbPkOi21IXBQGmQQdTDkxH4Y0fAd26zfPkxZZpE8VRsk
AUEAhsKr0ViVE1Ya6xJ+ziSj5O6Y8FLTVKAac/rvc3WBlbiwxBeAloSVRBnV962O
Ugeba3mtAo58Vr4c3T0ONg51qGTzAsiR6d/1nZx3OTaAa1cPyc7yG3+wpFuTwYij
RfOKIciBMWjDqjXDgv/gDpo07EQIyfYOU4whR3wzrUkvCudYBCrJmSPp4B92FkL7
R97ToU+Ybp/w/dznnFILf6fq/h+AKoP85U08DCSYlgN7cDC+LT6miI7qPQtfl0QW
sQ0YDrukWHht0K3eH4iMrsT/lYaC0lUc8/+/71jUGR4rr+ODHp7kt1Lotpw1cIrp
6coLMalrsEfQjJ/rSqSb0Kc5hupho0hFX/KmfJtf2OUYZDxNRmVJMaAG5ooJtEWc
y9cpQH53mQXzDWu6wklDW7zdz4nlqXtnd0acOClqgXHFBT0WHWpID69IkeXJB6I1
5nkmtlM04++zHHnXNodgG0NfxOB4bO7hzQ3ukA02N6zEgPuFcYFFnOcwx4uC3HTX
Bnig9UoAHSuk8g8jfmA1PJC/CeGO+FwUNuIO+uCZzXctk9WU0gbTL6tdhTg/mU+c
xXlXmcbZVvSrIjXY17vcRDOm4ZPJzn8jiLSrDxQnKQnOEvDnWp8M2cPHJn5n4CBs
3KMKyN2uHlaZBPqJQn9IE3vOKguwdPxFggleVp8MG6UoCD4poT6mBg2xwGv36olX
Tc/M23Z1goCoQdlGyoZ0uM8gLAO25aPWIEUEu1qJneHuHIUagIdfo12AY9z/ZmOV
6sCpdJf97kSVI22QqUZ6kXz3WlI+cxuOynbuBRawExqcmMf15Wy4kX+a7EeX1Nxv
6jzKh3MEkelbtptqhB5vqOFqq5nXvapAJ/zWpL7WsE/HuHmJgVQKqic0/tlUnQWt
gQHhba3HRhXxFYXyOTkSCFwDnCxPykQWctXsjBw50T/vD7khjEiRyMpg0/bcakgv
ufofX2i9k2TbBhsnmpJgMgc2GI5u9/M8UKDCyf63LTNK5Up+Nh7jK/rTgTyoBA1n
oMPbBF+5XvHsdeoALyYDVrLJmlsBdJ8+GXWTvz97/Si+GZBi9yUp5If2w9bhw19s
d5vIaZ1eGj6mNwu8eN/j09eLIH78ZAoJFHGJIrt6SIbvgZeOjEL6qlGmY2l+aVL7
GdH/rzavl++Z658BeBsjcaM+RLO3wmW++cMwKVlXZtczGt2wBlcfFwT9PdyP+cup
zNXat46Bgr9GsSQtvutK97jp0o0gY7+kf9nxt1xYELOEiU8bSG4uFDTP+k6xNozX
tUXsFj/qLZzvlAs4sgM6R4MH3OYyW+jZvuHvH+6Z/Eh0uBUqsl21wKy/hGbpqKeQ
RH0Y24rjoL8zjZ6aYSVWrW4BwFz/H3Kp4z0dJ+Nv5s2f73PFW0nVTwDGa+BOeO7I
mHhEgnT8+wnLfaxfe6488uQqck9HTAENyjFPow/kyMYqRFgmXXYzwqZ+5kRHF3Cl
HdZ6XDyzm0oZ+LxxAfdxVelDs75nqDR1BGSSwFGDRGZkSY2BLZKwhHAeyyv5rBlQ
cFYXu+AobRRkuUDuHrzg++tPhSfIcd47dcDyEBshihXrHgEKXgEKUq35PJJRGbKu
cfjZRVwTUTIRea8rZS5wOG6GqGxfNilna85sjlPeRqkpcw6oQcOaNAPVb0sz18/U
aLI3sb2VW8CJwIaTyGy9XB/KsY4zVfez3gwCGwWpGJOlxoeCZYQuOTgSqgyQH/vo
8pgYy+j/E5kjOUGwTDNCABvIClzYiF6ikJ7E1k5oTtRljUShGEUpOHNA0A5z8ix4
P+Y79mog/HA3uotgNqsbLkmLAbwtGytARp2mNT7LAvNiTQ5IdjMKDmlqMDFAo8UR
cfNVUUCU7W7p49tw7aHs8b0ybQ0V8HsXzF11VFcHXz5VGb162PDy2PfY4D9kjGqL
0CuitHjwKox+mnk+/cUffZosAnudx4LsoLpd9rQ+V8hNb0XVLjvnJ/9p0p5AOQVJ
2uG4YpuVrDfGlN0R97wY+kHanr860dnK/PWnefLWTpKYRl110ezApgG12vmVOdKa
tzjMrDygmEC1bM8CGT9EqSLEY0wJnxMWGz71H4XEWgwihIXgPQCJbfa9OKfhDzTA
wOn54gslnfTU55GGTvslHVfc/4LLfXINzP5YNAXOL44=
`protect END_PROTECTED

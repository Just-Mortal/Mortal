`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eGrvDjhoKEsU8jxWC9ZqSLMv2RNLHZChdt7U0BGN7bUhVT4aylkTY8s6dnTHBHRg
5apIi5BNzUe9qN6VH0RedQKMUzN850HTtte9OVLv26gARK9qQAQGyiM2AyxJcy1D
gEgpOlZVMcpg3LOynVqj7z8EztYYKTswhYhg3m1K6mxwMbjiiumX9kPi4JKzfiYJ
3JKYCf+HDpW2D765Aqr/nNnX17lYPZi3kUxJtPU3zEV8Hg7VY8OGpWw912xmWukG
Vhmwn+F8zFxV85UNI1wkkjN8pW5r34IutWFFx+mus6011unm3wg48PgQYm+PpSKr
b73USNzCA9rE/nTSSMnGML9qZ1Qaz1A7qvHrYrARxOL4JvuSb57wRyKXnXqO7mjP
VYq0XfQYSkMS4UQtrqZ9lVGBZErL7LIFMrwLbbmLgD/CMQCQmQTExk+YgPVn9MGy
0pLwS9uUvA5bjG8zIgypkkepevvU2tBYkwjujQ6Mk4tlRs+z55HjM9gCjov/A6hE
vGPYjQRjfzxRt1AbBstVMKcUUd4YUsqK9z/OZPDq6zYRASYbdctqyNaG2QR1Vk+9
9OOcfUZnG04d3+F4YL8/p+QEBMH2mRm1nzCMDSEmzLpIULEGRt7OMVKx7M1NkKJs
Na3n0ZoODHMyjsjYifwNkBy/spHZj1Q7DkYHxjXc1MgrMQUEIb63y0vtIterGRtC
5LS1XJLKDeKiTkREgQHPU2rwuffvc2YT9yxhDablTcisKpWNnHnQgcqH17aUGQNH
AezENCEMtZX2o0AbZ/dlKisjuY8exVpZ3e7qcyyp3BpdhowpiRla2Kp/dPEjflVJ
tkDEp++vBJAVal99mf7cyoatumYU8qf8v9UG4A7DWTc+Sj3JdH9Gat6nXlXFg2yZ
TJRGcBqpYEf5TLQ9QewneXBcBebXKG4eBe68052n4Pg3Q8jHxeBNJLSUuCImxTCY
IdEK3p/z8npJKFXXGAf51e8/EjvKxu49Ib5AUNVVW6jv1dHf3z7Ym3RKyYDOusqJ
Rt+DYAZw3BG0AMJT6ye5D2dxGQLdawcJHxrPIEqu8sbY7jdYwV83UWGAdq8xu1m6
8Q+oZGUrNeZp2SsVKe5W4pp/IhkEzdXx6WYxJGxRD0WshJDCbNDfn4DE/MRh+y9C
xFLTs+tKOWAy9U9w7vR9/A==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GJnGFrtWgns3kkHKSSmeBueM+/re8SHyH1OT6ymCvRqmCZ7acutr4aLmujKUZWys
mLKpkXKbhiaCOEcc4Iq2INAYoEDPnAJui5P+/9CgwGCXzspChPfkzVurS6mKVxdo
vBb072gs/GHKH6AvY64yj3LHWwgVXpKXbLZ08aau4OBnsEtwaoDuLmBb9M1SrHdk
LBBZPfN8aG6TccXJKveD+g0cjzkDpBHP3XYG/L2meFvvR7DVGZvAmyW9e4mEZ/jZ
t3b5tDYfStAlzCsXTZp4Y8vFusI7UXjawbcxiFU8dZaLF43D1W2qusqkLlgxTaSl
Pp4DxJu70nNk/FUWsADdnxPcz2W6ldIZPARKtWuc+TBGnxs8I8VhsuH0Y5u0EqgO
fC+sgK3qkAX9E5YeI3zVme4OKiffYZDy4mxIc+h/mEYHMy+HveS/LHDS1dTjMjcu
MjaHU1QvqB3ytjyYLC9CR8NAq/Uk1+hZm4pHT01NQw1nw19LmubgbldVWINoGazt
imz2V7l7mJXM+L2yG4dQPyzcJAs7LdV80UElQj25eFA0ZJkaJdSkbEapmHbJe0qE
X8FJJ3vqR+I7OjknntIl6dy7vqNkwGcpjA99gLk5mgmgHoSEqCUYaugpBDjOQ3kE
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7xdVSTjjuro9ARQPRvzkFlTU40qNghMQuiORa546Y4FFMKFYfLqLeDXgyaoT877
wMH/wpzSlIwJImppbyKtWl+tn5OJw8NdUtmCwKZkzn88W6oxvXZjCAYfDzZJn5Ok
wojoXubYbTFVtYis/IFKsqYpYOpLBdNU7DaMAMjC9OXoqDq8UEJ3aIrMZ1FgYUDp
SwJLlV+I8FPzv5Pn+pfDCRaxoaMLl6wbVdk/WVuZ8cYU9NRr2LPX0dcq0lhieORD
vc4Yay6PsiyJpDYu1QRXPMjYFx4iYQShnF37EcrW3qlVF7adrjeci3FLTTpqMLaC
9Fn+1JtlGFTdnHTN8l3LgPmQ9OJmdZPzYlpspa46NW5phJKxCqutWvtWYTrwdHSI
vdRsRPznKqzHXQ2hpqlCdZQdEQJfhHwS3uHLccI/Ic+6x/Mkit4u4pQKTqXHikYf
opOINz9LSR4wuE4w7mAoNcnC+/F8QkH3DJ7IrtPCeW5AqTW16znBrLq3V7HRoHat
Ix8uINO1Zr5GNwC/sxzZOOb447MKZ5scHTAJnakNsGUCcilKvyifR9ai8VlOam98
+/F7yi5e7AmvsJDMZS580O9ovh62G5zmB/fCoEx+v8cZUyA1OCT44h39GhabYkto
utf2IhAjub6/DHw9IjoM7u0PcfXZ06DO6yMLrhJyl5z67n3Yuy6tkSiezAsv5S4s
ANn/xKHqqECReDNNUGfqM98lhcTew04dt9bdvAgco8PT3CKTZAmCmkSKi3H0pvYI
An5pSyOHuaHS81BmYyTiaIlaNjht9XGz0vg02Yt0IZupKR3gxApGUHhbPP2IBoPS
i264x3B7MocUtSvrbuqvnMOaRfw4kc0L90V9mYqwIvz5FeI1gQqc8ZE5E4X6nrm9
JVQpC7TqKqYI4Ia7JXOnF6x983DbZT1ra7FqAsMP1AxPucBE4icg2pfb+8AxZ6XF
MJYLKSJ+daiyjenCizluhBKt6AeDwcb+sXOtO0f1ViVGbYK01d0pJcItWuDz2AKW
LTCJD7raYtLpgMgfzt7v4oE+o44rfeajlBWbYWF9j2UrUsnbfP/AlPgyGsf8wVlx
MiPhuQB1PHJXK5Yqmg71kZeQsotMklYnSiCrxIaogrl+MQqQ3cPgmw24rvSqKrhV
grV+Uf2ym4kvP6wQwnzFqqC3nvq7zYpGPuF/vM8D68ltATI+EKDJNS0x0Kmje/CQ
AOBw8aENqjiyzk5ESgIHXb3pZAEwGbO4Pqmds0HWUUYrQYyXDbl5taDRm6M3f7A+
VuuPmrcQq3vg9BDu3fc8iYD08eQ5LQfwe1Zhqa8UrLConSChw31aVc/udfx9Mfq7
4EsF1nbs8WVosl203hzoHUQZGVM/FuQVqpUtbpI8yogvbKWWoS1qNe28fhDEcPBg
RA5rM9hD3GEPNGyGwI1opNh7KDH30Ili1Tj1er4r0HPpuEUriigDuxFYaLusLjzH
VtvPJ5iMMmvrNwIecaObWjL9Wto44z77pcE/cwSciM4DfIdOI6VyKOWMMAufONQx
uaf2nMqmhdJQ41/sptPC/qPQ03b7GKT9SJKq3INBFNmQsiByQc3OV1zUtcOo4PKl
cUw+SlrLoC4V++aS1yLd8MbUvPl8JTVGtSrOclJVygz4menJgt6JVsKY4oQ7ao/c
B6/e4BcCkzkg8R6S0cRh4zNGWbo556Aipzcp0eS9fUEfJhiaFBUlZO1sqR8ZN2qj
9/RFxzMgcG4/J0PqCfMOIs33A28csSMNdda84EsyMMOKV7jjAuHrff3lh+Ln+yL5
485omRO3lA7qASc2VHzgYcNureSkZeHCQR8UDjNNA6p36Sq+jF6WaZil0d26FJYP
+++fRuHuYcfnGUslAtoOy/Ya9jHSdClBVHdCdEhOymBvOLYH3k3K0veTyf/ANukn
Qu0hB+3F/74c9VYFb9Vat8YrVH2ldsjHsDRqNulcXMxInk//wZRXfSz4snsb6UPf
MmhyIBJos2kBRY94tM7skR2+zgEeeGL1t2ilqU327WlBHaD2eGLqr35WDqtluYbx
kvo8GgR2ZgRym0S+ETizsO2u9t5mn0GJP1fywjS9regaiCWxIk6c0dJGBHMwTV0N
URFZrbk11bACxfXsAG8/mpw7nOcLtWbMWvA99GVTrxJxyIqyl93F2+TBNFKDM48t
EKVNbYLrGd1CMJf0y+gZeqMfVTOscrOTMIltPGNbsXV7kWanD3JMyAza4jjctpIr
Vm3tPEqUSEc64cQd7rRN/ncYpJXVfPk7m4LORB6we4uH7yNA6oFO6VljapIiK1zo
rh0SpzKHbZ2MyXKZtQgzIawJDKw3CCxC74nHPlg2svVzECOMFiLD7rqZsowtDwSS
Ucww2JmNaEeHegHt090GVUAzbn0yArGtKHlOZESL5mgR/XSL3ZDxzprtDG+IVM9g
7H2B8+9ynD7HVOwPuyek2dEvFZ3VQy4FbAf+Ka8EzdwKuzCRw73fdsf8CSCyrdOI
bLJx5HCm0GpRU8E1nqPYWcZJ+23lDCoaHMRJHO/BWtbGPAShv+T9w2En/9Sre7TT
Hz/Hj1bFIsAE41opf+GAZfl5ZW90v1UgIoJP+6Gc7AMYXl+Tb4cMOfQ2i0A3PBCi
ZnD3UbpxkmGPPWgi8ZX0D28vV+SaljAGLRJwdo1LknX0RjPBpLNkCXoIaVtGZfpy
J6O0ysBjCNnl3GODkuLdbIDp0psvXevWrFBgfh8+x2lYymFS70L89pNKiGJclJP2
B/rdunt0hHfkxPCaSk4AxSZmOMwYptlXQGJT+Dwsiwd3NlwDQjV6f4UMoPQrO5U5
8hYDDyfjk8rxvVVHuQY7+slNQC3EN0YVal24PiBFIEemyOIiJrg+Le2jZv4IAnEz
IpRYeyWtV64XbuKpsCff92nKo4CswWzoUApJbLVslZQEojvO4umrbeso8WeY9dQV
VpZakZX6wcTFbGPtxuyaB6s8Hd+w4T4p/+f5tdhfz2xeK+9f3v6dkbNLQqsNYekj
t8aSRWGQPb8v6H83mrD8QKSMzIOZmfXlSKB1EJo3/QljTjjtN1KxS6skHMv9gG12
KaMUTEpnB/OWDPV6CwU4DaNKmzVzreUaXx/+s7iQppXysG4KtrdkWlhopxQ68dpZ
iOrffae5qv1GIV5HcHaMwIVw+9JzroyvXwuaNzeQG06RlL8/EsxgzU3d/yjd+Qh3
X2M7iu7CGsnu8qJBhbDid6DakFzVn/c3lanafWB85EpbIb1x08E4A7KCBQ5bFlVj
FFpGz/OmD9M7BHDLtzmkOlo1tTN/GHeWHgGGhN+GVpSovkdO0XwfJSqAAk0kCFn1
/lUOt2VWa+u3VvbFm4plppM+ScbnsqldV91XsaTWq1HYAyH63ApKrTTjhWTv7J9J
0J2OvfYgTOv08J6g9ypLmHRHEW+KpzLelZJw6AF1g9kXRDXoOwHK2yDQa0vZHi3h
1MFCEpAUF5g5ymvc4+KyY1P8xGvBFr64rmaFZwThmhGB36cZMy94NNaubov75zOe
Sfhz/NTSzGLRWnpX2N8w7wV3YKw32hzQsGKHd5xNMcad4q5UzljIIJvwu7b2qgfT
KJWmGAmHFJaLczJc9+vEBOC8nv2mmdiPIGu2fndTK1PHFoTOJr4X0tsM3JRF3Y26
7g/KqwKgOMO6f41nUnDp83znksIVtZcezvjx3QCT/ILYfVBwAUrIg/CKNxxOWedc
b1J3RPSPpn+MMaPvtjRLbFWgehRPR/VzG8QESQKr+7DS10oZih3qTuSWaH7d2Yfe
OgaaMRO39VA+fjBQAkbIsQ9zxRLssYaJBKYOvb8P6xdZ+zhSkMox6iU6nP85i9dC
/Woot13P3y6p9F7nFGPEQnR39aZicXPvCjZyETdb9lCZq4cNAT2We1q+g410Pian
MVuz+kvJQ3nkbQ3PIKpg0bNIjFw7h6sIQsSA0sSERBKMbzygZXH5tmtcfdwGSNS2
wQcmLjZsLhRERRea6sjkRDLFOSLewpV3bWnOqPKKNffDtuBu65iXKnMVuprhAGE7
Q2iFGZ4xYi+YY38eE1hNPbJOvPFrRPewF1bjxorzubEo9Gx0NsaQOmzWnG05Y+VB
B1MCuJXETia3ZLQD5IyOXqrUXGAGnk96KmhP4sA7QuvWqGpJUHpNd5ozdBkgkJAc
FtECwXJO3chxf7YkOzSzR/JbuwG0uVpgxj00bhda6YwaZAM+aY5bxXvDeT9jnC9r
xJ+0+GV1qi9Pthq2DdUxa4gyPWovsuWhstgG5jwe7Wtm457CIEcaCdpeeLG0mC/v
ddY9B+vxX/cl9v75hSkZrcAkiTr/hDJBILlB1ei7pACpz1H00QYX+CmFQL77nqXP
fPj82N0GPnX4oUT1ETLM7tvNtV2ltMrCVmj/PFhk0QtnzpBRKXNMlKlgrJF141EO
x70F4Fbt/dRQTa652wWau8wVIHwe2E2ZBoa9/MgD7F6su1JoJCecd+PASt2t+yhT
c2gvbNIqTT2LZOY09iORMN2hx4ZqqwkM3CJ8MFYQSJoKVl3SRKbf7R/QXHrTxwAl
waOBf8nicIpWl8fmGkNUq+K3C/d9ggXInbNkY9YxKE4dkbKV3dAcWHQF0Jh0IoaQ
waCP5i+k0jECv2Fa4LWCWypyvKPVkG4lVOi0pg6aPvIh+2tdOnNDVOkRO7kPnAe1
vKZoidApyTGcS5+XpqyDJNmiMznJK9GaFzikwEcOjv8zyBWc7eI8LwR0zhKWC2OT
T1fRu7+hBy/lcO/hflZ/5OAB30k63a9J40prWgWTBzvv70SA8yanrEVUY0BwJJXp
i/HGi3OeRki3wFtHIHUndinqVZAx+/G5yP42OP6t0z99e6nNLCmu9p6wZ/QeKm1i
+VMalDdqmSKPm/oxPFtuSN03ooo8GWYh79V0/aMrEVRGgFLK5kMWiab2u7uCqNGV
cA3HYahiB7TKwLaGK2kAabbNx6whRiTKJdkgJDNG4LOU/zx4ycoCMYxSpgy4brR0
4OsJfzpbClarAng/rONDTeED8muVmj1/vlLjMIWsXL1+D2R4NqMKjQ0t8TTlWASt
k22SkzNuoiOQlPBfJoituxffLwBVaJC8cCUnK7/zbSsQNM1kb/pJYCPEe06GaiJp
rVYl+q+stak7ARe9VbnFcHXxFDJGkezuZR+/Ojy8v8z6g1z2gDl+b4Nu7Hae741R
argfcp216zogcllMY0pncyDDttSUs3NRSuve9PZI6zMcxkiyjQdpPf52UkRGS6FK
lcibu7WKlcY/UyunhprEg6Ks/NRDIAFJSpWDpA4DQew0WiyFbp4tfLZeGMMLeOFw
HheLkZoVTyAccGRk3HDQgVhuKUvJCAdmHJeOSq/Y+7jYcC/6ZMs4r483VEUwbNP/
bTde2+Ee7WsYA1jWI6iHaeTWxVyi1wsQSbQNJOqUvyA6iqCla56sLomOVMv+47Sd
HbIF6AJkNOWHcenYrSBZx5vkQ4fwqAUXOuv+1Z6jHBiAuEDvCWIXOhaBTZr7dKI0
dRDQZ+tQnurruiz+nICLtg8zha+chTUv1h6ZnF6WGwb+wyKRBaeP0xz8tOtVHYm2
uP/dHKnGLDE4QNydv7k3fyOUTS13LcPiwSsMdH/lh2LJyvlQxki/Q4elVDsrQ94m
F/VMJn5kOrb20pqFzYEVGc1e4QF6CX/ILa8JpQtOcd+0FCjvJd/5JKMafxq/KJ7Y
27OXzAyEyUERicnNbyzunSglGNKbCnOM/x7M0IQUzhlKk6xNoreFF3pQxxAgofc+
JN1dKvNvTM2uhlK685Ng8TgCF9GwMpk0ZfWkUh1l8b43iLZXR3lL1D7kjt0uWIqa
a8Ey4b/UD4fHCDpXnNifop33r1h8qsS4uKnCUuUQJEg00YlRFJJAGPzwNKAjDps3
+EY843pq3k7XIfvBq4M1Q/qvhWeNirX9nufiyvPlAMho0NwQyBjT9Qow9Mz+avJE
y/TQtwGye+AaCj2U0ufF0lWugk9vIrOx9j1YGdSD+BGFekUpGKiatoOQnsaKZzDE
TtCQL+ceJHqC9nCaDer5SNW5hLS6At5upE7Eb8gCrBdheM96vskSFCO0nBjbvnhe
sttdVlLfW8DAuoI+Orhd3olhaqbAfbSID0FY2bTUWpm5eiT/nfn7CidIfbGT5d/4
neKemI+3Jy9zLdBEAZrsBTaHs1hjrunuqXmNQh2CXGof/iJiPZR5KixqZY1Vp2dA
el/sxqaXIgJhBv3h2VRJqcMFtgj9/Yj+LVj5IZMo9Os3EFR/eDdiJl06756E4Vz5
pEpwIS9UJWSpfMiYmOqTIL8zNq6M6eXqZFqsOPgm90mgMvjcVBxf6XO6jlhMHBuE
+wHa3EluDSAGjwsly93HVSwStUlJgdCOlCa8kUmjUCWOSpbYxSDB+ppSJFLg4Es6
C8qx6Ru31Ej0ilBDZOfG5ZPtkB7DZzbHWmDSOdyhNDIlNbpI8bdRjB0E54NN146f
wwpj+lhOYIIKFW/Nlf5OB1hColJbKAte9JhPE7jBv76dnyvQPiuq5Ui6Lh/xXyqv
q7zmod9CEzAsJRhkd9UBQqAUparsnG1wYef1e8JIQPPbAqqtRm5OD/dZRPR49/nN
207akQLS4uW+Zvgm+e+TpZCXpOhufvI40h66UnLPhBYSsz/+2RvS+YcdvhiW9CtY
3fn5n7XhGMh6XSg0PFsclbcj6vYtyo4JCiqZvKCzOgSxVz0qYg1rOlnqjcfmtUh8
noe3XZroepkKwmZmagam6lOzCixwNnO9Js73J8NkkathqTg19ZkhWYU7BrpNUDVu
/FGFcjD7sn9TIhMAMClxZfgWxk0TgBT3p1pHLCjh00kUPBP9QdZ/skTPYryUab3y
/ekBlSio7k971TV0VrSOh/XSX1xGD4rk8y5qQ151dPUGDmcvvtqzml36YpmNNHE5
GdX4tYPEEQ+1sY+8XqMS1c2Zo16VNqVaeedW0EKfLORl11W3N8yO8FaL9YKLik5u
V9FyTTxKERlDw8r6abbi2L6+hFxxe6OP+C6q8FWaNhbNSPpBgR9u2TcE/8l2j2+O
VEKqrUokoCpIUdRNeFDpHYLY2WFI7H9sVrFiPWTLmZ/K2xYSqzxP9Vg+miiQpJZH
N7rUExGqxQ/D6DHedUiol9ubsEP6GxrQTKwWy6G6hx+ne9SIVVicDaLZB0XDmvlZ
sgSczPtn/XgfZZYwpe5oAyQsQs1IROHBhvF+0bhTJzl2QkicSoZRx2TbDiP1pkGv
YY+vjIQ0AvBlmiT0iLpvH5KHCKTFiOMEnZLG5vZ/6DwMuvby2TLlwkETcjlWYCC4
Va0N5EzddyinOjrXl6SaB8ccsiP/htkcFT2ujJjCVQ2FGQWhYr0hE1OVZLSOL9dq
VAJVPPueA4C1r/De423klPomh0Dww1ZnPB1o2ZQkbWanjo9bZcDzSxPNXKIV/QId
FPxh5/nOneyEpkJ/F4LUePX1ibA0GUWevm03dMGXlDUAsH2GhC2hjVxGmBbV9DHh
AtW3PSxq8NUWOzhFB5SqJs0mPFooj1yZN+o4qbCHEJGo9u72WD7ea1CmtHORmdPU
aHZcq0myw6NgSKlg8Ntvoj22J3u4BYmnzq4wQdyQ8LwlABS9c6MPdiBDcZCXOOpk
oj6XWKtgVTqgOQWXG4bcwx1xeWy62jujl0+oCu3rHuNF6cD3ike4ubqir6yJWurm
4bVcS3CJo10L5J8iuJkCyc3m3mFiSxynIyK2RiwMvXAJ3OkfaayXJrjvBzzucg8t
v8BFCwoTLk/dUWrNdZTeo9ifaFVwlM4sAOZuHHvYYaivzcHiXusukOuuG4Ijw6jR
CR875jVtstBQVa73t4J2Q3ev6k5IwHzq5T55TC7jY24LxFokNvmJegcaDojgJ0QJ
rIvkmEVe7W1bIiuTbwSCOBT7NYl13je/Zsba0W3cBzwbmMCB7Ctcb+RsQgN2aEQo
vyN5MAz4e6uvnQ1/ysKWzqYbPi1Nd7ML9kNJbPKKgyWaixmtzS7bXf6mBHKwZRq4
FX/flaClBMUfgSQ1OUuSTz3QZC2imA9oBjXUqHs0NvVJ09SnzDXL5SG3lt3N/GiA
RDyVOWPGUYKxTXmJfS68JeAa9YsGrHjvSo/p5rrS/hZg0GbSOC+1LALZgvDpqbZ5
Mfmsqxu51H7QJHmP5A+NYJlVn3D3GuquZ/ejkUKUOwm268V+8H4ds57S5eLp3Nr5
P6FImd9K+X4Qj01OXLnLCFGRH78fi/pI5Y6eWA9mLU3GCC9yjjqpZ/yUTE4OV6HV
4AskWkS/ZsHbjE8dzYAYuqjig56/Sb/ScfNsb90B5F0bCcOB3VXJFGUISWhSdHzi
12D06fCLulY25STTNGc1Ia8h7NLF81x54pBuLltDG85yhDQFsqAGjF4NqdZNB07a
gKcC8r2os8jGtgjssrwr2GHQtRN07fsReF0NIZRtwqAdp9RW6LoK/oeCI+k62EEx
26U8DF3UIsSJjAvopKFXgvRFA/ph17ct6FVblQu4CDkYyTyB/YcCmyZC6TOOeZ2o
f7ZMNBZhSWmCg8KFY+eHmxopMUHbziDRJtzGF/1EyWXQqiltIae62be+l0sMo7mF
b5AG7EaZD9fWQzoZ6WkUrNHA4e3DnSj/WErcUE0QwizNj7eyXKo8T4q26r0C8Kx+
Oo5N/OD6F5Xjhse44FZkQr8+5mHXiPT/fWlLinJObqV6A6pMtNVkdCSgnVxjt8+e
lzz/nyjUz0DPF9jBpU5erNt4B1p6SfjrdE++zNJcc3312SBniHByzPp9KQBSKTU7
r8pqhIU4CcupZZt0PHQXl5TpZ14OeBD+RLdPlzHGCDpeYAVp6z6CTf/YvXFGsN04
Zx6YAonefKiYWe/JGhXHAP5gl6JroY+rsT5Mx9LqELH3BXm3QSVzd2ZL1hhMOVxn
ImAe2B+YswBm1C3coLDdmiia4HdxyhCQTRmhSlflbj0eUuoxFwjZccpIOu9oCYzn
qBzBgJKYArClunnM1ouse9X4fgnVqdvKfv/je4NKOLxTj6N8az7bm5STo8b8DNr/
DIPrHHfeIMenS6xPiDWbD7gKzQ++alIy1FYBOtZ1adZgOLDxL3c6Q3XXeAkbCTm8
QLTLfW1wqiHwjFwn8+0WDhjGKvYazM2Zdym5uOwshVAngGz8nGjAIEmpkW7wua3c
dWqUbNZDCMOstkBxHuS2pnT5wLfkCFq1fqPvUP459idwEfXkrgOboVTWY8DntScu
fnrjDBTnYFBNvXJFSTPbBiNJSPmpqba5BIFHglQ+K8zq+TJ3yWFM/cf52esaKtfh
KikQBWeWlhWm9e7YFxwYxXu9w2fkqLXnmJm7N8M7w+eUencRgSWH/PHJEfWbWbpu
PvTAYWLkhh/80EtawklmtsFdfclYVCj4wWPgTuGw9TVPuxmTsriGdEMj/Cb9HleK
i+v3VMzjbGozV6TkcXdj0q0y6EfE4c+rcRdEjAh7Fq8Vx1LdthrymARDUCRVxbbI
3C2ClQQ0/pmp7dUN3CmWwgoy5nQfUBz1urkvgQOmOsZ3dnFlB54+ZyxOacGCJeks
7DIzq9iagcyoY0vAaxJ1Q8COB0BzLgWKu7VB/QDneWb6L6X0LYWaTEKDyRCI5rNH
nghNUGPCTHORdb9zYwIzTRDln0A5c6AgWCLHggs4pq7KFf6WnDaOMYjc6ypeZO1s
L6ibd6nt211kQQgPCeUjb2/11Rom9JxOgor9qLYoxa2veThJLn+5G7GQ9klF86I2
8oRxMj1doCmHaGtprHixuOmh+D0eaZnx8Ny+xHPrJDQ/7/7tpPogWoxjw//1u+FD
e4vFIUbYfayzPecg1UL7U0D7zJ/KGjYvWjmiqNqSqf2YQfPIUSqSPnEXadHoJpG3
pt1vDHmrQPhWzqeJFLagY6uW62WE1ZoFa14mtFvYEc1igCEt+UWP4/d5mS1Jw/5c
jvEQ4uN1YquUxiujYSuKnZ0/ZFJoJK5wCGhjAcHF9SyAsTsif3TMmIp6Gid6WZPe
tBZSJS72U3NytiQ+hO7BVfk3vH5F5SOUT7oUNX8unP/5XohfahfF1mZrZ4wCSHTA
QXhHYmL+jIa7PxiuKnEXwkRv4vmhHeyJxQdM0kJbv9u9eryID4j28SXK482b4n4B
F75P+9Q0eEu0P/DYt3jRYk64a+Y3r/IB1m+zupy+qu4K3lxjPtyMYISwm775sUBc
h5HGZpNUy+hhFbG2YF1VaO6Dqu5CgQqQU9zeIalIpHWGdFRw1aPN8/EJDMjZ7I2x
mr28YLNiFs023lEzqxh3HO/Y+Sg5YDF7X+dzZSU2e4SHfDYgS8u6/5ICIHic7AbG
iuCpwl20Iu2kw4SQ7s19CNZwYzq9ZsfU9wm+pVQ6yHe8trALzwOVbXZWqrgEJnVj
A7hPVAY6wsQPi2xu+3zTwciPEkSYoKjFoBU99pvOfain2P6t2PrsQse0m7Ww/xUD
RAy+jdK/0dPSK33uAazqnyzu5PaqpCTFjZjEfng918FYRbUCtg3Vzlc2UpD5BfRR
enwQ12xig8osyP60rPi62Seg6SBWCvZbr9QEGV/6N5gUCCxNQWI2FKPKKfkuYGpm
eM8J2IEXGuPS0v59LXnsajj0bg9+Nfy15TS4WuM/BTzVdQCIuBCLzDKxI29R4cSs
Vll6aUtVZfYo9xWscJn8wywk5G7ZbproLEVVXaCMfG3rHlFY0dVS0ibu7iRupdcZ
Gn/N33tX+3bo9w82b8XQGmwSlSHpqVjk8RNqCemOjE/0w+enEkvWfJOBlDN+6DGg
TcmHlvkf1wmsKDd7uhuXGSVkoU7hug8wHUU0kU11JtgbxRNACPXItfBrZXSC2jZG
lwzKApaezULiLfiB34sQRTMc5ju34jXuZUA6sHWooT7hhmiIkFBnBj307Wxvayho
sPUSzHfb+seSyRkzhydVtFzJXUHobYYAKwaTY01uiUQQgssPlbrPAxZFG4mLHOws
LHZfqoUy12x2t9fjMSt+hLgO6+144cKPiN95kiEUA/WUUdUOmLueEmRHP4h8Lsoi
faU3bIon3ZHWR6Mjxc8K7UuP78E7ZHXvtFpbRUgnHA/TWXPJEWJQayGld6cssjOt
FZ0ZSgc6Df0f9PGSlrST9BkSGcEUFqpnbzZ9S/eI0AQTfyc8ZjeBkNX91rqSzqBl
C4WgKXTSN3ZWp5Y7H9zctTaR3KNEqNbHDmuuJcrelSCQEJdO4++dm3npEnL/H1AO
KGz0Km7R3ZUJri2Fk2q8Rt/yj3OFas4ZDe39G5XGCXF2VBpr5MnE30+P7iSKaq/h
rATvYRAq73Jn7jqW0gW4Dgj1GGMAaSokAUu4bBV/4f0xIM7Wqaj8UCaMSw0pnO3h
SoUodhXAaQ6E5rBSzXfiG8EHlwrXrxsEGSyaDovPBwcZQd/Icsv5Ptg4zSMoidIP
nKBZrwhRVnxtUX+zLtkl6uF7OZSNKtQj145A846j/VJXkNGo165yOk4+Xk7tCmOA
6cRek4gI9L4sDNUoxss9kSrAGbiwfw3lJ3Fi8v2TxnDln0mvbULk1yvlWwMdp8DT
xGuPbnW7tLffX2yT15nmEiZmwb4umn92ECAKqyIcItUdHSaMwIwuK2e0weX9/OEk
/3psKdh6JWWPOtd/09Aatk1P8a6tu++m897MgxQacx68zxNtdwG+W0QUYtMq96wW
phChtefdYgbsGGGspug4TvoswXwpa2AneNC+H2WXFnTlHwsTCdqUWLj3YEU1WL00
vTeNjSBWakU08BYVdl6A6NUfIfVFHY57wrVdt8SqmK2uhZ4fOfykaJsnZb0F7HfF
USM5wT7DYIEWvoNq514pc7NjsrQSB59e1V9vB85ADR7a2eOnHm4dHVVkArC9Tgh9
Hcq/0v3HHNYlTgtztYlcxk8P0nh1vQD9PCuo+MMjC4K/csEORKTyTau9UF08lVo6
IAhIeoCOPwR3FcNzXgpj1QSWVyKr/LEUpoWf/anh7Jlct+SZf+/Jo58e92eyRIUP
xVwj2sw5q+1yOVCohffORQkZZF7+S6IHFpI4cDAjk5UKVaESzCS51T4ev1RiGHq2
hwKFuNFerXuKk1Sq5N/eVO8SCSOGi1fljXwcLpjlAOClury3XuOLj4tdJ/sNUA3P
el6e+sccprKfabw/xyqPx8i8vxaopBZ9r1POzQ3sDeKekEoQuvN8FhtGpgHi0XCK
0n3dkMFewBsHZPKI9OQp7wLTc8zQ02olH/8mv08TYldg7tPFl8J5YKfr97gEDKJw
Zyv/T9c7K2oqKXd/B03r9Ms5ZGPVnttnJnu0HwGZdS6+mj8BGf0rPXwFfTy/He3C
kShMi0555e5/upbOUYF1QexdiEwghqXhcKVe6wl+Gy1xMDixa7fLaA2MEX/jGj8Z
JifUAlBj/KzgfZaMBHg31m7TVuTYrdPJTXC8GA8L/nOCjByhUUIPxgfzGGmHHAPI
RHUIHPQtRo584zmvuWZTdd1MwAC7e0kOFxic9OCYpO6SWwN2a4eKybVGJEAWpP+1
kdHggu0Y1TvEVJMNE0eK1G2TCw43Mvc2JYR7qySWqiBybR4UdkSoNDNBdQk4pC1v
m1JMo6sJcEtMCI4g0aHnvS5fd/Cq/jwF5II1CvoXbAbqUSr2pVaFm/yv22auLSQj
T4h8OGD0C3/y6cSj6D1rBDCJdIxpPJHq2fe7kThCxArre4UcHd5Y85bQ5GF/WvEZ
+NxwNlBWt5iHSWoLgS7IB7p2iJFJdRSovYZrheTCH0f5zb7mn/kEZpBPvdfsaZ67
pOr87rXE4LAQ4tbXJvVWIMl+6GwbeaFpyfVoas1fTf6f2gT7F2zmHcM+ACWnzdSA
pcOIfkOTjhh2E4iZO1p6XFW7KFBqAelSWClo/EV1J180pHmiKP6/u0vPUgAi4BR/
F/RlK3aYsJxTQcit7QaPWUdpRj8ZoOc2pE6KGn9XQ4uP3QHBJRwueKhr3wMRfEF2
uIhrDQOajYSwfT04yENBaMdwkv0GT0lCf3mUnsPo63omNXBkD5sdCsJCfebmUvwn
MBJ7SnqQyWJfnXfXwbOiI/Tvn/EGYImgthGGBxLYox6Cqmv8aLeM+CUxjeDkloTD
Zl3zLra2IzZGO6FnWqfX7nf/6h4jHKEDnPSve3LuE2to1m0Rpm2dbDLffOazdUjs
DOCQu+D/ClRbiMXyUJ5UDWLYA2huv2piykmxqUHlgB4oA4pfVHrCoeSgi5uEUfwJ
EKEE4HYusTc+Kd5t8gU3Od26NegUGjZJ0rVYq1sUMUkdFOAisacbpYfklFvo3dvH
QrzS2w1u671r+DYxT43bkZXk010No9TnKkJX3jQLRPWrYX70Z6vmSXapyGag1ePM
BF6W0gyXejmB/FjyxOSH6GXntwyKRKRz/eYhYxADRnMiJzQBdyaJ5KBiNubtLnSk
cb/wa/DNyg6sRK+0F/ZUWfP92NxRiKYqtGra2vM1QIeR+8YtFJfNcCIKcjJBmF6b
ETXee3gvGgd/jR4jnVc1GsiR52HtK4UvRrD38HqloeJGk2xBKVa3q27nbwJ3FbFb
STdAAU70AoXxiCNYQ/E3PmOINsleD6+PeCmVMnH3iWS0EDwSCsCB5Qu7lsItHZYm
zXtStzMbOIZOIe7HLciha/6Vji8GuDRSIQzlNEhEpTlSxoXNwfXd/Uprybz3AdGn
+wSGfBbOqE7QKgwivU6SCuGUQbDzmwPKyCNs1I0P7RQ9/++WEPdNT0ugw7v0HQJk
2gRWXBoQFNKc63poBDF59CrPMEZ0ikhAnyvRo12YyJiFl3qXIxeVZ3ySDHN1GAL/
J6xSWFXUb8R6Et1e91DbGH4itLSJJm8MUrwFScq0lZk444kOePSPl7ECKmnF2JD9
WSDBGphHt3YAei7F3baCNHmh1UesOvPICwqyn/zQCsU1Oidoks7/+C7RQCxG4WXh
g4mOKMZHwK4KMWPMHX2jExldIX1nv2AWqC+aMKf9dKcUe3nzRLcLXJY+d03xh+LP
wP1CAavYaak2oO4EAzjkun4QcmEttAG5vbsjDB9ToHwmT9V5PnE+PbkZj+Gls28e
aqSMnfvGDNG7VPl/68iRuRqM2kQ1ieZEaN3sJPyfj1WM+VnroHAWC/3CgpGoCZYL
/s8dFXfR9+SM3QfYjkhj0h4mbTUlHo/RITZ3V1KDWzlBnJrQR40uGj7vMZ0u3u0f
bttmVAtHUh7ymHqHyBjD/I8IUL9oTqTQONuG0I+FKyty86kGiIgaZhX3yPl9QrlH
d20wfjNXluvpGmD16KFY5dHzxlmAbh9Agn05h/lupy3hgsXuugYs2Aldw1W5YSi+
16+WdpHqzGNbfirwvp6DgEG52i4MHO1IGDGWe8FtKOtUyJyro5lRQ0VbilHLEZeA
eBFmsHP69LJOM79JEbsRHsTdoMGlFwynoM9GOYVKhWG+OBRycJjQLkvH4kns3TqE
AtTkEDcKadjF+GFVZeq3lcVNK3f7Z/JEckgy1EhXEhQwuElwLPjpTXTqk2Cs9Ba3
UnnxU1KaMM+pJSGJ0Ol/7oz+DDu5K+kwT/P0lWgLiVevFhvkz/cYr8PP91xHCGUN
VuljRzZvki82HMcptW1G7rt7OCSAYmkPtHNfTRvPZ5YRBGrQ1Qm+0zT6TDKWR94A
Tj7IlObzZp7GtQ3kcrZKcmRAV2Kq0Xk5VL/Esb3xcQAkqUwMp65hEfzPbRKyPHuH
48zbpKrAKFZ34nMxajqqRNO9VlL0LWAkFeyRZL8oSi/gGilvl31KpSgzLVf0R5FC
H/uACEpBCi7U48l6A+jxIV7TslIbecu8d2hDVPMaEQy+FBz36gipmDbfMmT1QDKJ
FPKqnGLGYdbBipb84eNjCoC3ElQcaGhXT9GMrU9Ry8HIjTqjREgtrofPpyqb4Ekd
II78Wt/TN/DOy8o3T0jIxuy+5/9VtWN5jfmictYo8+8qOfCMDGXWrvYEPw2Bzfqe
EtGwn+ufRhgkrsW/kQUNPfXvAF2XDoq4rINeUPfYP/fQKJYGGUNfq7o1rCjl3RMn
JbIcWeiRsTjrkuNk9oCFJBBp2PHaulzCpScO/K8QVZ3+G0A794vxzhyQS01l9KpY
83CPPyIZuMUrqJ+FlxIbmLaPPRuwpk9YM9wlAOUlfe5wL+rvuEjrFnqs+nSNfHfe
OICyYrg7qb0r1C8ux1GtRUcI+KTBDpwWG1ArhzZ+1yjbS2lCNxI0/hcZjJzG3dJ4
xW50o0TDzxnEgtkqRDJ3osveUX9MoIr14LR+v4gC8Wv5stbnUrc5yZSotz9R3qth
/sAMReKE5x7FGByVx6niL3exa3MG0dH1hOv+Dft5KcjeXQPdbf4+YXlhhaur573Z
HCxKWGQMaQM29j/mjhJXdLWY4bCVnFCKpt42cagsgZPzCRmWcAMszJdy9kwYaRhl
Jj4wqSqDCupg+ALHJkUVDzQ2E6PKO0heMO3NpOksJZETesWnSQs0vnjbSVXy65J7
IGeZlwky5yX9PDkU2kH/2l0Tdc/TKddXQuuSinqZHtWNwRhETmkKN9mMRd5BaVUo
pCA7Weywlk35ml/cKcKMatEgKlpv7K/Y3aPzvIPgIyKJX297gG+vphmOmBUtPasW
NVdmZPl3E2wDFgSv1tFnTjxOupEg3ZHH+OKDQLEghlrJs314HR+dNb6C9GC3by4V
9jZ8pk/lDy+9WIxmEMRjAmaPzq7MTwrSLD9OUQwT6san2KGN25kS7lBxWhbwEwZe
Tn26HF1wa1gyoJo7gkBinugm2hZZTlHeKMg3vj+uWOL2NE3KWQGZ40BwAIvmnZX+
IGmb0uYIcPhRIgewQHyizjx7EDcPvQy+qiNbCwwhoq4H5UPYQhJSAXJA/e5XeQiK
3ZmTztnodXH6t+hNv6EtS/tkSyiTapGhbKo+KFUgNRy+0xq3i0Sohzn12ZchVtox
DJEZrIEuSvXCiWAh6woof+LjUObfgSLWI/WEmpVFF37T+VfBWcRqpFv7a6aWVDnR
Eclm5ukYQInAj3KozFXzsPlYTxh3tuzraU9drgqdowphfZ8KRQjFAwYLUIDCNR+7
FdH0rC8OGPTaA5+bVYVjtIM45aeCRg3qeOx7oGDMDxJqXHdSn4TbYaftr0IBG3jg
80rBhgVBNz6VoHhDrznbnFMOtPEw6d8gTpH++UHdF+ebmdUtizrOQmUp3XTmnVuL
K4qnl2OyIbRD4JZcB3w3KJDFqgacjA453hBi4xdN5aEM5BHS+Wt127KURCZKd05Y
Y3mIP7qtRDwVXokrT1tn0SlC2P6BkSvTDvENfSYYC30XLAvBgNVj3Pz2D1vE1HKY
gNcss+VW4UwIQ5flEbiR3/W2K49DIm7H0Ado4fd7P6YD1CzIkRgU9JhXX3+Mq/Wx
ikOXLsDfGzzwN7hOzklXlH2lHTMP/eIzwhYEo13yJ4AO0zrd3X5OlN9lSYPIeI5M
RhmtPEVrYVMeUgZwR64AspzTvCHrbiY9I978zpUS5s5892VSV5O4pTO6OOud7wrS
UFhDuSIerJccrCqvGJU9E+1vp8PvU2KULa9MJZ1MEC0ta9MmrPrV9hV7NnqRbY5a
oTktR5U8L8t2+j45GY9JwB9Pd1VXNT4dpi9ZprIf5sXN0bqdVg1aL5fF8C9Eumo8
GBzTt1f5HFkUPrF3VxJoC6Kr93Uy5tCwvOIoeT2nf9Va6oNn3BvrKJbKmXNuj27O
LxXQw5/eO+Jpup4ekokPea+/PCbgscTeyObbPegDOX0SlNvXyNMRU9Yp5yI5OUeR
ILyTiuMenhl7e+8beuLf4fDn+hUmfWa2T43MqyHsE54mw8ZhKTj7Axcz1BIIDZdK
OfUSprvi59hACUTu8oYXFw639U1wzGaYkKqHQ/pbvSMCJB7cf3gLcI00oj3FNGC9
KGnQjLvzU8w2visEo32jzLbHgMiUvbt/2FGnI4OP5C3mn5tDprXzU0nur2hINoT+
aMQarU0twIAAzAEmE901oR/iwg2Yh8BSra6OMN0jVZ6YFUZ8sjWayMcspLvrzQQV
UgpfhE6084xPNKbLYZg+hDDTkdtmBogqAltfsvZoGIUWiKfrzwBXTvP+xNDr3eGo
cZ2+P5dTgymTtgFZjzOqE60/G7YIqILWHRKc0xiNq5p4oHZF4WXP8Is1/GAYCUvz
lX2MpYP3UXeNtOhcPwwX1PaXyIHU/Fgtd2HH1IB7my7P8knhacJAPk5ehA5LhGTd
5bPslZwOnihSNmP9BLm8pKRMh68GZAa9n+a/VNI1Nugh2aibVnqwSaIUipAmr839
FaVJleP31YzHmxez44PqVNWMQGVsAhBZh/Ar3X+WK8F7z6EjmaIqAPm+vQMLDJYR
aq0nYCbDkdUxHmV83ptV0PksJ7xzifxkdufafLdCKFbD4XyhsYDQFwGZhMThY9Lg
vEOdDS5Cw+t9pZrQ6VHYBL3xGOM4hQtEN/yXYbZK63MzK++ZIX3Fq4IT1dwi7l/R
pwT4IWcLWRoLSYV09Jv4UopUnMwDGbYUS5u7kaaaUu/P+W9WuilspfFIAk+6xsYS
qptjdNYz6BEQQItdxMBwjmYGCSuoWQixM5jWowVT9pMSMD4PlSwH7BffMob8f9bM
yO33VNmgXepr4HnbtpBSW1ypmqUybNt4B1piy0VyZdwhsweObieXpwNxkJM6iNu8
z8lDuYkGcZ6eMC9+f4aTNEXH2WWYF2PePgxhHUnjmPQOkF5AKuVr9vi3+QXpBxHK
nXItwmKmNGJOMC97WxnUPNRmXkueC7ClDGajOfwHtA7IvUbQFcad4ZI6xFoNhpQK
BC+OVqSZeRzuh4pbIQ3pvysbdsu+qanxvVLCXfzEQS2pK0NYsICMnWE40e3/MDNp
+Ob0/grCH+G1DN15dV3xF51P4rAS/23mUqOvU3uV6+518Zbd1y4UdIg5Sj3tsUtl
mENN/mpBsIKyqPguIXrcYTnDwhTEvxyxlqLcs/yTWUBpIWODztZtqFCRG8rxWkW+
aurpFZjpKkhJAjJ18cZs8ZFZZqDwLmx1gZobJcb0QGTpi/idJr3t0Tc5YQNWU2FZ
cxIYZqGK6/wxJ8erehzVf2kluqqXI1jJcbCFsrs5PAwmTqkw54xgeozl9J7vHILA
OsfNoZ1PIm3kxuvx1y1uNNIMpGlI9UXXwLXuq1WmMXL3jETzyqvsFXvpOXHCRMeP
6KXq0LVwuNl775IFmB0FWW1ZilfuXdGMva2Hf5I1k3nX1klzFITv/yELU/rFxH2T
fK/BeHR+ou5wCKaBgpDXDGy7eX+d0Z94jyOdSU9OpgXgM1bEr2qDYAm1vspFnUaT
3wabdf0QIG5Rr/1mN+/ClRJqVAf25qzvvK6SHnKe8vK5xdjD62Ib7IxJWOULfc1+
MjEzLuPdhukKJvL7pKnfhzfiEWXkiVI4wmK04imSSiDQE3rbcdB8zAg4MNWkrkch
0GKWantcI6zuaEvUzca90V9eXQanVV6DsGnjj6vC6OhnGQxbiiaVtd4KKPtdHn8g
rT7I3BHdZYsFq3Y5aH1zwztRJVDZx3gBIAu34LMTxJPgG8LAaeOGr5RxQgQbHuqv
s4D2cKRSJhfE6J85vuhkclk1hndGpTg+qL5IdW3GKfnvrwy9381sP3b7CAs2AI/w
mZXOZRZFtIBIObxgyqZYyS+CX78vWe3VMLKyBemMBvOWwHt2Eb9P3oy3xqVM+Ryy
FDBMZsuXk2YiBgS9kpuJzVEMMNDCtSwG4TrjZZgOTsy2WdsJSeNM1rFDaqnTNJH6
ruOh2LqMAyvw5cGybqBqgqwt6vLX6tMZhiqk0fIeBaWOHxxg3hE3OHlVCccQX+Xq
ceI7WxmTLh5d6obqS6he7tB1LWnx5TkJy95LrHW5d2rDecGPea1cXnEhWyahaUPq
GANYLk9j96ifSov3NE1x4ChqwY+AbOt88Q11iYtPxsVMH0Q/dJz+y8X72FiUi8iM
yenzKNP4gnb8ef3X2yeCE/kIEignBZ/Og1K3E2Xglpn2sbgfGHMFG3jD0ZAUPylb
ya9ukX6oM7v+uLygrw2v6iBqPu/DULfs5p7bFUmvpnfGjn+uwo+rdodZFjVT7BCA
J0DLgCTuHDSZZVTry2UARmkOY4+xgZvb97jc0qY94yGgURHyqPBGBC8ArYP71p2T
VhVaSof3kZqnsfDnSDbnWyiyvrHTUAKpZmUPkdrBMB+eYmYeAWpJO0CfsQb9ig1Z
hsDpmc/azrywe9Ne9KKs+rAM+e3NbevpZBhzib3LOyi7BBm+Lfz6qmvrRbMeyfYN
LqyDnj4I6VpUxOIHHrh/MGfje7GjKC1uCfZO9ECA9nXKmVJJIV2is8FV43Xm7QI7
LA5V46kYop2g2TWomobys4HVd6EI9peKYSZqzMiacw+Ai469dzJZaj92DnFuAETU
PuN62RaH0XeDKdX8eOp02X49hKi84BfFY6td6uoq8qS7cu4wp00YG5HPE4evObqq
1tsPEPHfPxpNN2qC0Ja+5RPykzkxZJ3ZcD/YOrLyu7ldWl1c02SMbzwiZcglZ0Bs
OCqFweOpuA6XX4l4mOAm3OpLHX3M6HP9JDzgGoS+5iJrAXZyPlNHARRqzXhvhRel
tHVACIdPZUn49NkjvHeoENQ7p25DFr0GC2/7PzROphEcEahLtdlzWNT8AA8EvZ9O
u8nhDx5VPU7Sw76nDQTO4qQksOonExZO+SGfMlbjdjn/hrvMPYol5iVe5GgXRQJ2
kauQokSYVi52OSeTXfLAoMq8yZYoawW4kt4VZ2jABT3cwliJemksAGi1MCrn/EGW
x5K1+iBG+fOOp082fxU5CfRGxbzN97InV1dCdC/bcH0Q1ut/WMVtqM3qEMNb7nLA
TEe+rd6yz3zWKt46hkHzDH6ySPQoYPSNRH/WebB5+6O1rbNzDblUjrdAHZsQGCJO
G0ljaU6uuAFTT8CH1wycOY4Ygtyi7c3c5JmaC3xqQeHLwsrBnU5uqQpT9VtccdOG
cJ3QeJ5x9uzN5MJ3KUxgmG+/FaXRTXwB6JG9eV8NIeCeyjW9iVMhtKsgchFQF9cL
D7ffHc3QpQBEE65rFMEpp67Nql29mV44bhffil2tv7kygwusp4ynTy5rKhSohx98
JKeq3/Ze/rhq9tT67oWmxUvK6t7nQupr1DuOeeq9yc0/UBkl5vI+m8UUveqtxYx/
+RShLDoFF7xg/7TT9oseZII6gqa4yVGk+QVARjJGrPFUKXgN0c/AtAQ/jCFy+6wN
BwwuZtwFyCJlTYKr7O9De7RMRl11aLS78xYoSBynZTJN1d46iLMYOpr6OboZiTpe
o5Qoq4XCP9KaT15AlILworQoG9mtxW+H0g2qaNf0xJz5FDFEdlyqbnD4eUYcZHOT
GALgnfud2cv7WA6e5oCp2dAXVy3dSYaAfpPVWent7tUfoJS+bQ23nvOqXhcKdwKK
32cE+QN/hIxS2+pWo6tPcA5sWteH9xkjA/OBb2csp1ABWZCvlpTKIg9bM5Q7uAGf
I2h77TyrM9iGY9lLeSi8ZMA+8HbaYPfkd0ip9HaEWs7S7h46EKQU1/vNw6/f0bg/
kdWgRKVh0J1p/n4XYGSzA3vMzRpoQU3jELM0itpSIxdBKlHwxKG/ltHSyaAK5vWi
Cx0iPXjyoXANWGds5l/7r/Ml+/Ck0sebE8N+esLzvt/UVTArWcBpWOqnRlgtCPvl
J+wdqP+bRcMpoCIK/MtQwHQ0brhmN88wieWJrV2NC7XWDDfRmjmIsgT6AYUtbN14
AAprx8Uuby8QvVQtZ8EozszKkfykNgb06L/PT5Cf+AJcWRWHgSdtT40L88f5q3dw
Ov0o6ilegqDr+NSXRPksV/cMBJsaNOqfXL8CCSr8XL69ncihRNWUODEF/J0z53Ty
umhKQ5cVN3iIvsLFM6U2rsI3La86i9xrefiNu6fRvvLhcFNzz6GZrHv1K76ps+M+
2jFmqI5eVBM7kLOOtqIaW2SM5IANDPXZqNZvHGSna3nugm56FvthXcRSnD4PbZ0u
bYk/WjugFgD8GrnqlmHqtopzDNTx6+EMSN8p6BA0zx9M5G84FhitsnWJhGSkNNKn
kkfmQu8+H3nc22X7kh/2xhYZYFgwFaIAOWEjAI1+4oWDdo/Gc24p92DmK/VaX4/O
D4k1nWnfG1UqKVVRZ33Sjn67hXmo4Ri7EsZbHAgaiNeWHfmfqK2oxwY1hGVVzjBQ
BG7Yf4QwY0ctimbliY5bocVJFhxGeWFClsvZhbQEm5gw2x+Krnkc1wQNo6iPa9W5
nMt3DGYNZ8yJM6dAS4Xh0VvgEGqI4ZVkKSjZtj80ADNC8q9hxvg7rivmopQmtZO7
cZg/O90q8ON5mO7Rc/DAcS8G/5BUt7zcBQd0lDxxMgkXQqZ3VmkEzZMhY/OAkqEd
VAur1SKA5+mFvqtCLT4iYs4sjAyXZVcDj99EChaZkPIQATn45T3s3lYKBsgWn5UM
QYEsohZ9hk6JLkCm5WNorqCdYzEvpmpX1faKO7J1Vxx6O/I6IBmjthSix8wy+MIu
XB8JSyNh/4fSqmU2+HMNd43p9Ee+ETH1dVStddoXGhirPQHP9wMfSr6CGVgfIX4E
YComGKOoVPOQskI+we9CusB2hpBPgZAp8DKvlFJTMxSL2TH/gd37jd2Wg4ofSaWe
HsDo+u8dYpvvbRDJPX1AVmzexsU7bZ4Vdqkz3kccuDsASpNh8dMeviXZO9gaouxo
H3fw8ymPI3c7KeR0A1FJWocdQE+3KLAHuqJdNzVMt2P6/p1xJ1Ld9wf34hNvCsYM
+CwRJCHsYQC7SesQEzGB5hHIqI2LQ8+v9oim7P++/Ej11A6+5zTrfMU+kbwdz3C5
6fkddx86AOCSrO5REOWKvCcty5E5KHfReXLHciqEHuTCMDcEsCeRei+pEt+Oxtr2
JMJZFsKI37GsbqkgfXdiUIIPW+cKhRgkXgXqPQBWFODmwT84aJliZi4GM07aqnqX
MI9SKmDtBM+CsiTzp2gGP+4psfPW4Yk0sEGU7OAtBuywGDtko3LjYf+7x6PMF/l9
wBdVZStVc5McQTlq16cCOmnLOnfUVNn9MLl0YNnbjHqWts+rROSUUVfxFFCsXhMK
1MejeohfCMkfxs1U0Wd/gE2LCN8HNRKxM0xiVwj8g2+NEbxq34P1eFEo/Ei0PzkI
Fnfzcknjf54/FVY279p2PTcjVs2a6SUD4X970OkmCnjzQbqeERtXJWqy7FCASF+Q
hLoczULHk/5r8uUxRXaBFDGshagnMewdOaWlELZ7QIYR4jYd/vcM0Ftb4qTjG+ew
Oev/eT1WmfvZDRhAKkEGYoAHLvruCebkpiZ5ahGtaHTl1qaK+oyJ66d1fzfc8o7S
SRTcrlrmkmZXgM1biZPM7jp7M8RZu1xzsczJCgTj/N0LrYK5Pe8GL10v9BFbBRmW
1SM3M1lyNhB1zi6uxBaAhFkDyO0rrkFMId0S4QwCa0swlv0ka6RLytwUILIvSGXc
D1b438o1PSj4KtvDnRDr+B1uH1KzKSeErKGXOFnNBE9p/NJrSTgdW85g1zqMOY1T
t1LIcz5emYd3q2ILJ21Pf9mE0+vsGJhvBjsS1BrVn2QwtBHLKk+dyHwels0xAa8m
ValAQjws6NCXgi8eS8jKfzJSBJyJJwOZlBIAkGZtWBF8Iryy5qsRcxzfKuIBZWvc
jSjpMHNVNoD3yfvusY8Od6HKY9juEGypSZ5sL2mCLVi00pXfB7Xc7mUaEhcCigm6
xhIMLYug/qBUI8k8Jt8KqYEtsrO/wG7WAb1divhIa4oaZgLiY+yTjb6/Dm8VQy4V
Y15yOIAZwTlAY5chRmNBlDAmlGiX7mnGQw0VlwFGyQ8Py9kh1d3UCRv+sYfsgU92
Mzl8u9iAVqeC0JrdqY43luuPa9kMadA61+k8fWtWX5rD5tj2WQeXg0BJ/UFwi0Vh
0fh6jyldhpKBCwAtvjUY43WsepTqBuSnrjFj8jSGdvdfvhtj1Swj0delVQ6nZCBV
YG9uYLZKxAL6wCge9YlNiTA0U4PB36DLeIj3iV2PxhFiRnzSp7mTt70RV99gAHtw
L08vIidVsDsGnxJF7g/DKS04Jnx2rVy12t2xOXIOwJxTYIdGimDmPCZdVj00dXxT
pNRap9scLlSCfhhCuVIVi7Qe6i32+6UJSL2woQLV3eZCVl2ghpv6+quKrO8uPAJ9
c7lhRQRvMHNOA3YvYd9BJ3V6hjiS1EjBa7s9ouZwFVh6IkmOIqQTOqTCBs9TA4Rw
pj0SefAfoiGsbfv3ch2TNk+LmFIfKtjcazlxNIMSxBBRn5nbzL3vKuFn9D+OVuAo
ALajlNZ6ocOzbR/p5iFPvSvqXr1lf+zoYwtgiWHKSCOmhInYSeBUBOR0cUFWR/5r
OangKprEXT1LQY8+DtCwiKMGThFdRlkAK6ekEBOdKAyoBCJFUMA5euOdfVZIwzBB
s/f5oIUvWurP/h1gFRncRSGYQV7U2nXlp/+hg+oOpqvdj46UmHpw1l0HvWfwtmiU
qu0Auz1NV/PXNyweCHL5XzgaKMm8F/pqc5Uhv1Z026PxbwiZUF4SIW5SHAypdzcr
Jx6rRw+stHpz0SlSgIo8LNO6YvwG/NryTs62J7McHjrh/RFUVojKjNq2UUXppDAA
3R+iuXBfRjEZQgltSkeOJYpKLt8xRW3alrOCIP/czEvmmk4RiTy2+hk3L9fUMBJB
3EEMCGUrtMTvELTdIGzlHCu+8e1lqDC32p7LwEsWQg5kxQAQ1Ly5SIfBkqHacECa
lfxuRYJ1s9l6XMzp+md+PdiPOneAbZuWmBxH5OiRXxT9o2DMp6u6CR1rORfGH/OS
f/G6i6/ZeYXTjpHJ/qmbPkgdd3mWlzIC+hzf5uX1OAD1r5XGQik1U15wUzctUYI2
4E1jnzClFTPmdgcfT8ZIPMIqDliuXMhhWk1ISrZ50/ezIcN1oTEXjn4OnX5uzWsG
0mQQQ75was41au9I6/pQbdEOi8bThjdvirhJsWGbar9Q2HRz1JuQsiLiT2WvWlQp
OLLE7RxQq4YzZ7HHrKn+oCiPm/L8UbwElT0n0WGAtgXciLh8NFmazhorxxPHirT4
QPsRpfYY9mB1Fr7qSddCzhJAHgJcrGi4K7AXdNCtLLcKJrw6xAFUe+mReG0w3Lvc
owrOowJr1OY2obBu/YUZZeDf2cQVWSxvo3P0ClTjpm8n5a4K2sRdwJUeZXm/zTJG
07K48tmFGHE9jwfIW64A2VJam0czPH/jbbqaZZQMIP7ECnvePGiAfGvtqybURFgj
+AXh2YgZXNNqiSz7JfBIu/X77zBuqbSNSpW/MPMe7uPGmwJQTBNSiWHRyLibvefW
1X380GeaudEtoe4TgAfhdmPGSaHnjNUSZsTuuBD8sk7Rgs6LoP/wCYAZGdGwHBZN
NB6ac9tt6ri27lSwj+t6GyX6Of14YAAVfiDKK1bLcLrXmLfdurkjtd0LRmpofP0I
AdEYFWg+BNSXQWJZKVIjdIzVD6FmxTsuaeBSbYQVHprz1atD9MSbKTrz95XJG6TE
3J00TkvanjRlEEkwjqMAqIEvPWH+uS0p+yA5N2mQiAuU3nx4Gi8LxfC0OrHUxw4+
gsho8da2vIGFKC7DbSUdhgjloAyNhEAzYrFTn2UORieAyeYCbLLf7goi97aWCLZN
oAANROCZ19hPFCHCyL5pykies329Gt6cy1bLXNfF5kUJa07Z1TqfUrrk3GJKbo3P
aaw/hhgqblD4hUDwbKJkncbWscQp1YO8u3RZcAsmPGyuKrRwGEp9F+CLl55/1ZYm
7EJckvKuD1WdOG7DYrfhEx6ZCyNCqjgbuadzqMEiaGPYdVb6SH4ygmdolGO85Q+U
w2B1KI1kooxcfS7hUhbx3JNLqUACOvRWJns/WKjbwi2krdV0x2Ld1comtlZBmkpc
XHtAxLQ12kOAPV1o2OW0xAoTrNQH1lTrvJMnohuEzxmoNL/FdDnL2LU0Wx2l8Ig6
2Tb/aRlUdd8JJBraEGiOJqCRjuxmBAWXAP+0l2KiB0v/rRllj7h+PZ4cpXk7BN12
80DQP76vax+v/PuNf27009EGCtxCXUwuRd/PAsyMqkOMRnar1eXLHWQ5cPzYIYqU
BUHxh19H862HRNJmtJMruSSbCdf36fvZ+TzI3sznAJKX6syqbV+vXrBPJ2f4zqgl
q0acn9/qrvrM14SHmjWIQXuLcsLcPfMGG9CZY2gamZ6w1VU8W89Ud0zPVZ2fEGlA
c0S6FLvExKh5AboxgpBPOWH917KX0M6ulIzSr7gq0IeCdEvPAZKbIP6hUB67pNh8
QI/lCxVEDrjV7rfVDTbzsjVNbqbjl11UmRNrFd1T3IQx+uqKWvGN1npe52ZQKo4S
/f2yKNPxSEgNV3pncccVYagtLgSemNIO4S3B5GqSnGrST55BAs82jQXprgWRIX1t
Ft0KByb564MFtRkUd4kjy9XOYFOEqKsOBeB3X1W8UxtiUqxwfco+q0EUuQE/7Lxv
RNxCrxwPxYsvB40D0aSasiS0YUfEE5mlwMbd3BDL8cfaz2ni57eVqE4HLUBzgUHr
kfN8PZPjPkQ5vSZllmurtaDLNoqmXbqRSkWmUFCrdC051JRHwCgMJNuy1jAoi3Aq
Q5WM+PYbYNGrexY3/780gq8BHqxEboPIthLKcpCpBveKYyzkTxqSlE2dGisKv5pK
gh0wzvn5uI9sX3x9nUG6xv/Kl3YkXsrn6vFcjUAFZc9ALdKyumrVejneVO3FmYRy
IQOamLQrd+Ovc0+kPm0rhNS5GeLLRJMQ3j/h/6z9Zk3uFIMZSPuaJuRXCjGZurl8
DXDB9K4+z468HOXIff6n01whPZd0ENUc/03Qxa3rd5WUhPm+jH+F8WdO0FB1WbMG
lANW3iKeCdvdzCz3bMW3cX1jyt1gDGWH8W81SvCkvA3PtvxmredfacppVnoCj+d7
cFqo6/WC1qfisiwvKCwOOfz5BwLKq9L64/z++aGwHVL+oMXdFLF0qlqgzbZPGEOx
Pw8M4Ai87YwDANldjxClmvaU8PUaN1lsJMsx6yaf55MZBWhOnGdn9MJbgGT+1ytT
WTLnwRohirV6qKzquZbvPJeWyb0+NymzkNubg95CLfOTGuseHZn2DGy1Mp+oMged
7unexuazRMr5B/0IqxpUlc09i2l0IMHLnpiC1i+F49C3FRPwiS+lfCqWa5MrLBUz
dFwKW2nNmkzXQUCstczoNohl7SR2xt8xy+BiR77fy0xPDXuE/FR+gCtkQVC1gCPS
ic/cnaIJCF7PdzHdpAOlNty29qyRLYc3Duw7EPJ1ZkWZjrjNUF0IDBQBXlL1/j0T
uNR2soNdfM4g1X5/2j23oD+kwzdc9zaMzh9nDe0dVUsyAFSqF228bUvB2YByBJgV
XIOyneCChYIyP5KrLEFi3UrxV+ZmQOXqq/3k5Y6itqcgox1XefanXjfJPJ1GIgrT
VEv0lwzZPTnH5dSsot/2VA1S7+uCIOksUxgmIOM7nwx7+JvOBiH1zGWTqsLo3eHm
etyp2yMtn6VKCI/1fsoVAJ8u8GsBzMY0LNCSpTe7Od3LkMkXS3/ozEhIcdCseOJ8
Gh+t8cxSXrGw8oKMT0kkoS5W/QXXL12gWHMR4eAiX+8VB1pax/kwQQThieAJaGvp
WxtZ3DwDbixIZTYo7ZJuu+TclonWO2hY5FqQotro/IjkVZINkzjm/l4Qr/JIxTY8
VcALVbHQWxVCjknTAy2rwKbKg2TvE1t1//gXDAbEwdnLy5FWLWBEjsvuagu2jt3f
vv0oZaLT5//oyO2wJJY2/m6kqebmzcTxsfsYiKBWOzB3HUxivY97hBE5ZRMgCbsN
nLjQnWbQVZrqfcsvTxU/0m+aI+67Sgk2JfcKilLFzG+I6QXyAW+o+cqKtNWLfa3f
lavd75CV63gF5UMnLHPEzDr9jdvmvBOqTq6MOdxmNMVBABrt6JdH6CJrSkO6Xqw3
gZjOHcyuW9Uex455vvuR7ia1dTLNrL/hd977lMJkmQ5ujPUTd9teYOUxoWpiRTEE
PsBEIvhznbxiJeAspWKmZb+d0bEX3c3Z2GwPO905y3IAbuUmmCxXvnezbBKITxZl
Kwk09qE0416O7SJ1uQWAWILhIlRNDMmfWaGVC3W5wlHZVlHpb63fp4bOJSmlN3y0
z8P20J+XDTxYGHvfTx98iq6tFaAjt5szaQACqQgd5LEL0dV8kG6sK9XWsNfNrs+F
Sk2lE8F6f+hD9QrOkKGJFMCGc4KqnKZgAjkMxscxCSfYwNakW6qki/Y5bcZ27QON
7DPv9YQjfh7ZEiKZiRZNx8Tv39/kd1wKVe/WMUzQW44INaYpQWUo70C1mijaZZFM
C9eCmUJHZ+21tAg8ef+gyrMUU24/I6tX49suVVLyXD3e9BTe9fUplAjLRTOhv+Jt
DP+L1Ez7+Bnzby5tcL/1JX6mZpixj30lopQdgaVRE/bxhvl25Dbys5e1OZePb03A
kMQ1CA6IP3cQif3R4cKR7+EC5Eanv9qCpdiiJ6oPbgH/cs5av6isyWOgyIbX4BCs
xyDYwlTOI5p2mBzaUxqEHes9tzFt445H96mujSzKNyWoCKVePFj1PViNsUTFtdKA
hs68Ts2oDIrFwdD88GSFbo2z1sXwRJxxOo2oLuNpL29AEJb2cj+nwCKbC4lBJlkm
pfSOURAUQkE9/Y03x5tEy5kh5qko0Lkmtu4QobcJI4nI2Htyr8YSxHYGQXvn5YQr
+Hhj5Hq4htABw1MypnXdLhCOlwqrmtrO94lT5aw2FcN/DxLnx3+WwCnh+QLGa8YS
dHvnbBxs/KSpYGIdiRzR/f7bKgvwkkSiC5NiQbq1PtshiUzU6JHVVETmmMWBtW1d
rKuplXYIOOZcUSVjRVbR9aG1KhIJDkWdbnbWrP9u8/B7rPWcEVFI++3lXZwFg5yY
rJp0SgvZpkKplXxaHIq9eBw7mXw9d5sSXCfu8LMNPXdKBMcb1zZJU5VKp0Xq6WP/
83znDFGMIfSWfw4Ev1deN5h25nalCu+ZkShxFJf6kwUPyO9r/6+RBC+WR2OeeUId
Mr2ABsvzr5AjAJlEsh49CY4ya3uyDVQ/BBGH0poJYwcblKXSIPwoKiQuBmLo/M40
d6HjvrFpHU9UIzTYqPm+/negrOV9XBp3OFhlgLsOnN+xcv/z56XXQRW7e+1LG86X
Fsx0iGL+8TqOvNRcSlgRiD0VedeoyZ1V2rgMKFsSwNdpO90Z6Bu57adnmiQb1dq2
UZWj+SYhqzqp/D3Wg0TPvoINm8oJxI69wPuZY8TTbwSbYw3EA2rAqg9BflrjVyVB
jsQWHC003MyNx8of6LUF3pQjWqma5WpJYGf0046t98Ta7e42fcLo1uZI2VnnOwgW
y0hCsn2neugXsuC/xFikK3S0pcSytUc3/qSlgIzYW+SpiX+W153KKh76vsTzWN9R
A+TgkGQQFdCyvX/9fUd012YsoQhc2o2nsQy2o3jDo1CsmRNANPXlvjcxTA+xgXlY
DJQ7JHbpdIMUQuWO1QVxj3dJ2FLo9oP2RAKB9v2tbziP9bicUrcf0rtI7XMFCRun
f4qwN6N7Pt+IE3LuENm0m5mSM7/Yxr83CrlyZSZOwpcCEBPb8HsWVX2jxKdqzmuw
elBHhR8OUn94E+/junhVXrCBUYKxsZ2HFZuO0987s54B826RK7+0VfpeGj/qRqze
QNj6kadHd2mbnv8+ToPx865XtRTHBEcY4LCmDMWFdZOmXBed7cT7MzxBgYsP2Wfp
l0XxhTWnQLr1DGUce6o6tmZcRrv49DWEoWtqef6wgH75uzdIw9gH9U8vtJ6T4Ptu
c//eJik34JgB3BZQPXNm2yk3OOubBSzYDJ3sGmwbrIn1mhun7ZBHHoQBHdDLHttl
sc/yxuwuWB4Yi6+0nyScPz+78KEfimHHO/u5LGlhLaO34ie07leapdbm9GLtymOc
/ANaxgUG66DwuRiOvDq4I7Dx/qfgHc4lRqS8AMl+dkJAb59inPMAXYI4mTP3l1sX
wEMwGxkvEN1/Mq5Jh34GeCW+sa7a5OiWZJrwbfksLnpRR+y94HkgvSoqYvTDTvsT
vHfadXD9kSQTUu0eOap6WhNFl38KdNJnPT88BB6IG+tr7MMq2xHDtIHnfWjSEDbU
2wHA2qB6T6Tg7aot9zUU+7wDvP/LUjwGzmWP38YcXzdhzuYK8xcZcXEvyD0w+o29
E0HoegngL4GvmQTm7EW2JEBT5aURNGJ2+JFj70B8YMYNZH933xqTCgYo/Oiy0UjC
k5LYgIXltNdr4AI0SQRifwlJa5jfa/vc+jmaxOfHWSLcwuCF1hOyUd7imN6PEks6
iT1O3EGBOB0jrfHwisk9ZjCW11MQX0OcR/4xYPYakpvvWuoS+/VovI1QmxmWTJ2+
rBQ5oWF/PgFT+zi6Kf8ZqrQUKYni0NDZ0pesQkyWPESUVvPWkHcp8vwSaWunuvEK
1hdznIemPGXoQCbNjXSgPkQR5f39VSu4NS1XeK995L9D4P+OE9jtRVTW9e4XvNvP
yBPbdOrMdZNwNGt2rhZ3dj01f2gSChwS50QJndPKiEuLmrTf1eMAx3xYo+MIhbLd
uvBFOVRF2RA5fxxiGoDcm7K3habBnD/x9rFdvRtk6QE9MxI8ajcoS/xzLtbhc4yh
j5tXvpSv1l5BM83Yy1DVX/0wv/gbCMt6W0X7zIZfq1S0mRI+JDRVY9HcRwdUTWGC
UQoFZpi6blhnydPwwdZPv4h1h5Z6NQVRzCZHGjAZVWZR2g8Cy7pu7bDnav3agjgb
v0Irw/4Tudevz9yWHFVf3T0cg45bwjHHAbQwA/Pr4FcDS1XuHd6EwOx2g6WR0/CX
hBAlpLw81N242YRwiZwrwbLiDQgDHuinn9ioNqK3zFTMqqLo2HnwKMm6C4hy6EVo
vy1Btc1sFP7a1ZFpTJOdtYj4SS4sTp5oHQ34kv6w3fXT6voPrGzO2+P3HwOQatCI
+dQDbA8zu6AwMH16CK6lYCct3uA6ZPagMe+qAYfZ+yfCyGdNgKP6N4aHI18Mllp3
ke9MgjRnf1uhZ/2IG+ZTinXBL7zpFdkWLLlFE25fHQAV96Fjz2PAwRLBkt+9+A7u
VR2r/JUGxANCAeLk6rWyFhMS8p0MHi95mhS7pa4mTZrCkTIOHzgv1c+2wDlWaGLn
6sWS4mrvgB7RHd+soOUsLBX+nAlmqeiLNSkFuVSEMiT2Kx6hozlPlkh9CSNPGkh/
pLhsggs+oQzSJ9ydmg5IaA3JOg8z1caDkqeuv6QYsRiwmA5IURROD3kwSaAZHaGN
9JxkI4Q7idzfumLr+YMjrCAYkJsFd1rSDgvj+TEzzaXlt6lLk164Q+LrDh9CIcMR
B3Ud4AfjdFKdEeHj+ljU4EaEPWyZLF9R+nxS70DKpuEhG6lCaKsPZYEbkUEKO5hF
sHeMIchkDAZ9VXAaDlbP8wqOBxEg8637Qr8QkegO14GQPIUG8KnlxBJmf0g2V+Rt
hktiII5QrKlYu+Na+iv8YeQPoimMAA+fw+dOkAfoc3gehrnW9zSpSppPjSRskGjk
VBrSKRiwirH05vrsU9ltMQCt2a3iTI2RGKJcevBg9l/qIqI7b5dSxR4siKLCVGf0
LtsYBrEtvCm/MiEvlIRLHcfZLyTQlbr3/TNuQeBfTqmuKsG69CUZ532IS2mlKATB
SaNgztja4EPQFzlvIN8KsQRVU8QhOEzf5jPAEOdzpqmQtCfguDLytNZIFJSyg9Wu
pgK8AlrYIMvcIez1haDCaBCUNx2C3TwKud6EWoCEAbXKKJvoSisFNjF9a55hBvr7
JtJRW3y9DlzX0rAPAoDYLX2WNbhqcI159xqXOMirjq09GepTl9rjScT9m6b+TQaI
WwrYkXOywsm0QfD2cTkEEN+RZF9Lgy/eRrxF/5cgdEALnGeX2rCv5wS3Ix9aaY2y
S/edfZLSXoALa0HWe1z/ntCquBvNedSM0L0AhuesgrgngsBu2AazZrNash/nE/gJ
M0g5kAdwds8F5ANXBnr3tqdk7VCesv9ABk5vQOFPytXkf7ppNiWwADgVK9+H4D94
xCjqLyn7/9K907w8iBJgMbCw9VNgMI1QcN8hm9VdtloKJKTyLQKtAuAE0Fr5o1Ao
Zv3wf0V56C/L/NJS82Qdp8yC74Xo/xMTuaoXGjPipn8vtbccwF98IVJCQJL2PNYM
AIUnMR6F/M4b+RWfV80x6Ja5OGgzRkX0KspSC48xcvZtLZ/xaV1nak4nL7zn0ZMm
YFTC+mcf/Bjczzv96yRTkNjOjgkslX9GnBg9u8m5O4Ck6w0pXwWuA1rXzDUAUNde
fauvAHPcy/KRLp/NXIqNJVgToc5ZALD75AkF30b+lU+lP9gKWKzqCyMEhWQenm1v
FdyEP/26NT3u0Zpe2VMMicEvnXVVmUu23XP0hrzd6QjifOB5W6ypenMl9gRdOOg7
jzxxWgAzM7MaYAivwMimPq6Nu/BivaWzpXtShJ6p4Vb/i7doihYtr+qlRucjb494
eEgjRfWleH+8tcPnN+zIF7s77RxCianekn5rE7X9Wi6s9kDvhrvSRCWWvwcIt7Ci
mByL8gSZwdQk8iNknXxY/JQUFjos8SJQvv7HGcC4jquoQO7t+x96GWRzZWVnhVBS
68jNFk0DNdVcLH/EICxJK6riCjS9MSyKB/VY+CrgD9HEC9p2iUXh1K/p3wbthJyb
Gfu8nsooMFTT1XQtzMclU2ifPdmhfYsmC/zF9r7xDN+GsnsnuRyXcAxDSiN4tvdR
NI5T0G4ept3TYtbPc751dq7GHkexdfF39LrljmOeSwXqgJ9Tfn6LcUUrSjVhxYJU
cyVm57CYDGbP66jcoQDm4GtnKGsKuBclnjQzjNWxvufDNUX6w4wJkFQotqqSSLwC
m4NFmYc57wyHDkTgk97k0ZTguYerR62zNWBPEM1Nrl05tIcV3YoKEnKHLVTzMGdW
WkiAKYCl3RLk+0l8iGVLXO5vpUUNYV6JyNONGpOBRuk0msefpymC6xYH8w0ALeIj
DAE9iTv+Z5N3m4lnZva+c3/V+iAc9AkcbuGVuY0QELuhAom/mMGTRQwjWE+SAS0j
kOp0SPOsszsYRleZ3qBTRtNetkPEi/w5uN9NS/tXSJ9RZlFko0bVdkrVEO1TfpWD
cyW3nQ8y7JykidoxZChIAccCZV4BLJo0dOLIEYx9XIw4QUv7oBDWtXR0atkIuGDk
0qUrXRwCBNfBUS72oAcDWV5UfPY/lkoTTHRgRrpso8Nwd8OLsqUS3A9wPbH6+KyU
viI4Fe0dfD+fzcAosjiaJgQIUn2fAOimZYNs8AgLdWs=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
toM5J1g8mxxqsangkBKKibCX5iGUmQG6AYiXAwMVYdIltWVep90JQ2YVfqc7rERz
LDva3VwqOFMMp9jc44IU0flWXU5J5lW2X5RJnaQNQhhxjW3rWBLdAfT6ySh4sviU
2JZYPlmgmrIE89nMMSH+WGpF7s4Tt+EG5mRzg5pGVMlhGUIRwjsZjPBxh1RsljaM
ifgZw6qZAmSntwz8UTGDU+3k7nxSkJnakEKOzACQXjZXzZoLMtUiqqrSF2LFzXUX
rK88XH44oE4nLuL72swNZ91dBKAu4I6U7sfdP6pbVnSZitRdzotfyMAamWG/v/ue
snZO07e4npictmaecROAqAhH/Pb+f6balxGSfXLcThn8OmqRWG88SUrLnjvHDJXD
9CxHP8UmEBAKEjnVj4LCmqH55J5S62OtDm4GnkWlEIkiiSJuXg/C1Uw+nMpHFTod
XRGYWFRCsSS76bF6DjZj7ZOFngSX5Gm5CYrWzHjLae58DnNfOMsTHzuakI5Yztw9
aydXlQ7xyfW8mLqC1D+KYtyz7fcBUsDHJfZ/hTb3WOIDN01+Rq9TLUz3ihwZ5IYo
BlezSVJ7ATjDPXqRJPNCmRdPePgqu/kJ7tA7OHceCtWqwZj/bxdRmapAAvd6P5rp
HTIRw1D6IIZxfDc8Gi2OcNINPadG6Xd7TMV4wCxSubCUkVXzVe/hvuh2u0BBXCRG
VKgP2zJdRVMoKginC6WqR0cX/S0UrGnyc0qjBawZ6HHu0p1orNX31E896l7bKdcN
/B6O99L8V7DlYF7w+C4YIi1xZfjD3ccvBpwW2p1BlPqQrQ2gNEaWTzeIdLSmjzPb
/rQppz5ELT3eNrsAIZ0h3/UkdQDorT7gQy+XFsJZ96mUIcpLdL2qUM46LPYH3t62
3wU7cC0piSlm0+hLwKf7lZE8JHrLlNGZM6pswpFi5KDqy8UArda0p6RS3auIRDWd
wm+h5R2d6B4H9OsgQ8KTyBgSESyoaHjd6C0t0rXxXK9Tc2BEII9zobzTkPCskubt
4gig38x6ntLeHfgzGdDkmKCV2BjtDUaYrB/lq1skk6MjAGmtso5nC/RhaNhdmadf
0Ghvbla3pCSCRMCbhajknepT97PDnZhblO5moJe/Ur2YFdhDHx66l0INnUR2Re2Z
SkbXOO2u9p7ElqkiSDvs3ZC63b6JHrDTHPG2Nv69Rntru8zOmEtPM4E8x9rk/Llb
9t7JKZ/tNljBKVDi1/uHN6a3L7r/fVr+WWIfN2CNRs0PoToj3lZIXuyhISPQfu6D
VaIcWKQW65l91c2j6sTnb+qIK+IUEsvNn2iw9/JMIgRl6VZnK07Lf9nGwbtZ77Bh
gufdgkCVI85z7sgM1gMwqlKqWC9sSXYyBNZLCWXrPRogzbTbYHGycGPWI4suvGQQ
PY3AZ5ECHAjN9YiPVS+cQbtZMF8iFpgxLWn62lBWSj8vqRxfdShEZJoPp2+aoRQj
eLkmMxifIEIzQLtCg0JM7lNVXcwPHiFBMyTGbZSOcsdofc/A8ogKHyw0ABcl9XF+
KHCAuMQItFoU8JmGd4o0zKpeDOnR7l8YWoXa9tQWxaUiCRzbohK+636Vo9+GjJXl
L+sI2pXkmJT+TgpGgZdZPP0aXHfrQeH07PO8CvSHWdJVVCifrybim0uiRWj8FqbV
/DpBiLWd/Rdk0prh8iHEiLCjC5m1pKNkEIIUSjX4m5yZ0W21LOEuy98zpwMJfuvo
mFGemNvTICvnGg+16vv06c+i4txlys4HCXiLuAZfFJHhsIF5nHMBLTzKQcDhYRdO
u7IKBOyQFTvZLiXOmjlAwZfrZDBPgdSt8apXIc5xwpNTlem5KCicnAnvc2ddkCrf
trxb/kzGjTkQnVKY0j/kdaXNGKoQ38u4RHu/UJ8sFIq8RF1YjT0u+KUzbfkxpeMu
ICo4zJ1Wik64gheHDawYRa4wMqvaehfUaI4Fb08aT+e/eysrNgkXOmcjzoK+wzwJ
FAVGoFrFqJqaAzMiK/GKrJMOYL2B44/wuCSN+6g/XriEPamxGsW8534MHVzslads
bp+ez92A7V98Awb6eCNilrOnS9czKtyfT3rdr1sKcFn/nJx4zZWXcP/aDn+Hh/2W
/n9htNcJW+jgUPwQYYq5u5kfDemcn7k/oAjWJ1O1lYwh0vA3hGJ5MMsy66i5s26r
pDaYUu6XLuvvNPc/WUi59GBs3dkcbsneGQyaBdOAbTNy5r6+MiRXTLe1FLsnmHsZ
Z7+9zPX60Zxg5Ihz2zFoZNSaP+ONNGexqa7iknYluTmhUj44nwPDZH3RXjVQE+m7
BNJBBRk96P1AX3mOHODZfBGSF2TuuNJlywpCzToH7gwrnu6uiq8SiMncuyCUVQnE
lH0W3nTLcVEvE4Sa4IHQbNFYCNGSZ6iipXaWWMvIMu0nLymB4Y8nbbggCbzl5zqT
qf/V/l3NhxEpYOUtRQjqYlSdQBzqzGKJ0QlfnjzTFO2lgKu5wwHne6TWNtzuUs9/
cpwN5oJfxmdgUqbom0c/YTHCC334r7U/rBVV7O0fewwndgm4RSU/MfCvclU2L4LD
7XcWCbWWNXMK7DMGL0iMcXQ0fuvBxnw/rKmJK15+K3FWfBqbxUkJ5/YuaoW8o8aW
75pZ8R+Ac41ai9jKx3orsAPNsm5xM53PzrlyLWqbmaEIh42H+5PDb0jxXWwn8mgW
qu546WwMmwNnx3oi8PmhIZibPfLV+uFEFeMNMauY9HzVUdKAXfJvt35CDtU/ZrJs
yjvA1hKkCZVseYwmnFDc4hbE7aI5F3Wy59tdHhHj8nfGvbxkeu8vcHUTupOCs6YD
6fun1Rug4yirLmmE583lWUfdPwkWb3HVXpAGje2he6EXUf5XQCU9Ar4NAyMvC387
XpaPdJIwyMaT6t7ZERO6DEwQRm87Y1XXvXk6XmekS/UcXs0/deHM1eDL7BVQwuJm
ljAbiiC4uj/bAo8mDawC/D4nCrWyJk7Y17dmKosMKH9zRYLAc7urA+BugVeTu/uj
3HYW7+6HxOuruwKaBpDYql5MIhv8C7j/LJHD1h2kD0sRosvGiXHPXzU2/B5L1Q4u
3nuLeuZ6RGa0LwMg9jIQYrHVuNiQGWcOgp0gRLBXB8o97YsBjhNyjXhWDsa1rt9B
LBe3VbQGWSLUJC2ItmzvUXO+reXpIdz03gUrsii8U85UQn6s/bN4cwufW5xzOD2C
l1ryju6LOqME3DWng1VSfzYlKhLfQuL06iV1ZzwyvvZFutBlSJKeAbKIwtvbVZsO
vaTG4X9ALP2IZkmjqkabJs8ffr/Pq+r4HtSSfkbpose0TMiSulJYypqW0HJneVda
QoQ15PgkngfxGLzmRTI6RH9eGQfVwDx4GPnELRBXI3OSROnLjEmDamKhSqh4QxIW
J2VCawBaXMvsZBw4E3z7ndgRDmnqtvlRO7sEmfYAGqFtPKvR2qLNSLKgQlzn8Yff
SzKByghW84oYf/5/4cJiKhUc0/DMJIeorjEaZuebcjO3HFTLmWz/XPJQKKHV1042
1KQjTx154QfatkLAKxINJACXrvBZn3M/z4cKnYulqpxTeHeyqRrqfk5vNP4bBSGd
6fdLalPCi8OhahTlb7a16/29dWBzqJ5DCzpWYiSYfiQNJSAZ/804qFWXK3UFInmb
5r1nhfH/fikES/57bey8UIMXbaPtdWAbxPLoFQYNkDwf3px6vsx9MLWgZ1fRLvBz
KT5tvHxBEAw6D8vsPJb30xczAzPXNO2khdug4QkQh9H/IjGQBua1zFX+pomu6sTB
tPczGpGDiLmlECqQeE7vlgydlNvfDZf4naGftl5QGKL7o6XgjzZ6omNxA9EpYdSd
0XLSfnaABak9i3RCuHXZZQy7bdrwfwFK4LA6LXu/8tQPJ0J/cWMQw+0LCtKt48bS
p7OTPbbGBwAeH3+LJ4XgeyCVp4We6ZotVas6Ds5ELkuLCpMzgNevYG0xS58RusMH
MXnhKy8lk2BjRh+uUS/EiFettpMcWMX3QQqQXV632S1p9m8ZvPzTzPuHvF0GuUAB
eAPik3Z3oyH2TpwQ9L01uDBx0e/tCXyTbe2dDo19CAvtwMn7xpTjluzCW1WOMdht
d3P587VrD2zYEtQrrXGdCczNJm8ig8gyggd4WMnUknIc77ANHKb+/V0JCNeDmLqT
UavZnO2OiwkXUi0iGQSWlE9YO5RnWBXcJK/ZnR0N4UlpBoCGqBrQ20v7fxxvBdBr
0LfSWrF2kZFpVpnJvzVyzUeNFpMvzo65uA4TJnuwSMrdoYgVYObEK6WEYlq0zE3j
rqaT+o1Ebfgz5qCLY169ybeiP7TdJwg0Od5GUY4zF76nxZBOUjbkvbjqJF3yYi1i
DVEAwgnDDWWmAkwhoUhAr95F85vvFgBDVFrOUkt2hIuHU1D1EHFbgp6LqHHKVA7q
eOu2tbjRE1aKHfyakpZC8O7PPY6CX4dz8iqadbGMKzpafd5qzx9d4ENnZ9D/QEIM
p0VfD5wQ5SED7fKmrm2Iu+xxzh89IxLJna/DoWuYhKXdtluGt3dKuPdU75I/GZBj
nqjv1S6lliq7Sn0ZhDH31ayrnVR0Gy3de06lsbeI1xB7nYgvidgRsvsXf6R0tEeD
3wzPOQ+cMwHPJKHo0cXLitQE30mBlhhaxEROlOIjXedEUxCUKcYTbubK8myfZAwR
JFWo3sYrnkw+HJBAASfC7wTe7WdtUxRDaopxZmz58iHj4uYi6+Azs4owyPwHnZfD
bBwkOyEUbvW38TEAwDOXytDO6jHMeEBcIHl83R9Stp6gCu9U+ZwkzrSslWJJ2UWl
SXApP71d4jFJX6sc8luRU+BzVVKJRBlZJ0sX0nwgd4WTHq3KvC03mh7fvJxEvqVs
cC/v9/UtNU4YADm6TrdHIjxla4lcSeFIcBWO4gRz1Hvsr28Bew9V6sD/n51+bKv4
+iwziAYVuDlCklcYe5iclsJMbRNtYxHUJqprKSTOpBubQp6E37aOi5NRVU1Zb3rM
ybWeE/15WCPQvbM2pRW6Lylvij4JSnXmvUTXwpOIZYbnYrxYGXjnmdx+zIDyFzOX
8usygNFHc6838zbTX9au0BnwUDwob1snXrExbG/NO2ioGh06PZxrRus7DEj9pZhk
X4TgIqCQ+Z4y+bmUc+XVParEWx+mEr3XdV66dFjjCytwi0e91CmzlMjKNHtYQl6H
z0v7vAGGXJxtt+fzC5NHKkUqCRcJGM37pN0DG0nOrZfqVlYCTw70L7kwvYxjy58u
a1Rfl/V6Of0l6UbhVAH3yCXidcz9XFQjEucQyeuZx1zYnCG7U/y+jNhUMcickxr4
TskIVesH4dKLb6gwxmIJf85unRm83ciDk2MtOEg0JqxDZZmysz1PMSkQZUxPuTdB
viRMtWGaWBqHxnIL+0vGnBpAi4nMi1/GdwGmXjJkKwgZ0z4mWmdDfkdkdC5xZNBR
XiYhIkjUEv06KIe4kjtEoTBs457e2uIes+ZM84FCDcty6fd2pU07FZQHAuTwWxMK
4vbzgN+q3t/d25em5mYkayk+XgiJ5kRx+CEDdiy4z18ajFPtPQRtzLQXGXU8Akcd
vwebd1vCjlYkeCLzUN7K+2IFkQzKVnogq2BgKccAt7ju1dAJCwXYN9c3YGmWyf1k
u8gvMJU7XBr3LtqUrAWbOBiyGGnisNgr57TMW/9SJW8tSNb0UR5Vp7W+BAjqdrVE
0nSCJW9FyoXxfS1K0sATCKc14FrG+CKatKi+46S1fc6xkCQOpDb2Cxej3CwuYG2N
9mCWLDaP5UcJfWFrR6zmF5+lcMN2oyUH91n0JV3N76M/Wa3Gf1Cx3wR8tamjH00x
V+0yTo7vTqtEsA3LmaC+p4DT2DQ0ycOJIbEE3V71E8qibEUiaeJ56kIgvZj1U3Jd
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cln3iAy8w9YhD+bdqA6PciXvyMdMu/sS6lxI7aP8ejIFhTO3d+UNl1CJ3FCG+0XT
D8Uvrjm1UNH4r/kseHbOGJ/gUkpxy2ugompmunJFAmzRmJJTrSago+rRoMvvGjZh
Miio/HhMrU2lgzwsdQMMFnlcRWq2MRDA2/av8BQ+lEU/Lp0G6C/Tv0cK0/wVsrc9
RI7dbTXVV98qYU7YhPW+w4kax8ol04iI49GUVhxsG3kvpgjwKwObd28e7R4BkIcH
fqdrC1RIBBePcqGomidWrXyCYBkA1bMq9WrzFtzfgKt8I3YZXfKqVzQamn1fEnCP
v2xtan1TbYhYrZuELuXmXbFZpYlKfG5GzG3v9TLIVPMa6Sg6mIUR+iqHus5sxqyf
`protect END_PROTECTED

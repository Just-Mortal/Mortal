`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hw+rx7lDmjpwc5bT204cDxOPd0/eT4qlly6alwHEHvYqfM2btkmfQoOmpp8K3XDt
swf5Xrc2yKW12e0LmpZRn6H92joSgAPa+dhe+u2wK2S8rbuqBAr9OfU2VusNj4Jv
cIaUjFl4MsyEPCbjF4jR0cY/rSZex5jqHVhN/4hoYNEvAlIphYqCmivN/dJBsvQu
ycEWZTysgluEh4Roi14HKOEIL2bzOn9x4g4MYWR5+mlBcrlbW5OVBD1WIdFUBk2Z
Ja5L5xGYxzarmJeTXRvq0r7i4Q3VLBT3zGus7k8FaKxhfKo5Q6jRfvGj1vlQG0kU
D8u6NUdm+k1cwmJ4qAci8FKcBSCy63s1AtO4JUt3i7EN84E0QBTUB+3Q1HV5Z5uY
DnmuDXsayVA+LIkezr8IjSI2u3cvzjESgeatczI0Q43uLev9OfaMzFMjOwXImbSr
yEy7lAYaxb3xPmvhJ7klLHTHNmjwMLv9bkXrhSELcFa1Go1zZlQSOrJyuwHElToe
Liy/uMQkxLNaBx9BOPWUcIBAVwzhBZAV3u76yICN4o4zHoSfun6VTNtRs46Q7JlB
wpe5eFYelu9OV3Obu5M/UBc65QqwKPUXAA0kgg+TMDd6HonhTN4AwD/Sdc48oQnX
lwLkJ+ngeNcNRKlPhAebjVtDPb9hWW2Rag1/yOVtj89xwSbAX7e511bF5/WQGHRG
qNeIgA1MUVOrvIszqLp7OADy+S5y0llYeI2oiZt8pM7AJ+NhIx0ZXltZB/WMDU8q
Hf0oZUOPKO6z8R0qBv/GP46vkgr3yseKntw0GLFX2qYjlGcXtR7mXp7X+XiUE3Rt
BHD1UdP9CciyV/vxjTGgmvuAsBjyso043CwIDl7XaJzCp/FId/4URXrpgWaEHwWY
/o0Ey+y5yJoltK+7/W0K9LVDNRPtIGu+46TWmGCQymPpN4yriov/d6U8FMiBVNTl
EDM2xw5KPqC75oqBaxcoM1uH5Z7o6aRoU7ylyRdHHPh1heCO24F3RPTCOtEZ4djQ
uH4WsIall0GvEzE+9hzVxx4Wxwl/M30eq8o3EBzsUd8oglUuZWGLB5whcXzF1jUv
Hz+npswjuSpZYxdendphnrSSat7kjZHFPY3AsOTaTCd4H/HXzr2o7viJ3AsLcYE1
566NpIG8wiIfpSQCj7T4MTTnIOgAqwXYvtff95mB/aUjP4NZZt9qGe8G5IhcN0H8
h1jW/4eoPrEuFLAU1ZYOnmlLjbI6V4MNklLVlAHQJWZzoraEYdq92mjdHLtDYRd5
Ezc0qSpjqwa4gWQufoCpr8VYggee+RRkoH2PNPnKdtEcEEuX35FlmRYxRvaB5Ur7
UiVQHhCV5DQTUrkTosLy6dgDJduMEmonOErVHyc/ht+sXGgAE5K4Zj62v8bpTIrV
AVke3M2yL5/xl8bFpT1+VRyUdoGrZuble2ncDonwuHwwhWI1yA84G/Gk3mu77Tpl
iIFNYFsdG7vdWPxklBQg8YFyBh+zJKzy+l6yrlBYWVC4GJBOhZh5Ko7W8eJLnrcg
B+pHVF5Ww9ZMZgmLjQrPBg4rqJ5DpmTvHRdglwvRkMUp6OT1d3atxY7Yf7p4TGoD
cBlTnLEySrfQeiWN5TRyiLb12Mq1p8D9RPByjhit7hbpiOYmdKODCrxR7LSY8D/t
SsktMcRgL00BLg/ygE8soRm4uqs/R6LsA/jrD+zIIFIyOdOowmZL3AZP7moi1vbG
9iA5DaVg9ynIVvaAaM8a9BVV8Lzz+Ckipp2s2yUtNZ7EdDPGbvIVvlRNmC7D2BVF
qF2NeMXMwujJAIt58mx6Q8gG2rnuRfrw7DciZKVXwi9hxQhtn8/2w+M3RrrEb/Ym
KOvSLgX0kY4llUu/nUSQ4H/6QU59fCV8hzYHZOgP8cLAd8oqx2471EKaIgjQ7dDU
pNW6lUPPf1wjmqKUSbo11tzvx5KWtEEyq/x5fWts2EmBU0fPOXefLWxY467Cr390
HPPxWJ6VKBk2YME7n3U2v507kXap3p6BoIT6hCTU22H5Lt2Y4Av7Yi9iz/vUhGx3
45EPI3zW1hxPp45HEmcQiIbZuXi+RHOjrF6aV46HlZG7uHb37PZynSIKvvrYRuSb
bhEclAmAofRk5j72UvLOg4QKt/akpq/C7I5u1wXg+bifn8lIo8eAtayNq01XerXj
C4cJRMEudaCFQ3LpncCE6PWpEiZQUJEovizvZmJuUMmdL/zF2qjksV1h5rgarstT
l9qIihWyVLpkrerW/EgRzPk+ZvHS7HjRGJBqnndZIMbpjHz34LEaUi2faCNblWss
5891OxFr9qF3c1aHlNgPqRxjbwYKg9eraOwGdh7WKY3EJN1osEv6dT80cobRBKU/
befeXAdQF1qTfQrqyFB1U2mIuokwhC+dMDsWxEigHSqx6bLkL8TbbotIMwxCwBus
P146ysROw35NfOXLbUCSGj3hEcK3HGpjHUkoTE37NYcn3WG72EqmRrWLpx0l+uw9
bTgm6j1RGlpD//bdFNtRVcNvFwCKOjJaGHu4+MrPr1z/Ej6B+j63cpzE2crn+vZU
vmAzDmr23l4h7Lhx+pSM6MXdg7lUO6tKuzKmFnk3+BFhhE0eJF8H7fiZf1+lLddg
pNXiI3uWDoiwzad4GjqMQ1mHRzxlgah9ICRfm6z7eq9CGu0KE1XLkcbdEw02M0qY
ButG9k6ebUTfXwr154U7cdGCHTeyjKZltuA45AvZDfKoX8vhR86Yg474Zs1IzIMO
WRQCpcy25pJiwyDi5NnKg2ahpLaPXWl9bw9btgagliMslrzU6OQXir/7czD+DPDK
Ps20ownXlNZbhgHP1FYERksbqKuzUR6D5zNVkQZkSshR65cfhkP45Z47oPmeoLum
bb6Dv2nOnkJcR3k9R7+IGMb7OfUTSy+xtVFjFLM923gg7zagVTgqfDAg8HToMKyp
SzxMwNc9NrSbvHy+giGeY6jPycLqQTgKIxTMTN0mYsSsnf3ANn3EafQtrI3xhcfI
zmjaPTPQnQOfk75IvxOthmmZgQsxlR1ebGJ52fih8Rxpx7TQZ6K0GgDTVYzVllpW
eeH7gjIinJimnwN1NE2Lg+UOKNvrNy+OWgh3zNHH6FN2g9xHrTE4+HdKvC1oqT42
8B/LIrsjtu9AHnDsPDoiYdgVPhljp7VWejU2w5Rx2ulUp/UKX9s8bzxwc6rSe3La
MVqy9mEsvTM2jAcjUov2aL7vDkxu6D2biw0mZcu0IzPzS0/L3A2jDhGQdPSUbwwV
7wIW6roe9CCj4dcKyumRnmc0SItdKqSXBREZFb5pFAI=
`protect END_PROTECTED

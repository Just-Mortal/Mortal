`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yxmkjG+aOJruZDIoLPc3b62wbBL2QcZOhBrFEHcg/eCCAvXnb88KSbpP2+0vgu+C
1ACduLbjtUmIF4Zo1zT2QXKzUvbW7kB1A3bqV5s1foilz0SmbBqKN3ZOkEplua3n
tL45BpYBs8tMO3tXPHDfOTg6PYWAQp8yPL7Cgt1x9d4uvPIEXT+htgCD6wdN/gLO
nEx9cZkhPSi1J5dYtzyTZNM9yLdPq/7ArZQJDiwneA7OLjVcx4MwLfE7i7JaCdNg
5zUVWL7ohxEbUpky9y+TEp/KJIA2jYt8hQOMY+9MP/BbsR2v2NPEQhBBZ1XJLihM
Im45o+Lu6c527hKT3nqb7+PbeRkntoE7gl0YkWdE+v/0zw0SKx53fU5HrtsGD6qB
SF7/zy2A7O+w6VuRBn9H3CAw/PNbBe59HDDcE8c3Ko0fVivlbL1Y2MkfscHpPP5l
Xae11pxDd85UNSpaezezWxbcUxQMQoBuvXmbzgn8D2fzYllzEo81MzV2NzQSn58U
KYIXJZf/R66gnJYqhgpfzvOdPOqtsUbRIRfAqT9LO9LJYN225EvQQXvLG4jVZ/CQ
KbH/g6cMArlDH4Tp2bo7bierDwE6OoLKfoCvsMwTq/zkPZalpP38o3fbWmFhfHBa
NZAPyMzB7VKpydA/EMfqxAE9EDYE8W727Tc7jF9WPU9kHv+ctVDTnJjeoYJhphUg
f8zsLM+xGgyKzNdWgCq/Lt29TTtO6MGzkg6R8xBXFt61Rhvbetq0OXK2qf75ELNf
nChKV7+DtcKu52pMzf/8YmXgyhgSacE9Kg1AabxRZAJCGoqGugTz+O6g2UwKQqk4
FVY/5P/283vfc3RaRrWdeaAXlFUGYIO2NX8OfxOL77KKYC0FxkzRcs9RM9BV/bTs
xjm4kiIDyHmWSCM1ChXvEn1wd2DW99cfqfguICdz3f8=
`protect END_PROTECTED

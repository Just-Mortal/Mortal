`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1ugaJzYiD7B5Af7joGNHHPLkFxdO/F9lgHs0HGJk0V3UdoOJMNxPARlo8+XEYzU
yPQ9ZsU+Il/nHN8wf2gymGwvCYmoHGBmmaju37clytLDNCIdA7cSXPgjs2E3zI1a
MwLzPbz9yO71si1EdDqdb/WLPL6WBejchb97EHvMuUtZby6baujG24bp0kNpwhLr
QNN6DVzCI7CdrhSIUcU5v0hh+xivfl7WGBRq8kJWz93pOsxg6BuoFajvpbBr6MoV
n4PIuR96N9PjDYqH9JfSb5NMLQREYlcMgLa0EQFRmhzeUj0HiAXCe61exPeT3+Gy
/cueOoYOo/8NgfUm1E1XwscRKidbNca0TsrMrY24F211AlNnLdZgJQq9yR7rsDOQ
/cGXim729OFrWvzW75JUG8WHnM8ksZ0mFAP7lxd+ViPReWSqOvvRG4tIhS66cFHm
TKQy483AXAq9sOVHPqVUIp5WgHU2BE3SQwgO+zKQ+72kAngXByjCE1wHdxdwucwb
JNfnFo0mFrXjb3illReq248a3aV4KLsgF3qmxsPBdefhkf/bC2cWvfMtMMsMRnGE
0f8gNsj+lkMQjKcgMaLOiosnhTYyIH+/hT3qHlY3ZROEpCqhVfB+8TT3C6nLYh/S
tWgBO/JF1yHEpvzN/AfOuMzN4lEZTlPSBIssH9IeRHBkebvSoVI9YRo9uohaq8Ii
kiqMRvfZG5foHDh6ioSRcU1XwS62KR5WN5JbjWaXW4NTbOBZ2kiWZpechoepvN3Y
yU8LGWIt/wXyojuGHWreGR2QRm8Uy5UOtg7sQpGafuInciMrEXtQXizZ2S4GjC+l
cqazA+RGKPOvm99aOOU0xK81M36LvjjbYngmTTDaDrXnst/6fvk4xuxk1suC4IzH
8Pep860xkgloBVGfKCHdPo8XtgyrWzZjI+nkH3ehPXgsuePdyOZiKz8NwrH/fR6D
PyyKQdnctUH5I09cEklR4E0T0zmjAluQoQ36/Q4tTm8/+Qol0gW+eJ3CWWq5rlXn
NuVVIs1ylWhbnzBc/pO83B0+JTX1pNk/RBzmgE72RW8mqwwg67jxrSr9n5RVUiid
7mH8qZOOnkKGSSuKPOf33yhynYucPHMss8UpmEWdi46G6gsH1syAtI8KI3G9+nzj
Yz2PJNYKLSlD8FaoKvZ9fx9EpJo5vuqIAe1uPh8gqZWFgEEOOrZUXnwAaFLFpgnE
p0Z+WdSPxSNcMvr4piopyihZNk0L3nrcQZ4mIYBSECDfylz5nXryyRuBXav/dUe7
cOONV3bIwSVQR9N9esd0zRRvuXIn5ks5xRtVHbIJQTvIjxwnxRGW2uf3hEIx6i+z
bUrgbjVK9ZSs1/v2Af+pYS78JtUyWIdqVbOMZ0T5f5ox9U0Fn+nUDXnci1norpWW
RipNGF3PqsdbG1AYgNDP2MNCSViFGsv8NLwrVEBSw0QbxhSkF4Tv1aP03ujaXYvo
ZCmE3qFMiyZr71cRUiutAGzbIhbIyndZ0RMjzKvT48Kvbw7TFEpV700C5YX5UZKI
2h/UoWQ2ZfybZqnCh9A2tQJNhhZvAlzuOJ5uLQk/iHgGvIuKWUnuWOCxBoAo8jaJ
xiKuAzyYscN/qZDhGEZkekBkk+R19WeeBjP79oEe8C0hf0Yr4Lc2kg4oKcN5xQUS
Fpxn2z5UcxmriFz3hw8jOb4nXdXROVvq4kx+GU16z95PEu2OZMNRQtrtGg9Kzkfi
ZAjFF9177TecyXiz5TZyKz9fPljciKnX2A/pCUaoOsHdzpv1vyggSN9GPqOCzPIe
V8PWeAdQiFV3FzYjVi3bWYDEEQA5Z4WgnPlhPl5035DqSUBpT2TAxBjDe+jMuo/o
Y8OU5FdKXxF1jr29wWe2X50/fI3HQpZO7qiVtgwId1zUhd/GBzq1ohx3eo4TCreE
p4XBlqA4941JYeydPr7HFWpCRS/t6QiSGpAjGr7PpWb/xqSnFv8XrII0vGCw+/6C
AsDvyjauWHPeoRUrHjsHDdjuJXfJqdif5pfZnN7liwzsr2QddLA1vwfZ2hNvq2pl
tFjLU2jPY26YYqn7YpItz3K/X6jMfC/aJUhIYZBb3p6U/QAWJ2RDQu05qXyuYaHE
RnozhpALnXqUNcYOzop5GkpN/OZ9/LKeGLIlMu5/V2C7IPihTQPi3nRpuMWYQb/V
fH+u9YT51aZGrT077ehSBrgS7dDGssZUYnZqm2OUh41czkAW+AkTpJzxs9TI9HWR
xKRmNgyAUMUQCJQiqMjwW2IRwqFXJihfzqigNrA8hdbMzVfe7WK/ws8fWHiu9MJl
xQQSeFI91jqdCqOw5TsuOEoTYAWaBlmkIWJJJEjVSKVuEGYxKL2sSTJ+DSFa/x7E
rQ+y/sv/NGnnUz7PhXfljDBADIqQyHlzNYGqh5V9M9c34ofP3HUHeCJFb0ljlwVo
bX6bXLd5zkUf3/ZKiaqIbIz8bzqdLdBD49i2gyc7upLWRa2ogBxplo52BftVP0/Q
gDTgobt7elu6WnV8mo9dAXbRYZCZwmzPxjDzPD9l9wDyhh5MIINK170FFBwHdIs0
PRbovo/szVrZ3gHpQI/+nKHL1Y7gWqL0awF6GGgLllZOJv1IIbxeSiqo5cc24gJJ
WLk8qlCtLnD2QRSDeefp1AuCPHrGvPnxCHc4sU2vjgMpeqRHnmGz7M5lVDpccYY4
j1yZ0RH9iFHaovRFkCuVX9Y1F9BVBcxbZrZZsZfY6hGNrSa8UYfi56lQSeweHJ7w
TmU3bU/wrIbx0k1d9uMcx85aGwNpZa86vaJ3aIzKPW+Wl9CnlYs+/FfHYNk9PVQb
Bsqj76nEP02GvQBV//pU3zGYloz4xmpMz60+sKOGBzthvy45JWmVfpLsKjyT9tVc
3cdx8fDnn7Z+faOz1ESHKplLWvRXqUGq92w+k29E2XIn6oDkdPf1LEtnfkl/5dy0
w8oxbM9Dlsfp0Pt489h15smbxGPT8tgPTvWXBDwZzo7r+GvrbwhFe6BZa+CQ7az3
0ijyEubh47Z2TkAF4wzClqLXNSZVi63c/60XYMWXLN/xIO1vvUJPc355BK+QSCiZ
2ald1IC9YNhstXaxRnCNuP81Y/mN1hBaFiAGiqyEyiTw6Z2UIe+S+ZmiISharHCJ
GwxeKBXWpSMLZqTnbrWOxc1C22KK+gG2U9O1pyiGTb6C6ibVOQlOOJIC0jpA/mt9
QlVjqTWpVkFnYB1eOyVpkObEqEwe9Wxt+ZzAaim59xl2X7K6LuM14IwYKCnZG/JY
nS99sh8kw+xqZjsZ5DfLf2b4cMGEsTxXrjoWZ+YiSN/xSS8rR4X6eb3US68ObZYw
t7Y2lD9bWYbeYS/WO3I+X59F5F92uEFg3FIqoFijmMXb/QRzYkNKREuKWqvSRkax
9kHf5nYQF1M3WzWSuVU6llXhDl360/ST7bKrOnyZ6/n+fw2B7jvDuBP+uV6+ZqK/
6gJm8EMHU2Y7eWR/anvia2/RP/iLDj4BhnXYOiwAtyoDmbD1LEv2YELD3yasqIcD
kJSnFyfgEzI5BOjsR1HaY/nZa5SR21tD7DhDTfhJt457l1f8ae3thsNDXHr6MsvE
+d4SBWy2q7g1DfysbZ3m5VgiNUFX9fKeZBZ5BRmqFOY8f6DsO+x7oLWXMN7gz4dE
WnuQKSqq8iQUdIMjoAs/Y9MWYguwJL3vX7bLSBrFMrKGKU4/qTxpS/gWMLWmev44
0N/utcCbwaIaAQOcDv7UIVO5UAJzKRQVOYkNLW4KpzeTrJkzmwYIQNCh61Vwiw2N
Xt69mew7afpTWHL4Dw0V18Zu1k/PeI9qC+hcONYf4NqV9UryaNBlGTHON6C3wYgS
ZXf3RYDz0UAQzvlUhUFfJxkbP623MLRdILx8CkyzhZ+bOJzC1Tfpy8i595qiEfHQ
qs87Tp7Lw/J2jw78cOzyPxUOir32G8CEEctuYeSi+e8iUoSjnBpjWGn38jcZ9RxG
Y1o/qV1MtZsZJW7EZrxuaVcXrNTFoE1e1IK33Td0XykqCLay4Bk4l2RmFIEbaGU7
9yZZug6KgjzU/owIx0AbrpMGsgD/ifMyB5w5gNdil+0L3utG9+c3CCChffKT7q6A
uH1UF8ltEcZEwyfGKZ5K0r5/t08PVab+huaLHlhCahDbGC5BGwVtXvVVbjR73qcA
hJdF9jiVDdNXQLQPuppd4zsCwJF6x1G1RLAtwVrKvbVyDdidXPTwpCnSshKlUaRp
yuW+gxu9ktAcD8UTR7uwPkSU+jEYR+jMg0IVFh9AgRWnrMTfvc78yN5Pf8ybK/Po
PxLR9tyzKu/v8eglp07PvFqm+tfFjQJ/aGCbeYVbTgg0+GQ6RHgnfQgOaOyF1ReC
NhND02l7xnxy/YQM2NgQyyRFJT6GXf2pJjmhWwvSMiKkBjcqa1w9AhF5hGv7CsqP
q6dSwMYziw5S0TOmD1OtXejTqnFqXkL+oFummEIayZHyXKNgsPRvqvr1v3jPwACn
nNVaJInCUzEokEW3S1tfZhZ2IhyBLR1mLtSsQdo9ztEgH0sb1HOpN9w7UxBSgW7A
xja2fJs9OlO+iojNgzvvREt8lsEj3CxKbnWoSLe17xWG+1TRiRJRilFClM1dORRg
xw5kC+p6+86kILWm/oEMSOJ8Tw67bkpKoTTTWEWHxhXfqAG2MdQBy67l5AlM0/qx
LzknFgeqwHD3vO8GsS018Jzc8g61rMkc8q/eX2xDejZySiXFHEaLvTeD0kuj8/p1
X6Z98E4W9t5QLHZn0a9p0OGaTW8COD5DWpj0UQAwNG44Br35zRB41oja4L7cg6eP
zq3OtTwSzeqWztyaoQZF4D7QU/1tNTbJGejJYhFzW95CzrVAPSo7hrvWDJS8Djfp
fOLpRqVkHwPN3KxMvDekboviUOk3oe539Dbap1kFDNp91KYsOFGDtj9S0dJtjzKu
EoAESHPxf77JPaGN3HXNSs0hp+iRmmGgXLBL7Oat1q9iJ03XzUzXGumzRN5VMbAl
KA6LL9BkmnizXSgrDkxUgqtLxbkiNkky5hPg7AY3Opwcryr3ngJkex8HWzojW3kZ
3YuFGDQvWA7NjaviwRgKdC27D9EffV1KadnEZ0QLicjiq3y3nY8B2b24aXPHMNH+
m1ia8C3zoNza/28Gh9VrP96q/hgeZjvLOtRhWay5J+hZrTY2MkqIU6NftehFMLx8
RVYudjyA3HkaxpCN9YpxzMHMJ2judNav5IiuEzBwvMk5zGL1yoT9fKeMP3nDBnVV
fs99kf3wOgkXpT9JZi26P0odMULaj269MfuMiPQDSEMs7DsgXT9WulLFzOhuOIv7
7t0FU8Km0SLtZNNu0SRs0W73bJSHQe1rZb63Biw67FArQiE5BYVafD9qk/T59WDf
QhF+TxxWWBG4CbVEVizHskVwa4k2ey3L1YrsLsAsZ27HXG+kcT9WPm/HN/SHIGhO
YnqxrANZktQn7n4OvUYJxe+HoQczTlrBBharukyHJmdpJ/FvWxPk4jsHDqkrUl1o
nMSv5hcItZZu7HQivdUzD3EY5J6DFb0kLIxaqllZKEfzzTFNJXhreRXBWA+L40Yl
9AEKjlhnbpvR7eUTzl5IrTBSQLfvH+/QytypUQf7oYmi3g0fpR/nGSx98qyGDZOY
OwVa5E9u1PsfAqbCyQl8OMV8hb6hc4u9a8VspHFzeu+SMm8u4qf/X0wt7axR6VHe
DYOMFlQu8csKlYn/HzS4TtiuveiThMngLG61li4bLoqgAKzWap+EKXv3Rr/JVxtX
s0T/tyuYSE2zuC9uUF29VvI+2eIOtflCMjp1mkdDVjzIzRQhbRgi1/7G+OOHPxO/
Y8ScYvjKk+AWyjBjkJROid6/rCcqHo3bop8tR3aHYMYE4LHcPaAHCksgQl83ZgBs
ZuQYXfKv9nYZd63EhrrV7WlC0CnPzK82ltCbOLZRaNLUE6Ke1XMR6XweMP3E7P8P
GXaa+PFdEDl6gGo3EOVj/dHparD2Uugxdoa93zg5ZiAPZrMABCGpvpY48tyOV9ui
CEJj/NPuhpNK/4WHjFvRT44b5yPjaiGx+vLQjgRwLf42iJyJid50gJgDu1BOIqtG
QjLCTSpMh+OmAQtjDZQNpq+4QTiVh0DI64MjUROF1yR55EtonwPrhDBVNq4uJcbD
GtcKarJ5GkToY/ha1lmwIfTPDymuQhlxmZF+NOSlX6tdMDwO2h+Za01w+M3eOPzA
koE+GrWRYaoxEFkNMNBLW81NuVjXFxVfIxuf9hYLTw6zDRBs+HbTDIWyWs3Wx9It
tH6htAD89O8htK6Hmli+g0gITiKXItum13A2ycbUsndsMe+5+5Hn08zCPD6wVR7w
sHc3cNtVnK0G8TJotx/8LWTFWuWKzl6stJSrTBheICo+R6Rjq+LDHpyrj3DjExUQ
Rek8/PViuzp/6Fb3zRFpRe3gpoGxQBVPCS/tDpPLCalXQL/RcrscVY4kw95j5bcS
ZGI2379AKQtrxux6rguXbYQ6nNw2nIM8DTT4s1uoWYoP8FEEmqsADjN8c0LYz0pw
sJBTEn42C+J5NbBHmIurMc6fB7cTsmwGrk4kbKm7+/K2PQ0PoDXJYRhl4MjKiM6r
qALiDPisWRiZumqLUZNdAZ7swnSQIODpzex4jc5+bRw/bHR899NJcORDPp827d2T
fS30rVqN48/JmHIu1Yp10hc/EsnwdZf6Eq/JSQm/V7jdIFA7h8gDYuZN3B3t4rWf
7/brwGx5RqdkYTpHnbPdZDdHhMt3zeI/fQmzbLUDjkdiWky7cGMbuhCsaM4JYSma
TAbT2+bGuKSCRQZdfJXfyecusx7TIhDGBtfgpVZTfJ16q56v4rjftj8OFpuCLPON
y06XN8Ej1mnY4URDPu55ym3+VkjMzjkBhlLe8oNTGi+DjIjrpoyYuNXObF13J4tU
NM09creSSDI8dHLyZB3qqTfZTbETmX66Fu9fu8vpafnxBTo02qHTNUqpTQ2mZUQ2
9db9rhqO0SJuywG+PRsMuFIGjBFLS5CbViRy7gD4CLTAizWsz8Y0K28N2FCnHcds
SfhO/TY2lg5I+VRg0UjWsv4ejTU7tSK9gObJHDN0ApG0K02SFlgIf2WsbvlGMIOW
Fa2e9MMzFuuy5J6+9EcVaeGOnGSoS++n1YsUTBvOQV9GKDOHi8J4HZkpAOvEL+qs
T0uy14N0ojsZhbkGLdniTHfvwI+ZGj490GRHzAE8WVzoyQuS1V8DppqSIpGxgfrP
7fQ/tWYJ/VlQ1FbUJAnFoBykI18H5JWOzRG95l4oqBY=
`protect END_PROTECTED

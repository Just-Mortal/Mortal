`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vvnGgPd4zF7DddQDuL2U/twYfaEz/Hj+1SoHldg3WHj4sYE8e14CCHGwS3vrwDB
UPMK5lJ4tjrTk+csTvwd5ul0jt5Hj+wMxsYX7e21Cw7pxOKva22qmd1+/O5jNuHt
KdE/mk7mabzul/GnMMD2xPyjfxASCv/4NyurjKf3/aGczcu9ZwLqfxrsQnrzjF0q
St1XZTt6Uhadj2IujMPVqwsg34M1xDX0o6KDMwSjjD8WSAKlyU7fiK/JMc4bIE77
CyWv3aJgQ38SVVX052FbiU6RBxi+gsayfylRRIwkHpempIhvMHtjaG+GiJNMBy2S
QNaeoW8GKFz0YjAj2gLWVnmZ+jpLLZSY9AYhqYDHiYP8DviCv/aa8nEH4KI7unQL
vhOtRAF93bDJ1iSFgUEyY5Y1PT0rzpMjhK9Z11AFk4hpbfTOsj7f1uWZkYjnoFL2
leYwD+KhtU5XuhotYQeCdhWScmtAYd8HsGgXu+VWK0cnAq9GOg6wnTC+Dzt2o/zc
gHNQw4p2MTJ+qGIZaXnQ5Q4sKHp68P30F6ISjFRw4HxbaZdXyKgKFsUqlyGHV+Ca
dBwrjIoV65+GE6TiXYtcjOIH9ltJ3xh9SVw1qhyLmdHa9KVBaNQUdpRz8plB8IS0
oS4M8v6eQmfQRUek2Ag/E10/EdkFoeF+0QEECxE+Oy3bjw4Iecv53ltLYKMg6reX
f8N/jJZlRFtRGcpJOvQPGXyHAY8O9MZPZA1u//UvCvNV8EqpO/jK3LeNMF5ssJMx
GFswToTFMDARmLyLbS+T4lMYqnad13FqWIkOAuLtA218krb+bGLaLRsyuiLbTbgM
yluV/4TJcgbT6k8M1AFSBCVdEaBxAFJ9HYpDWM4d8DBDKPgFrEEI4eLa3AVVcJGt
eXsUnsPAvs8M+4KmZF6YDWN9QLevmWbT5wlp+QVsgJqug7U2XzTGp+Yt3SdLlCFB
Bv4leVB0j3QmJs6S7+DMT78Tyrjju3OucGxVVeEtoxOEAkBpjgzYMRbOGzT3yDZv
h4d84BRh28Z9R5aaVfJlW6pzyigBsnyNYvCvu5/96Lo9jlyfkjoNQsGR3yiIxEJE
17lO2Jx7z1tUW+2JR49uNubRBlkxAUk6DrCIyUtwOW+sUJ/kMdMKkg59ZV1zaZB4
GKQ3e963Is2wDT1nJZ5FfOf4TsLQhICbDqr+ryr3fchLCTGM1CJlNnICqMgQ0VwU
fqBcpBe3dAzMUJkJhy1xcJUbOANWbKugO8rDFPgRWPh4I6zeFvHV5Ofx8WPJvGQ2
PSsNL0oDyqPSON1LXZGV1P7AKiqri5JjgzpCF4chRBx6CwrDmq/DMmqeLleFzhNU
VvV7CeHuUWepIFvrOzGHyomMEZiFEE/BJ95VNs7MboRmtnUsuZSl9CDek5m5mIcB
cZG3uR2cIFaMjC1m5j1j8Hz9fqCSRCsxWdlOMZlJZs25b8oV0xTrOg//1G6kyrKF
wTSWMblUflOb5Z0BH/DVXwfZMdJbcICnuGgl3b/0P5RQBE7MB+teQ44ysn8tLqjm
oyr13e9cIUDUUaMqFdSdnQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVtO4Xn7uRGchxDNfqJdWfst+BZK0l4nyET8b1uzUCXD07CkZHUyVZmcObqwRMap
Goa326Qzf1RFBtWJAy6g4rndtDNvydFSukuQ9lJ3mKkpFXf5n7SzdhVqdTGPPmto
gqb/AmgKvOMzNGtt6O1PSKnNhkWA1/tAt4TtsFc+lDf/Hnna8spEzI+nXUA8uM6C
5hiyW73dmPxOXDpvy/wj0zFJwf3QrR2Avv6LW/kaP6QskvonNloFG0KBM99W3wry
3GBm34m9/uCrhYPPvPjp0YLv0Sojj/q2pIpEzfMHOelyrR280v/JBhfdJakcCjLh
5e89btLZ8X1UbaErv1IvP34rui25zkwol21g2u8HWGqdzbFuBS0fZZWchX7z2dFS
cxE/xPMJfTfOQMKffsM+vYE3WinqLXaUDIMfeYFrPQmXR3DdvagNUanW+gXQxiKL
yWOisZdBMmOVW9FXoYzEa4omB+QOZzXmO0OdrFIOiy/4HKGZ2RE8KXWOjCzMy5iV
mHQQWBWk41JcddJh61ys+VlfeQ61+cHjCFS+v3hXFU5TYJvhn+Oepq3FIzwJ1K29
NDqcFvvSsB6bmez2VIykM3mOK6EW7q2ojAtJG/vOzeJNIVGWBUdIEfM4GiGjvFbc
/lWi4lW9/ctfjvUw6w700v9fftx9pOpPcSnjjKOC/jcPKkO4zyBzOeWF46KyhLQs
p9voOgwNS6wPIpQAihCRYAXEgXSfcswakqB5gTVRfN6OYYa3tsZNXLK9OczyLt04
qOQZCwXUfAYeHPqkr04RAMsqGGW4mU8S2Prkz+KiU30lG8QPbRi8jxkj4bbQIk9J
NPSvG3OTWL9U9ueCHs203wB96T28gzEZFtJ6kCAs62/EZVA1WDSQQ0EZMNm4ZHTH
2uHvdCnZRstaJ9d9B8852WcHPlVbGYllnrpLceXxaoBHP73aF5WUncSghIkcVfQO
eNVz7M61q0JsUZ/p8ezqwMNkIw32ep9UFn6AJwUXd08vtpYu6d9knbH0lGSTJ8rb
Tjv5ftosGVGeT1lqBOr8n0mVJtpkf7X4wKN9Ci8bmE94kHXuxWhQ6RIi/Az4Yyj9
92of95G2h3j1ZLbDgPVeC1Fw7YhNS8fGfuYH+KTyebLwk9J0P0k+EtxbUN31BbuR
fOc3pL4lLhuaVTZo7u+Wtg3pq+KpfvyYa821mAhcPv/cOfqGO3F4MzWYLP01EH59
JHlaKXEk8eDWvu6zfA0Ej0HKW9WfnGYKx7z5yjW8Ub7sCwPUdkEG0Hgw71CVwVW7
hCsPxV4ZFlPjb5F+L6CSasI44Okszwb5ca7rK3W6hpAL5mN6lZYuQfDN6uZho18z
78OZpVmc5E8KiXAYgyVO5+LR4zvMJ2EynYbU9uMqL/UlxAZptq9pc56y1NrIy80B
67j5L8nOjAeTE3kfFPrDKCZYo5mSyzWDh9huWd91fP8bBrcgKA2W4MamS3nNcUCB
FtcFM6G0XLxMZSAwkagX9hvRVYsJrIiNv57B8ZK4k3rTMms39tAatNXNjEaKSj2y
NcHwuC1BATidmxTc1mx5Exllvb0KYY6qW86wnjTMr+vih/Y+uOlJ0bB8UBis+9Y8
q1TeP2uaY8uv2rVImYM+KsCUdQgYq3wy9I2v/0n3vDB6tYMvG99ZoBzslGpXS8q8
`protect END_PROTECTED

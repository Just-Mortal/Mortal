`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jk3eyf6BFznaKOLt+fVMTg43mA9iYlDiUHQ4QaCVxPNPiUQ8unVWbq8/fQHPZ4Bg
fE4FgtnlhIfd2GwrJ73CVEc0agImkMGQPJJP/fwGd9qLfObn3uTCHKjTFz2pWTlJ
gMnQDd/x4vcGcndCHYWiLGa15r/eKN5ODrc6faT779FUej4hkalSDC/5Us+kyI3m
rY/+c6cexZtU7dFhHb51Y0KwBXX8OXLxjbRTt/AbH2nNAP6/n7mJHPZZDcEVVrb9
FvhCZyy18fkN5jbmf0mjGFwNNKUSzzUJZoG347QcXkq2BTEFfCY8SCET4zAWMVEJ
ApnMmnbieUPTWNqBvnzzZGCMEBM10KlE8dsulYQho934L5XwJ19jlsHwF6zzwqSl
g1zVcGr5VLsK3yxnfBO2SbMejupGpHO5UcOUBteCihseSDRjsgbRC/aZdhUVI60N
t6J9latDwiyJPyAvHhtEvMduF+Z3pcd0lWIxXWfZnEe8WIOoQRBOGPmnLkcfHOB0
4k8zEcMq5a7SKa3ORr328U7XsXgElTyUw0/7REqcp20M5pMyDIK1TzuSsRI4YhH4
LxuuuqFeMrtLoEZaJTaODUja3V0l33jjoxlm5QhLl9n/aGnjZCNgadihXQRaSoV7
qpMP2NKSJy/jKR7CfEsjJ7I79a4p1I275RzQg5v06uK2nOLW5B+k1m0wiI6xaa7R
mnMj07uvxQPjMkyWvr41A4qWq5iJEviqIN9U+O/gJiKD3dBagvsoIljlSS9I7wCV
VaePVT7nL37XjEWy1ihpsKZrvmU92AFwnBxxWrNc3GiAjuZ6BDQohO6MGMSRclfl
aUS8SR4dgwIvK8+BqzbE/LJBNDQFEap+btIn5YzAdIryMYUL1MIdS8bQOgRX6r/2
t1XvTtatghPAOgkVGAuyjc9o4pixkLNDzL29YH7BfDkcI4AIIu75LwWLzYS9s07h
WtJJZSPr1eZCTJFch06JFcc7JWv5K6cn0r/KeiPXpsMLjY/X7sWQMCe4yUofwgkM
LcwfBuIX7nLPhcHY50hTHQTraAcgVcxc9cbvQUTYw1ifkugJ9G+KNbtfbS+VIm+2
+vmgfJ/vDdcTDxWEoOAyJ/8r7gZ413+HDg87GAhKgYub04qs+M0cMp10tqjV+GC5
oCwBD+NTQJtbvxduzEiKHgzeoFamin5vwgmt0KKPUxDU/YxEZ6DgYLk/6H3vgLZo
nHbGPtVONdnXG5fmSSObE+uQJwq19k1Z3rky0q1GSTGFbOmm3r7aLjnJdUyXgQbq
gfq5X4uB1340xfAOJ8FIspZRCfUKcZ9SeSs1AyMx0HdlbXZqwn8KlYFmCGIeWjqS
WIYdOOigPn0sSjL7tGuLmhOPCw1lE44rEY/V5M6RsqU5lBCAUKJVpF6IGb/H6MdA
SrLOFT44wg0chSsBN+43gEjDTi/0oRRsUiWFiCQkcjRYrxkfAfVl3U0uVfF5vuGp
NIuqsOHjEvwpR5mFGZIVtyf+xAHoB3Q+AN91lSZ0aHqcCsSrPHv6W+IftZLT0tzL
TrE//CENjF6tmrxj5g9fNyYef+hxT8WXtROt4+FLdgH/iSQRXxm55ci0VVV16VrS
QuQ/AKZoYxnF0iBUUbpYal7I3KoamIE8DoJ2tpJEL/LxpXC7hMwA7/gP6O4W9PVw
BE0+bQHyOQYacKdrB3dlaVhbTIEpMtx4Bs1cvf257/mPglSmvX+3VDhQkFSvLt3f
eMGnJt93Gu+zfzMiZcnfVi8u8+VDPe2z+5hCFszGfmZYTXV2aNq9yWfXaJD8dTA7
wpxOqD62YOdoBiCIsJj9H3m0uyl/VJagWEoA+JHdr/VD9TIaUZ3VawaMH8pSlRUP
3JHwZsInk8yMwgrq1MnTKUW49YWDsgsxrdQq2r/BZkazf3Z6dwXKm5HhmZwaFPjj
YbbmtHmnFXcRMaNNIQ3YOttGFnLqvm0ZGartumW/r8MrfFB1tykjMpRNVVHKZLdQ
WpuUmX5w0JlX1RQHr1FXjRXiADGQG9oaFQd2YPsFyPdabtiZkM9HM9fn9JV1yh09
Y2YKDH4j5siyYMHi2v5zCXBJUZBIZfNsTRf+ffLc40KA11lxETGkCoCHjSn2tWlE
Ofh9CjQpzRkHHBjbQL6txWTHQypxbKt8ufibVJix3N7+mtnFyyoqBHixZYjSWea1
ZSdkhhYI/DR95K0EpZCohHPWDAAhx+2/Bf97nVKSsLEFTT48bVpwjJ7jGln2vnqN
AgDiyH9FC99/M9nn4U1pzSJsaANgoSkncnEhoY55XYFYPzFp7gXvvxhowHHQ3ItE
qyjqrat7Etg9VzeGYrBwZVMA+1E5rHg6WQh0UYRBtvQa3GOBo0wLaRHCYZoZ5Rd2
17zFIPAWapGTdb6ofAZNcLa3/d2lpnpwHyrDnKmSbcwByxMHzzPiZyCQjtlKVlzL
tF7tNG3fg24nlMms4bQe6uxmugZaIcbfZxA4yw/FIKMV0U7x3+6LrRw9Rm6ryZpP
L4kHURDK5Lx45oRKv8Yyl0H34l7rTbPW5hMOO/+ClQDdlHbA2/tbwYEMgS/axrbV
cF7JnS3hZ1BCuiBfpmkAqxuj0zatgobBlgV6XapkKvEvIwpLydeOLjSfRIYLVosm
OpGsKYC5CwrgaMtuAD1JavuJwjtutmmTo12p8avaA85tsFyOTKcPMTs5tvaxssiu
YZM6Y84Q4Y9KcJc1tBT5TIjEmOy+gXE8CMu8QZCTLniHxyt+r6X18GiKI5tEvIAO
wQavNv3EoWTd/vR6+oCPWYq4VI9VjLEnV0PtuqChjFB9XeL6ZrZay5PENx4pC+0A
McDMoHmQwyCt8u0mRQWl6CIkEKaFnRo/anGJobzd8x6NBIFCtkLxdb+MUOFhJOSm
MqlYng/qfh3ieQFoqZK0AYFfM6RBWiG1fL2L1lGvexoZsLgPdYxUbLJ5MLS2Bc7F
16fXAkcyAFYrz0/Qagk1tESslydb8+Kj3VySTUZM3McS3t+HFbakVR5JKjrd4J+M
6RHUgmijsCHmu1aSnI6orsGVADzXG+JIrORYzwSd9Zm8s0aEu24AVTInCFC/U59/
JFNs4rnrdkkGSB3iyRlzkRlMryqueWFGmS+bZetbocSRPhdJ1SOHS6UPQ99vhuj+
W/TCerDH3te0U6CiFotePGd7KtjzDX1srtFmzHpxzprRi2BueIeMQ3Rxs0Dfp2jA
D2cVqZF6QfQTg3CiFKze6CUUh4rSBhCXNfEZw2DkG51ibbVZbpbUwyUHG6EGYlR9
MlWy6WJ7P1jAfXGJQ2yAIGVY6Vj0M7gc4gKj0nqvdyTUUA/y8Pn1XaR9x+tLtm7c
yFwYZVAeIx02/3GfQpIc3mk1nccJvrv3zag/hbL8Le5OLPrK568ymgD9aju/iJcM
BmKhmriVrNvek+aN96qT/63qyD995EbXEHnYHZ33Jd9MlC+WJsc8uzAgZ6pkr0c7
pLnD9MtJQ7pxNcJx3C0FqYpJmWm7jqLFwMfXAPUBxHxQmv1Fs2YDjNa4rS88dXfa
lnzI10QsZYSX0ota2PRouEl6e3iJ+YDK5MDNs37CnuOZ/+vJNhbpjROCiXcSgmQ3
t3Z2ZrIpo+mQRnmkMvEqxtDGioMvFfjinGXIY5EtfaHuceUXPWjyQ5CehTb4G8Jo
iLcxc2BnKcEHwLAJoSL2j2mNO27JOsjz/K7K4BSubn5mNvr4/XfmqhRxjydeIP2c
uS/xmbp5R4H/XIE4ma1AG63JIDSRvRkI/oZOPUGLbUAnMOUaWEYHIgqMfP2V3Pyk
X17/4clauxMXcloignf9/FQqRs8SF2h4+wgECS/xDiiYLOmHhNLwAcWojAS/ff22
XJ74KO9DamdZXAqW3/Br1FNPXpNtq3C4TyNE+blcv9tW6/ACAPSai9aKhsoH2qFo
1UMrzzyINycly0GjJIkJ6+tSuwXWkCNStHVESE/KfwUpeqTYWQCZRQiQyQOsKem0
w9Z82TmKxL5jw6wh5PRc2WDqYYoc79EKuHQMhp0o4iFTay7hrJieYZaDje2m5iAl
NUrwDkiiei4V3tT48rsZ9y5CKRH8xQ50wf3m45nKzzeAA0C5hEenhDalsmVQ/5JP
8Het5QiJWulO1ngdEX1oJeAhj9/j4ijm8xMS5+hPGWwE9k1M01bTNRTz37Jw0SmZ
yH2lkyUz6TwvN+CW1ZO1YOUT8eHf7Y+p4Fg4ODig8bZ6NjudGxkRKXoyh66SnSkS
qQhB74K0gVfdtyARDFM+kP3G7L8xIaXnFSJ+aqhHRTzml9Xo+tkgokodEuc/QzZ9
CS+oKEMtyDGQpvgSq3zTtwP/tw/MjdMuis3A6eUKjCGlk8l4fjIGlQVqJK2c8vps
7mWedkwakF4d5KOTGYXAtRXYjwFvfnngld1GEuTyuSPmfV1qHsIXXxkBg8eIFI5K
o62t4TzrdxDZag8URtndDekCHbdCq3Uvq7gsGifHjniBbUfkXAym6CdZpKDiqedz
voFnriuUmgDRSjxm/x2XIjFiEPpBXL0X9bTZbCfp76wvOZr7BnvGxoB/IDTmZ8rx
+wVteZMmgh991L2SWZcvM9khNVq4uzLsw3WazKEGq9Na3MIkxpZLIsUUT5oD8MoS
yE+8b7xoxdyjN9pf74QBzlD5SggYAWmElWHT1esi8MRVDjSx5Tzs2TQwF62jjQgh
v1+rJU7oIVIwWoA6VVp9MmljmJl8ovKblWwcqd++u77nq4EhW15eDBGQS/3YBWp6
2nSZUlrIRck/a6AG9dsiBWMClTbQhAtNQtxcOGkGZ61ITCqJqy0Bfad4SkQkgzaS
8qJ/PnRVe37pqKTkDrKYxma+gnE2TYpcEhlZXW01qCmC8zbU9Ht9B57XFN49tHEO
maJG/nnRsPfBsGnce2g2FRGY6+e+YPLhwCKNdVNrv3y8QNd9HV6oyHnQRWLzl0x/
Pp4B4oR9CQKmqD87UOhO1WJPtES5FOfCOEWYYyezFufYGHh4y3Kb1BZMDkp9U1hL
B6JplbPnXC2zHQSUKX+ti8rXZjxf0WfB+91zAHWhViMN8OgqMqsL3RDkq8ChVUGd
oU45b6BN4ZFFnJf4b8EjKFZf2cn5+UjtR+csC8P5g6W5s9pisT6vJ96pv2hw1koL
gq8UW+LwQhqw4amlO4eOI0HCvEornpRwr9XFPOk5FSm/xIYQnzvGuLFesxCGrh7N
mMcCWmXc021nCVG3+wjhvDPEPsND42TKtADfEjV7KABpQgB2yH5omwVlAEstcRlA
AzN+HNEF5m8mg0o2VgMMrYUd6DLt9sDJSENUfZ9Hf2EzLUWWjV07U806olSTt9hP
vp9oXl9HbdMa+VjLQAgoW4ABUeiGMp27zcsEB0c6PZ7lDmUtYi2IdA3ocEQCXRMk
N//cQik7R/a3Bi4z2mczDogizTCoISe4KkKbK4IyG2ln570ZnwUd0Y+tIZeNl6r0
fpuFmihYz9ynbh5VVDKHTj2qxv8fAJqdr8lYIj1SIB/w17oPmXNdSVvM9xpnCpc7
a1SYYoEGjFN94QLEbiMUYwaEa8KEAJia7JbYi3CaHmBiirZU9e5sBpXX+jVJMA2A
WknV8HJjpQp+jKQn9GpN8/ICjfalmycA9wGScHoiCcnQF9yc54QDfSD4B8moxFG1
K0xfRQ2o+SkbpdFtOepXnZ1GfE0oHHr1HiQIoK1sK49h6wuw+2SuORBaKDqJYJvx
V+OVhYVpsdviU/BbnFQ1xidNAN8Asigc5P0ORii/GbGwEK52jfN+lZUmURj4DTbT
MJzMb9/0GEiiN61YHpTd46Js7fRhOv3rJkJkS6XgmO102os/STMDn6EGfVBtiamN
pPEmiDPzv6hEqQxCWwKzm6bNBPNL00XmYQqomthlEmAWPuOHUz4zGOihHjwSNVmp
5Xy7jE6yCpZwhpamZjhV1JGy90qGNmpGSsF+i2mv1OuxBj8OyIFAJOAxtTUnonir
8+cSVKXkOrbHlNDLMChefaLsyg3H68oONBJFMCg8Ig6wdnH0pVSBlAi+Alo/lOnM
YvyBCDaXZJCAoAWWBA3V8B9gJEIHNVMbxCjjmCuqjO5BwD6FAGWSW3VBUFVRwmkJ
HrZHHo5sHZGOGzgYTtMTGIhG9VQmWJm143i7fxTU1BmZ56Ov1uEQ9S7PDOHYVnPF
tWKPsw58yjwxaywzR2jgTsJQ9d5+lx2JgKxljP6OZ6cMiicxal8VYNta190iLRCE
dq9b0L6MR+oa8KhM5MIXZuKHqgkn4aUSDJDegsyuuWhdEN4AF0fWgPkJ7Ixds353
96leQfHPPmctVIDQrZIc26gHg3DpHrhjNkorTNZQPGutkYp9beaO21dEcBp2/ukl
5t55aw/BQ+HV9S8P1IwUMg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+W46y3tE/7VlW+euX/tVGKqMctwYIGqgHKbIUR1wZFmRJrFTN2kLj5gmA54Ehxzb
cHMnAU/ybeCQbN7XLzYcAY5oDz+4jubiz1YSTjJTctgQHrmSTZaHVz5db4+InEDu
FrUMYd10dK/IS+hthsdFEZ0P0xuGQAR7zT1jI5HzqXn/3ASBBp+hc23fA+fJX2nO
Gf2zxPQRZXgxZ7S6CyqpDtjWXPMxvgdZxwdFcepr7tMJgBAaE6ePu/ds57FpBM3a
EAmFC3QrAeecMtM1d2yIEM+Rvslhu2d1hitTsJgKCFn/B0BVSKbUkZT1e78xKkFb
uqy0mQunnUpyrDXXM4rqTGrOAj+1eGL1UcxuROdukgcIqdFlsyijVhOUzLFRcuM5
jVE45j0p0UismVRQ42CebQEx71YM+r9sn/RNRAhEg0g4T0BTL0xxyYC9EirX5tj9
2yfpC0NMjWBGWAy/idBCK7HlUfoaQpObgfJZbuux8g9lFGGB0U4IU7/kaVF1tFrO
zUUaZtElZu7TBcO73B0zJ3/3aqd1QP28W8cp26rBkBDGFUGNjRoBEuMWy+5nrsTT
zf1OX55mtEPClaE0e1UCHgUnO97LZ8EWurfsX+Zj6t0NNTdUBOJVTGyTMouaWGuO
rI47Eee6fMQrWXkYsI2TS9tUdLuxNyi3eQZbjro7F8mkhbT5h4ouOFJyaCF9ZJbX
agyI3AWnelUiZXuu95tXowlFpT0aO9R6TdNUWhNzp6H8YL/Hsd1Qnd717gT81pUm
PMLTLvzfD+NEqMGDORJO2ZhJShVnWXF6t1aDX23k6f2ow6VoQurI9ZQNaZSvUjY7
4tgj3xMm8b2/rF4z3X0E/MMoHFlSoI/2HD/tfBrwET9QmtY7wTcUh2vygSpl/NZV
MMAhlnOC8kCOoNAErcc/xcShIaKafGF1ebTxBT1v4/Qv2U7Alp7huWfJU0Nlx+IY
iP8O+v5/FuNgGTMawZOr3SuEzqHVa4cvgPXXoEUTMV2+G6wFnkP16lMTfRXu38vW
ovKZh7xNCYWr+2YSBfYz7MnqxQlT9D7h6SLcSMQ/3eoRKGa9IijuQnXr6qDdTQSD
WxJwbrt80GQfUOCe1NW5yC4VmVKE0Kwi+5dXisCe+HCpm9BLZtJjhEcNNeY3IhZB
A1pT/FkIyHle4Y8BsIe82HgoY4RSz0Pqm5iqVa0VV9MQ583PEbTaDiNrA19Hnjhv
T5nGJs9GzNPg8/92VvQeUWgXiqCjcd2ECvVAfGo4bfCvCotkVVgvYOE0O0uNnr5j
9zaRUMP6HxRVm87w5QUvkTisZMfw2UgqhPZrfuVVE2XZN1z1bUSMEfp2jIpk/ZpG
phRkrpg3sP8T15LSJ7fWO2z1YhPuIPsL9TeJZHsYWplFAFkTXnn43CZIsHdj0YSP
Lu26aR4DeolTw8B8Wl0k8hBiWVy4EEnxK6HbaXZ2w6P8x9mO/1iekcCXy6MQ4qgS
/GnaRANyQ8XuqF81I/G2zy1l7qf+K5DHs6AIBHvGH7rOkdh/96QQQdx+xO2EKhkW
eeGCfihEA7p6tN/VGWZj4QgcIor9chawCdHSwl+B2HbfR+FGaE2sLhty+hVMssT4
7efO3YMEak8CU10t6SHW58+hAZf/HZdova+4qKPBibpIY/s6mVxa+1unb/HIaevm
AZDWiIZ5DnJx/vuu1VGkLt4rGfLhkgwjtPDYIaf2cL08xRaUbn5Y0cxBnH+jazKu
e1j22uc6C/rqbGDcDYfqqGKzjO0/YdG0P7J/uVNSAiGP8+w56Zrz0ZFZWne8kKB8
NA/3R0cGUloD87z+wl6tg0nw/7t/1xY1GnQtxUJtDMV+our+oD2SvOZcy4Ouu9/B
gD7zJKYWhq7ofHEI8E3MygC8KsPsQyDZiJn3dlqqbfGeMSXXrxbqKTuRK2uSAXoD
G1t8sEwQbhwccBUOLiofIXgpOwlfTXPmWKGcwxBm63JIN2pcYop6JYHy5Jw2LGeF
IY29or4LGBUx1ffdHFgSgfgZuzyykYcbRG+tA6Kce9WVRts2BIXTKHlWoAicX5Tc
XTtr8Glkg9MbXYkvuqd9XcQ4pHJvz2IlD8G79AuL7EzJW2gmYuasHjDi8RV9xEHx
fC5CzWrhXUd+ZRP6r1MtTbzb8h1NApAr2WvP9PQEWuLXNfhoFwtZtpoA7mgI5faO
nvnkQTARGPRAaZ6wMiIllQFvkH5WCOlgkedBZA5ZrPow8ZiipjLMx26U5FYTmEjM
dA2Q7pxJczqyjNgw66RAdipr5EUwwT8cnrDdWq5H7Z0L/OWkbXKK6rspi8EhhXl2
BwXXMsS6DHgD5vEYqdlrrmPoqtqWjXhFDgwmBwJrUX1UJz9kwXPusTC1GbNc6A0a
8gGMbBzamyRy2Nf59lymafSim0c+zfmmfUPWiibn0kY5M6vHpMl7W0KgwvCok0dL
OTXjRAO2PVx5VAKCoGmpq+8Xegl/PFbGGuFdhPPbLEMnAR8KgjzDd3Usn3YcA/TQ
aZSxw6FjYm3scMxkBojd+263gcNVJNDDRtpYc8bxzkHSK/IfdMWdWCcGRfnksGjW
6eT+JzgWKoLpFa59nv7KUhCzLgm9Rzfa828xmPzwAARYEMS0j/ibkVaDutfs2h3p
2WiSZFBF715Ch36hv4a90heAIiDGXKqomPsCXFmBTiTYdQT/aD4z6XvT4jpqeCfr
46MRNWlb45W3kkogsa29h2occBbCygkMHAZhdyyYW3Qs/Kz16aftAdrxWMwTHs51
zWLj7sV/0bRaeK3JTSvFz8JKnMx9r+V+6UNvoQuVqU52JbWUkJyDyy1ryoGLe6p5
jy1ozX5YudDUFkgyKAe/bdl3PH90rPx+Cj4c8lnCSjxCR3hi+IEeAUYnaSQci34U
dHtZ4cH+Y/yodlgOSFmEkQxSWMsw1YR3lMfjRz9zcpSM3O8s0QS18KQk0atG6OTZ
HLpt0sQSIpEStaIbk7BkJGCEU92YbP04zcw4UfmWc7NGaQjOp2e/rrBi4ICT8pFd
N009EwsjUzkJB6+uPv7QSsaw31qzb6GZ2pR7sKdlo5c3dgkZw6lf2SSKybOQDweC
34DVt/D55Aw78V10hMZCOc0Y1Q3BD1xbxQ7F/kXI1Ub6PWt2OfMW+tIY/jYSD9Di
+FY9+SzMJa1zpClBWam/cq7av3HiKB0HKK8G+CtYgSUCKpsdHy/St69QoADWbECg
9LINbBih1Blf2/kOUrXkiVr//9D7ljJMzDE4cGzXz51qVIhJfwuq2OW4KSKvuLYy
SLTkxdH9xP9rUYTY9WuXbPb0oO+ueFsycDvWC33kSBg4gyowe8bSvsTM9l3OzkaS
GUtq4AdJLdR4DLVivfwOGVeR/wQzU/A+IrjUskCWrfNFPE4BV4brQqaIPeDdPM63
Ys6ZD4g78KRTbmC50Gd7cw2Sa/q5GvxZi1kuTLj3TvqoX/XJRW8Q2pYsnTPcrG4Z
DinCjF/9LW/kNLTNzxbVTl/N01YSUkQrQjrdXy1ZFlPy27oR5hyoVDR1Axob2Gap
Y4dbHwewZDpy3YqYiplK7dbI9FfWdmPKdr2xI04lX5xJFih2bFXlnJY80veFVUP9
qp6eBf0Pa9PjCk0Ao4CpL7K0xYeb2I2Dd/2l5z64FXSZJsu6hPrQRah8ZDdQ5J+j
rxEBQt7pvUKrP1Jtlzysp+e2F3rEUll+BSwoApjRhyjU1K4JPE62Lbfx/RM2xr85
R/wMxSUxqNY1EVFR8EGFQS/ZYM4bdNhQyP7nMnaXR85yVAQ1cKHtwaJm/pSD0g/5
oxYNQ2PtqT7z1sylpkknUb2ozZhZ58ZMuqVEO7EGrBb8PPdGawDGtTz9/YlnAqwy
ZyePYi/r60+c00H2VjP3TlbKHNBKWOosqYPWcqES42co8W4DAj3Y/AS0QRnvc0qJ
CVBXGuUsMldSj4MMUwBFLGregPFOB+382ip53FUI+ANJ0IKi+96xf856D/rLRRwK
VKlik3b0es5ttfD8wBzbAjmo3PHHh0XF8r825oxb1tJHOCuFYYvOTWej3Ixkv3Na
1mut0g73+KEcEbGXqULcWVWFzBHvjM8cMmZQIlK38fhZTJEJq5QvqyeKyAoBSCv1
A0ExToMxasDXZX1tc7aANlkvWTUHpciWEu/Cqix5m3ynaQrjJ+S8ie7zqwyRR2tV
WcseAwOfrHutlkDweF4IwIazHdS4e92pfLTWjcw0SiALeJmP5VXLBWbvNxL+qzji
fSY/CimjPuB/ohZ9/x4QA6zFHDnboAf5VrdDa/Z1+Y2PKhR8RXQ5/bHV2NCW0IKN
iPnMgNUKGCOgKzuDjabflvf3+HyICGsJtjwqXj0ZPFZ8xj5DbMT4z3GbU8MTjkWj
6me/crB2IqdbRiur/G6wjGAhe6sEyjF7EiqADxFpCLQGZ849ZQE0qhKtNw0lDys4
VD6EgcqNYe+g5786oZtJUrYJPMKvOXSegfm2ZuJK2PpwWRWBKFwxzPZgpN5dd9qU
n0WpYnppfQ3dP4QxXqUJZ8gPSZ9jfajvgD50K2fggS4fPAQHldzAKzXwjFe/e10Z
JpcD//VAyGQ1npbn/dCJKjWiQnbNrM/N2ipm0qLIb08tYD5ofhvDraLZr4Dhr3u1
YQWJVJ6dPEVt7RTNhauAywNf1zYg/lufqyMUS/aozmcZMqlUezWtHSe32XDleHeI
ApoLj1/dJ5krwCmsHpxe/tEaaECA9x0Y+JW7JSem3HxNHmZuv0LPCbuPrrNKVoEs
1BFt8leUF1bC41jBvQ3oxjRtvI7ui2rJMYAC+DHOXjDR4/O446uqVzhyqPX9e7d6
2konnYaTHZSe7RE87SbEIPQmZYKOiXUw8BINT7HAOqJvlgQzbvPkz0OVGiM41U3K
c+l3/tje4dbbz6IMHq+7C5HxDqhNgUIYYuSNr0XEwPKnl8gNr0IHMwKfOF5r8vhQ
Nx1C0F1AN38bVFiLKD5UjEvk7vAEI7a+eOl/6tsoWsU72DjFv3BudrpdU5dE09OH
ckA47kYwl0TMnzSqx24oOluKp8PIapslzPAysb8sTZlgxXMT5ODKGOcBOougmtMD
VwCIPDu7rmAn2c1g4tFPEoDZ41f/Nz//us5p3fiKWN90PMG4Z35B+OXXXQFduOQM
nrPheoPU8BjFPl4+MlrU1GCerbIwpVFbbEZT9MKZkc6vtBWBbSbRk5T5+548Qof0
utofLESctCsYb/FekJ7OrYovNHrmrl0oy8zXCCzYs5GogOvVyc5sOk88+RGmSpQY
IkTdxItpYrqdvCrCthr4wf+eC6a9eGgoIN2kwmI5D2AN1P2z6OSQTntmf80c2OC8
qmME580alPI2RkPZuOUoCqkNDtdJlS6r1hGSjMvl6PDTePDEJjIOf3rrZaVu0qPY
U7SWffKSp2X3QC0pzGVLEAVhyTwZURBuqBBEIQY71rQGdCx42DDuslWOKXlMSLSj
EgQy9l+RVUt8eIe/P/3KHdCTPZF4YBbAe6ssNql8ndp3WTQvz3M4x60kcexHWjO6
8oQqgnzTIBszUjHjNSgmNuqUvxq/UJjLm/1pD7fHti2aiINRLVKhjWD6/cWwyvJB
OZOUE0LytBDPLGVfx/XiZwZxZ7MPqbSzMfINsXi8R5EaHUOvh/K/Fjy27O9geSdf
Zuhmhxj5J/Tt6vlYyubzW47sE3VrDyq6akklliQLoFtGzjocO0CreMo9I+hSPZzy
9uk6t6dvcubOaf+pMdAfRYFSzAMJrh625IRHPtZyPZunEydOLapE8Y4iUgx1pgx8
ZHMaAIVH5BPRo7ahjmjLmrGxHEIqQ+sbntj4L6E8u1hZrBxDVdnX62HzuB/OSI4z
KJ6xyyIPgQc1yeTs87pwY0EsF50qhW+qD8UEmrYJXnaN+YkrP9TNhTH3QFrJSzxV
86IB6ij3Y2TXFTHz2dVbbXbrEG6bLp7Qy4ePJj86BtTDRKUlXT6Xh35uweMFBoKt
2HZEfwIHI5M4cpnjaNWLxSNHO/WVBVa2ZBz815ZnT6xhXK6kVHgk1IHCpOtv6XVL
O9Psi6LGSpRKivEWEXGhY8z3WAcxXHFNjOuxRJ0A9iP7OIDcC723IPiEMJqjHXO0
xyw+kqRnguAAU7ysOWTpsdnU3NteUYfz3T3sR1L5MsZhGsK2tjQvL3q0Kt16wJXk
yZ8uMs1GIFfaFrZgd7RdMLtg3DhbCmsC2e32TisFYzCQLDNyB1lWQ8JiYEr7AqHd
X6IUFEKRyQUWDT3IIEDmRQ9yDq7QNO8Jyy3jDZ866wkSVLotrOqJE8Nt2yVlQy6u
wdsDcm4nBuTrxlEb1x8I6hVJKDou3oZ2yP0WZExUQO9mBuUEYR2s/tgv3nDCJXKt
a2EkKtxX6oPjVxChBZfJHrDZINbxcNYiEJV91jmCGwXbSVkUkId4MiKCgzJlpa+D
GSoFG67Y2d+AcU3UHeQKcX3bEoJBPlaXLssAriTHQijvzOg5QZ3iqMmX5D02M6ff
T2X4oRDHOERg+Ad54pAaInWHgTs8xo6qCU97QHESifW3p2MtbmsXU+EQoJBX0H04
c5/rdC2TFiOaI/Rb0LJCTBatNOBfvN/pWYQ/pn9jP5dIvBm+UvQWTmcLTOhv6U4d
iCgZdX+hJCHvkwks/x9oZgsEY3CPU9KBqbzWLyFA5/JqBitcKVRsCG/Mvxz/pNC/
VAbsLvT8g+bIBvGcZoE5ThKmlDrqeFe2m5gOCAFnjhFJoZ/8QzQUwATmCZf+ciOF
W9wdpba6+irMsufZYOwmm9Fbq+F9xGgzzFsD7r4kn3MIcYPqGbZki9UEIyTJoFQs
EoDERWTtHbobVyxzYvFmRthCShWztb2w8zEHexnvOK87Bb7bfteIfx2BaVDoQXdr
QA2acwZn3zTFoskQAgMdgcJ56Q1PRWXyzzyJgnruZoeU+NR2FfCLHnW1gf2Ve20Q
biYUTXjkbjA5eNXjdYNl52+RrlGnh0vOV7PgIS/yXryk81T9lYSJVQE+jSZ4+1vF
kB/aYpWwqsCdwejUw52NBGoP6kO5exeZrKVd3RchYJN6rIVaKlMpjfuwQRrMPbsL
kBgKqCdgzkQFeHlHcaFVS0tvagX55QowrvqD01TiosijZKG2d8SsA+00kDGnk0Gl
t7yNhveLMWwZXuqwKHPVFhQD3iZphTVO6WfZdPzo3XpIr5ovf8mDqs9+5xQ2f2Fe
+jTH1UVdrn3kiMqDvN6yyLyKOEg1mf9uEeX8LSWs5hCWU9qR/UMIWtm8XcfIJ9dZ
+UxX8bvq1PnW15o2G3q/7rEO6GdCllaI/zFW0+F280pwn2Rurj0oPQMMpdY4Dmi5
0E4uexONWnI4uquegK0OqWLHxcwy1VbNHCzRjeIl1Axmf+szDEtfsWUEcHLLqYZO
NM9SgNn5eSvl7K/Bbf7WMp9rhcXiQdKmDNnqQdngbLVakK1hPtHPCRFOMAMt9XW5
W8hGrw0ITKvYVYXb1345Vz9rWWKrpUcGxmo/11TcFePBj12rJwrVgm+CarkdKwgk
DkEivnnOpldykUwQyGttgO8rz1yb3wdlQX/LBO2lctAP/Bi5OaX3PfhQ+JAQZWi+
exLCpUnKA5fm+M9iSeASk1dgX3t2n48F+AD2JbRKRrSVPlaAlDLj0hFhMYiOQfLN
BvwbRXziX+F7g5HfSpFBiinMCteWe2TuThAVXKxdgaa+7CWjepUoId604m0Z0Ewp
GCNPxzunKEBOCPbh8FIEEZrQJso7nzKiFtgujn5mcW1FFmgCNo/LEjuyG2FIDGG7
1DgcMt/flXo22K6SRcLARCbtjW+DVJbl82Z/ZoN5yMQ8TfbfMY+bo7WFjciPCm5R
y/xSGwd8HXNg23kV+0cQ8FwHV14rj/WuiAn2728e6wr1Gwy1Ws9NIpa13OVPu1qO
DjHnWkCfg+ZcGiIsU5s93ZVOKVVUZ927EOwrCY+Mmdr7SKfpofd4n99BjzaSvEKN
nkaLtEAuyY/OHec69CnvE6iWuoPZ6z/5E6Jwhm40E5C8AxPgw2gXiges4y/YkSWI
0e/JjzH79jZyF+xkHjn/8K43WRqaul5jgnVY6P69Djz4DmWCYCrGOkwmKZnQbnOL
HyOhji4FqWSSh67pKqdmyGbh+kuDxydI01bVJf/YsneHix1FJ4tBNx2SeaPuJPjG
q71Qe0+tY/iwLChz6lx/K78eGaVLlCe+gpsu/FBdsewFBlbcWRW26qdLci9S5uQk
gQvtHAlyMn+hC9/ZwCQILqXJHusC+6bKeR8FrU0Q8vIiPhcwFkcX6M0WQnxwKOVI
5BPYsoRDB6I1rqZPiSTtnEgcRvvWVgv3sEGXjzX726W3hVOb+TTbnhYVYLyMfHy1
7QWdoVZx6xi08Xj2IEvj7/rABGQST+pHS2uYginJE1JgKYk6Cf7zkgym0HBgNWuP
xQoL5xbE82MRZtPhHKmtNF9Av9givpu/fpterfVDEam3qbvGCV1SDkkF9rf0RSs9
bcalIZ2XGOIB319SpEcNc3SBiq4Sd40N0tfpM2UbPNOLE73XfD/4stQ3POiPituW
xhw8jb8AbEkAXLGqMg+OmOGneIuQfBQEW/hn8UhANuUYLL8TG/TobtD++DAGA3Lq
9/K4sbFnlVwr0zEkLKi33qld40jd/AjGe3zrTvsSKpe83YvpIsgRaoR0mkl49JZ0
ZS5Myl3/SrDLctmLEoMig50FHC3pxTecSa8XZvf9p2kb6seKh9ZHgkSUz+EJmfwU
FqUa4ZhJ/8FNB3/JZjfohRxV0i2VZhixQgfEzkpgG+CCWfuFKpYWeCRY8HSFjSC4
6QEaofR0UsBWFrOIXdjmRK6iKAEiI81/y9VcG6sHZUYeANoNYU5vcklwoseO56ED
PzpJfcxa1WI7HtanQ+T7wJrZ5OwBKVwr2mCK9283tjV4rCaZL6g66MPiKiTnbTnp
xEZv1iisi1awgpSdovJPRxwBlJDOQes13x0NyBJ7wioc+OICEi5gc6YZmhlhpp2q
9JhRBD/EBLgqWDbdGz2pANZbWbKi16DDnNulQMHQ09zTelGoUYWPNHVWxAB8bSyl
d5/Z0Atphf+7kZRLn3YS9GOcg5ADv7kYrk9obd4LXZZ2qivjv8WkK5chMSonUROx
vbYpCvzxDWuFjiLGbQNTZwo3c6iR3pbAzOhCQ5LSBOZ842Ns84y2VfGrCkHJoeN8
ISnslLvT195kuD4tqqWUUmulUa7knB0SK7VVxKk6ExKQ/gfl4p09niz8CaTJZ9yg
p4njVbqI9tXeNo8x+TblyJxoRjRQEGnitkG0fLdj4vL56F9xlWAOdaHx9472PsWK
2vt/9EHzSMp8Kp02iS1zq6RQphBUJK6SCYWJPSPd2j6HMvrXt4uy6wXRFkOqWQ71
EWo1j7sLSsEhDNPr/kl4hjpyaKL44cvdCfameaYLMpboGxCl/OJ6JmhWF+sGV+Qj
+GOr+ZqTSlSfy0syvW1k6qGljKVItCQZdQ+Qsi/vU/aiuCrhmHEjQOHivIbHcAnK
yjogLEoJSvpSwztVu1hW9CngQphwCNoH0RpdQAeLAmJ3GsOys8hn0SotZPLiOPpv
cS5gkR1+NvdXqgKj0crBeTRqcIeO2Y999N9ZmEsKWOrNRHMpWhZNFNaBKXmPKxdc
GSv0tAa80tPxpzP0w+9dHIRWHorl1Q/FFuCUbNZbJ8oJ+iZmk/nw7d1wPQW79DtV
4TOAZ57xrSB+OmSRgM4Jg8AdpCf8bYgo0Kq5WfU/IWEoSxwgUtssQGMLc5vlevJr
EH9cJ/cAYp20XreUYVj6qcpFYqQBIl9rNTuW52u+hH4BT50GcAlE35wfAU7M5whQ
Pjysi3ZL1suzX0RkuM1V0jZN0qG+kFkNFRvaHgnAo3a59EAQG6QP4kk2F94+LBKc
tORnbEtn21ENriEQML7VEGgLMHN3MPXQWdulTNeUt3Dh/NCIiMFHMvrbzd3UPdUT
BPHsFiSHtKbN4L15yMGCIBSrRxpPv05h5h/sjUfp6x2CLdEJn2FUC6pnAt+65TLg
fXJs43Wqow6g9oo3cs0QpDbfAouMJjFji7aN/f0DrPIhyGWdfm+xtk//yj8KlFwo
/gjVzhWrYbu5yGCqwlgA9JWixzuJHstmUOUrpcHWtWDl7ppB0Uh6U/KWVwIFCmbk
eUmVxMQ6DT0ZjkE0AvI/R3YAV3UfbJQHm6OOBa95gt5eO5QUBHAQ0qN++GZdBrz/
1z9z0+d6jzaz2FI4TNndOD2bGKmeg455rOgqQaVffHpJqikpJ7rcDmU6b+LW8Q4v
ps3342XwG5D35KYmyd2tuNEy3YayIy+044M5xwwID2mpUl8tdFvP5HfJwkaBqckI
sLutoSnVlBY+4s1LTVsHyGN3O/KwtcyQpUbyclquqac6Efq200G9igahVdFu8cEo
qkoEO5wbK4R7IhwAQvuzvO5sS4bqCWkad2H1mZlXauODKTaEha1wCVHia6wxqkkI
1t4LbCHFuqYumcZFQY6ZRQucFs8JKT23RK1WZXGg759T2z6Q2j+Ase6TU4LiRzWI
rEWeGDSt7hVNChvDVwhvALx/PDQjLVCbmo7CgxTT5uJYUhF5giHmY6/lHg/sW6hX
ujmaO4OGI01nvbQ1tqki1TYYtu/nd67+Tmfqzik/C7kBiGLXxzgLQq8fTzntfdJ5
qFUW3yRyo2xC3mA7KrouPw5RBwjuF0A8Ipy/aN490N5ywcOfDao6O1WiCg9yedij
dI59NjdOygaOf08OV2iudg==
`protect END_PROTECTED

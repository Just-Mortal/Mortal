`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yMnPB5izGdHSZX1JtwYBoXM4+r7fTAociaatUKrVQ1IyogMEPiZFo3lX7Pvy/FCF
OPkKLUHnqAb/Ah0imfD8R3D5w14pequGdKbJ78lkoMdcaNZHr2WY5jYRb4U01aQp
dhKtgyh4wNGOIeT8o8srl8SIBRUUV0TAcmxHmS0s8Hbbd0Ke9Yec7QQDvzVyJbjA
uFkpdZFnIXZZu0nMNhtTD0ESlavlz/dKsVH25WtCgUp+cBkWW9FbM10M1EeSbF6H
uOOMZuHxTSOqJ6kIKTlR7HugX4gljPmZFdnkUta6Oqno5ETaFSvdd/A9yu4juWPn
NCLMeLfQrVzrt80hHsa7xv21BsRKqtYV8+nzxvY8Vo4Yh7jw5F9AF8JxX6mvkQih
t9GVtz7RatBmKVnfotATba9+ZkQsfQt3+WWSQhJQ0Yr1o4VZ/s8b3D1QEd4pggXj
6DJt5sFeq1B3x43Vpsf/3h1Khnq6BZ9oar8bRbYXgYe9ksvAHwPL7TlWAgZapAbs
RwknGw5wJAL4Q5otWbCOv944VUkDHgoACxXfkPS0CLLWyzHy9pBpVGSIEWqjq2Hn
FngedwLTdlD+uJgOx+RlQQRWAUdWRhJrqybCIoYhR18MZ0PVuSbUiLDaAOJwBzQY
kT4Uv+Coj4ReLxxaR4PdneQ8YX6BwpzW2SaaZU7szS8=
`protect END_PROTECTED

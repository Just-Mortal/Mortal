`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/0FgCUvfI/0b+scnurd2gjfg6+200ePRyHhDBBIb+I0n4/qHT9calZZ3Pmnqv9yX
HikQeiSv3wDhNqwhnpoTVLWBHVNC4yyKoEvZJzYPnmfJ27I/wQZUuYAXn8bWqSQF
oY3ILrNDuMHjSt/bHlUteGwwCoHeYstrj0FSVM2fRBRoCYgq1u5wAI3KU0Zex4W9
w4Ov+tLBrngtKj2eRXPD0GQ101/qnSfGQAURJhId/31RAJAukil8pfrRibSJ1r8g
IzuhSfSHoWXJiIKN2cKDGLQ+N9yZqiud4gx6Su8G9l7BQ01wQssNWDh+IP9M+kSl
Y6ocR936557cjBOqQ5y4PGjLmN16z1ZI3Yy7dsvfo8l83rcq6sIL0ResGHRpgrHc
9cu0T3ddzx1Zl2glFdLL9sRZ0oM4woYMgjSaLqei0kyCI4gqJIg5n+ChapXVaSK8
Mi5nMFpc0TQ2OmdfSdPKwldFj/9w4kc4YH7fi3MBaPPHlY3kXAxLTsGk8XX/QYAE
eCMgXsk57eSjwyqSeOFgJyay7eclzLR6RwkCWUwNBHlBBYnUyKThkhQZ04CNkhSP
jaTxkkqFG6wDWYQDdxiruKTeiQq1Aee4zPBnxJINMqvyA+f885UAntZQTn/jRblm
vy4hxbaw1vo2x0OlAUqkjHmRw6pnIratk1OmGJEFRNh5dJC7iz09R6TybdSX/Yzl
gMdvXCvoCi9Rq9u05vPUMmYNzs4HkfPQXLrZzRA+v+wmPb8HAy4duU7JrWNNuDVy
EYToyIn0FNNQKLo0xw9SIWnn7xZWJWldj6p0qoODOptfKWRj8zfd/2bOV4tUUaQG
`protect END_PROTECTED

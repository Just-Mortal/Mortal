`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0XJssuZt8PrDlMJQW7acoRr6xy7msSdyTC1JomwmhjCNzLbJYiHnaiUXS0Hnfrd
O/DufIXJ9T6ZwqmeT7G2zC+30piJwjaeAHwK27HSP7w9Srq124RjIYN6IVd6bxHv
rBH2uIRURqT3Y8gh2rj5FI2yLzPC7y6jDQ/ScL2LI+1Ay9R41f2ONV9842UxX6hc
Im7DK8eHfueAjBJZORscyaB/zIr8pjtalJT7OBk9zKZ8ajpJk8vutSdKyDbL9EGt
Iac1OU8PH+xoizPP5qx/I/8/fdzScTDfqGrXljrApgIjBUtRLGfTq3EHc6JVGSGQ
pQOcphBcy73uNdhaOykyzeScvr0PPJL8j8n90X1N+u5BWAb4ZPderNsD73mIW2rL
a6ctBkctu1XDV0UUwLltJ2BF0I14r+pn2l/OFpwJZPMYBEmev3W+Vrlp1ohavuPz
jKr+y+oX+2H9ePqz+3C8drsbTnnk0BxLb2c4G4c9lBssdK16BtXZAQ6mYWvIAAdy
tTPlEexVE0THdf+q+eBXRAtEii4UbhW6fJGVPNoq788wbAZnLw9tRyfuPRGjCj6N
CaV4CE7Wslsm0/HUrTJONgziWEk1yb+moCR5Dd4DwJsMTvCFr71mbQvRzC3m7cYd
p5UoyGvjAsvaLVgKQzVjjCBgVcXyr/Dr/VndcgTHsfk0BCKrgGuT53vOUK1GUBWC
UE1XPqOeGPLdNbWE1ZynAG7JafEvq2RnMSTgx9eh83Lrc4lna7Qd2P6PDKQQeMvP
lvWKuNa/IuebJlt/ZE/ol+KSwJHo99wVxCvJ2I1QLFR8IhlqDgvsPQsUrldBx3+b
yMe7oPGwTTsjgea7kxmceIIcnBErZSwrMOKYKbecqCAjUFC0XA1JLN/cZt5tK/YJ
esbw74Dgg6KjmQWIJ08Opock2UFUzex6g9Wm2supDYC6DVUx+cYiU7gIjSavnxCi
Jfs5Oa/rRP3Ved++mcgQq4z6zQ8kaiPlDtxZnWSBBy9/rgXBs3VLRjjDSbdJR6bi
GRj1hmLpDWHkqr8yPZqGuuvFf+wZdQnoA2KFHkd1ojzN8udYoUZW5jPgHdfoex02
enFc2q18nV/JXo23sUZgmUTfS3sktcwO3dPzuYrlJW9D4nNrGPXJgaV4jEVXViSN
DdNqxIxmbAWig4yzvUo5aUioySdTpiRuJQlNuIfyngVoBgumW2l3qD4X0oRD8rHY
+kkseRO+ZvAYwn6wP9kNaFuqTTKrC0LFeoWlNSRoUPOVztyLUFUbVfrSlNPhJHhT
mAuen9EZVQj4twgVFg10lg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5mNISEfmMafRHSaXjOV47twMJn5+Xl8HQzfEBJFg2JnxXn9LdomUmbPmFQvQInVm
zsdZrU5SzVNcXdOViQd7jif70/V4Al+nAL92MiuKSuwGa3/0i6APPM+JVOgN5Hqp
DNGvplA29TrVMz549MynL2tII1AVDLje5UOHRavL0vwbajX4h7HPVCn2IC5d1oZB
U17KwjzSxtbgmauSqY68XnyNQhtF1CEgh45M65FbA7mJY1XcusTwKmzdWKSYILIh
qDtnyW/QzqEyT3xO9OfovQVu/vLaZ4sHfUqSNn5Rur49aioWfHD/AQfDvMDYa034
aydZFJX+gFlbe7I3k8oxKYaKneQTuhoI4j+Ppn3HDpq4I6bkwy1Pw4f/NxwtIo5x
Fk7mbJmVfSmyTcaQUqrNeRS4Pv9zxI41x3IF0x1l64cXROg79FTGxS5+Z47o4rJ/
3NlfprCoKHEWhlEFXtRgxCS3Vk2RmUTuIbmRH5F5NSoNlBGJ+Xu3A453ioI8RD4V
rkdoumOaUmIKCjG49tAXxZ9sgf3wQO1cq03gGcVfzqNbrGiLHyrvH30CvITEC32L
53oCGNWmxL0R1LRIfLC7q8rXeI52cTUlaJXrfNb1Vx3DdWYyyQClu2iQd1RctMh7
kLtNjMyYXgIJeXBawbAvw1G5T/nS7qB+Cgdnyg7roPeUWipgVVmn0qOsJJpg0tvf
BhnF7T+oqOQJfcCUqUZrwKYwqZlEmO61bOSWXxHH6CGODkai11aR9igJ04aa9e0z
zR1badPQmY6ZIs0eLxfCqs4lF75Lm2pTEpaSV9ayfyr1rxsGpTBDfSXXMxdm9A4z
FLLEryfLBceQtHffyzZi+l1XbjaStthmrrIFQ8q3dzORxH9OJM2RPU8l+TbAK9WM
drpOOs4L6ZRn9nq4v5LAvEV2cULJalyXYKK4i6cqnu4=
`protect END_PROTECTED

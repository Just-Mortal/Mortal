`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CFcJGKni8PJmhylp+GnB8B7jwxLSJyLDep6xS4lyMkb94ClaRhpRhM8OwWUoiBGI
RrbynBdEcgSFsRofriwgGhc58EX+F5+Fe5jH0Bl91oEeWuBg89cL+NGuc2XaX+Gf
ssuQ4e/8O8VP+BPtRsbBZL+0Vg3s7d3WgU5RGlydg+Z3rxFkdzNM+Og5pz1rmVDd
rjyvz0yYO01hIui6Sm3QhZnas7v3oWn+Mahypup2PqhO3KQDkiUrMAGfyJsmfnME
b7UlvE2INQ3x38v9AYq/k8quFU0OVTV6CBQC2Cpxp0EsYPq1a9TP4U1MnVfphSdV
TwtesULxcdgcx+OydygyQ7+OMuiHrLclaUrCBQwegv67pX6Tnh2N4Fs41HxbPlRg
waqd1hj9owKkM5GgKkvdP5LVABvnTEUShOgaMo9Aw9MICPABOnD4QZChoSOXOEAZ
mJTQDRo8ODGKq+F7eYWAbbEhH+h1wmRUXQdOXrqu8y1XoRZq4n2Id1SsVsoedWty
6KFiXx0p/fDJU8DW16FdEuudvClYLz7/2kieTm8mv39ZRwtwlcFSp4Npu/nwly2O
gIRNg2B8CB/63xAu5BkZLZPiCceRKFgml6TQ/joTKC+O2ZKxTIVzqxf1Zo/rbD3X
V3q5q4kVIrm+SF0JOjNT12VayHhMX+2QOJTNXRyIdb0l6n42fMF0ZPkeEL8CSMXb
M4CG9yWhLeHkeaWyQYUfVbcBalh53QjqECYmYuH3+51GcQdqkm7/LFM3jtp02EuW
ptQfzgNfecS4ybb/YFxzbGb9wYWohEIJcK1mgNxlx4yhP+gxydqqn+aIXwAZHti3
LN/+i35tn5Oh7rOg8FC00Shh2AuGqQnbWo4CRkiipvYQEZEzgMyvkKHun5lE9Anz
M2okLc5ZCHCTQE+odmUOZL1dyIRQ1vBJGW17GiqdXIWSP+qnmkDbueWtxxtbhxet
bf1z+/BF5EEwZ8r3CzXJTNY1rOYG+dcnJmGCiCgsajHzAQDa7yJUOwV/FYS4JlnA
mNJRqvPEZqPT88K5JUXFC5+035fP2ZOau/Vd82wKxe/poZ4UKRQKrH1zGhPpXT+5
DhcHM8ROtHf87Dk5wA6ZFr+J7sISqpgsXeIo6xQVDgd1cBlGJT4fYR6hswlLhRQG
9IDmODFy23R8ZhaqjozSPsFSIMqMm+85eyIwQ6a7+f+D5Qn6AgUujdZjrv2gZTCQ
t+skwOJPRKn7AYnXQ29fLcItSX2o1XQAEEiHHwIzZvfXntKaoUarTJsHp2+Tw1qU
ln5q8Itea6VZvDCbnnOEFnj1lnUVmveen6fTkSHSO3KopV9vHobcRTSuBQV5xw6y
Wk2Ueg+jdRaJE/YeDQJoSe+VwS6q16E9LEmTor/di1i9YG3FdzMLf5En2gXhx60g
xfawutLRPM6R0cel0xnvgmBQzd3i7OAG1ZcMvUM1kX1JXMtKn6XqG7mgF8EJ8Hoj
yxEi6ZD7ZUhwgZq7kpRZFoXi0QZOKLWxEcI3KD9uRSlkDa5AenYCgVeNiTbafLEU
pU3ouU3Z0qy+cxm882EXkgN0r3esQBnATZ/Y8y2l5DKih/1l7fhHp46jczT+9YM+
yXulBk1DP8URqgnGuZWp49z1yjw38MVKreSxnQEhwbyr9aU5Jv0n/s7KEkpePVH4
NxHufp39JV6KRg3sASbJoDAcD8YADGF+QdcawVUtgeuVCpxXLLu0WG8YVr473Duz
oqHEfzRiKj0DQEVRqAaQPoRm0qSnDouLIFkFVieHkJVKA9J/HqU+nlWExZEI8M1Q
j03xuE2QyaIVGIRjrWk4KREQogVwYAeSew3C8DM4czxCw2slvR3oWLMwSx4AKcMf
Nr45wfjRKZiwui+Ogkp++LaQJ0+hoJ7AmbunvRBieA+XgPi/de0/NWq6ML56LlwR
PSlmWS3Qm00QeIdyVqACXiy4stphWXQwDWIJ2M59YvQ5ELrAAjxVusapFD0bf7EC
CiHAGfVT3z7Iu66oKheA5Bqi4ajCWM3roeNB22+JDZj3LmTyvOUQELPOYdLuSReb
3imRhGaLXE1Vhzu8mL/6+HPBJTb/GNWD/Mf4vwIys7jm8O+7GhX26edobiJh5vdo
rGmZtR6cPABsK/e398tVY4Dbq5qBvMD6nUGwJILF1yz+/HuW6ykOElrYKWlzQbFc
L3TXdKRk63huLtUGG8XOXa9WZ3y0WqZHYVaVzfxG1/uM1c3aN5gvoBn9ZzMjQMu7
UrnFlzzBLnwjlVky4BO54fUtt3e+wwRgrlbuU5xadaugULUi80/Yz2q83qw24rwL
LmChGh8w1fTMCgofZxQ/iShDiHOi/9g/9IFzf00ciImtSnOTokk63Pm51kwqGyYZ
pq+h0K+BYPywCb81oHcP3+hhLPkdKIFGfcqzsc7VTwlpgsb6ep5+KAmABux5RlZG
snTnhvc8gKr+VhRKNOB8RGg8GwCyoSkHAkfRAYbfM3bWQ04Er1lHo5vShbcokDW1
FqACJTsYFz1zkuXIV30ZAKzsrgyoj0J0jH7QXqHmlrXk6jwq+cmF9yJoL8AwksK9
AaiTeN9b4TouNpYhl0xcCtEcslVq5I4bdW84jWzIiiH9BGrT+0SN0qJGJfr1Klux
cJh7P70eCXO/aVW5Vx6LvHvsc8dzZ5h73eaJqflehZYK8C3s1N3WbrFO0CBGRmmz
X70ZhsbDR9Ra4rrEC93Wof8Ooe3gRFSKlbXEuvmIOVkZswVpEFTFYRmahhXLQ9L9
S67bsN33O6VhY2nHkm/EUvm8fOvNWYlihSsDT8fgwo9Yix/AtMSOMRC0Uq4jNzk6
uymt9YHa1/tAM97if8OYpLl3H/Wh9075AeM2MGtiXrjRz/srMCl9dUz7SflTtF8y
3bqLl3dONXyc8XBfZ7f5WwbZRewg/C4Qa6K8Wa/SF7CbfX0KwysFHzJKrEQYZT5h
DQkxOASkJSSJm5FFNd60nyWi1bpmylZY8Dxgfa49MnSvOxSGPu6KCYkYN3oM//++
gZbVKgFmJ3vhS6Hq4LfMEeOBFptLlv+PkRBVU9VbYfsQ5ZBhhatQciwXrw00uuRR
G63JJGRQbU3aaVyhXu2pcxMepiLjozSs15m/yPQunl/vo0KCj/JNetoTl6TicxXn
HFC5PIu/HhXDulu15lZ9+rWU5yHfF+dftZwEq6nzohKJyRpuSHB+DHsSWG9OILoE
KbXxTamYVPSHIMMuhQ9lENnlXHZJM4tEQPOwvXI50KQ60vUwI4ijvdhnL0wsSYDa
/umFNDl9L1IpzSY7i+TrnPRia2W/JGeEwuNzgJltsVlZoCfdvOW77aBVOoUC3hhV
Ua1WXdojd1v655CJrPa81CkLagYVARM8n8Yze96v4jDivl7Dp1tHyUNfRIV/M+XZ
+fIsAkF4AHGF/TFeF75kqCKZ21Q+OMGhaWTqYSLU4ZUNlO4+kcY2CWAyBgDJM35Z
c8BYnGtbYbYFLiqUtOtHv9ZJtMkWEbPo2VFWSgYLISKk3fWFzPtmL9/5EqDHnKgH
7AZUbNKQfiRYc4NziQV/2HBhqBYHJKpDgI+Lf3I2r7ZlUfr76f/rrQ5pplSFud7v
x2c6PcbyX6X3dl92V1QZDuZV8AWITEjG9NPPTfF4raJoxWjtaYiGQTnIkMGzE8iT
sSS9dbDjUkqG1z1NdJn28KpgSvIslj6XNwWcuZAtOYFEDkpjz0hoFYlT+EGlaQiC
+vy7Px7DZDClHl3/7lbihuUlVnY53uaRcCCw7nludAUjk8VIkI/m95mom5rT91qE
qSH3M5iNmMF3e7ns2cKH2yUJz8KnU2wxdXiLfKG4eoxFkzn8uWI5EyJjrk5R56M2
6YPx/dO3bgIm3zqxlj7nkdGb49k8Mpm7bqOcWiMNCpCnNzWHKoIpcPtPxaiHvKhd
hS6SmbosjN0+JOsePY+Pjcf5rpLbQKjDRDnqIlnyqYwYTqjFirmmVvAAQYTc1+Gm
AFXL26AcfeD31ZBP6ijTihQV0iebb/UOSUDsrNIRDek2xM3SDUbtMv1pArbaqNZN
/ONh1OU6+h4X/kGx6EyGGGrnS/zhF57Z7EJiFsIxOzeiWAxWcuthD/YtgLzDNrzy
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zt6l1NbwOuk7Ny6quBKOM6GSFOOoEB6u0izPK2IEEr7SlLwUxhyMgMkgqUIbxgoB
G3oJdRWUzNKmSR3qyWUWjbSziQyQuItnSe332fi1HNARfdNUP1+YAq1VG7zgTvUx
kzHQ7w/uPb/F7G3S3QsTX9lvK/8pPjv0VU+C6SDu73Hugy9W2b1UGiCaUMPxub9u
5fIwSLu9prIVL/IFLRuwsnDh/DfsqrqVHkjMpACFoAqiDZH7b/fouTfAlumnxZKQ
mDXzSO6SDPYxmZiBJoBXDnnCiAgQjcioYLTdPqJSYolwU20ld2fmK+SUFws2fDMT
W8h97MJQ2z9FNJyRspdh33Hraoe2XqOcAhewFFjGYiRmQmeYRJjwrkZrDQG+YV4A
rtrKnkAl5gAYyeGvVK6fJMDpvmxaVqfYDzV8VG1DmogY7U9kQqwYb2rlBxikF+zo
0A7n7lAmU0gthypFjivTLvx4yAt8ki0/Czf83jJzNFyJxE/f46TCK5um3dyOAhJY
koRpKb2RJf3nyBBntbIJPP/monQIfywx0XRFiEKd3SZxcS1p5n6OTNtEG1Fa7URj
WgvX1w+m+YR/fBOx8xrDTFzFXSSwfqR+Ci+CXAWZUWaHfvFu721zX/669ynN8k3l
pZcGWzWS9JrK718X08YSQ7ux3LmbemTiCRJm/qnrvGZJzw+uBPeZm4o/Atrr2ByA
ZZc8blOeiOKffvHgexfUdLVKM732c+oZUGob2Cdv91V237H2raCSKOqIaS+je84o
uChsBhk5e4ZW+0tpiMILFtOz3+c+A2cRBKx5+p4DsL1ute9HM2tCnoiJ45Ro8oir
9H37hoC8SgHEbV85apZTA2r+q7SNidPfXtRIXE3TT4D37ZkI5oVxZAXgdYP1Qi+g
sylIPsw9k9QB8kXueEcgmhWUoUuwvZbdJSPdf2Kb+YAIplOTp6Sd9pC0EzNiUbpg
wZ8Y/W37DPbCfuehSR6u1Ky0pJ7kCxAFQ10ovqaSeTIE6/uvTsGAaiIg0o7IemlE
zNskLpy9MwJlfxYtXizn1pYrlxKBO7vfmv4Ju1rEjI6eOJKXW7ETH4Vj+2X6eRVs
EdDiibREOpiQ5Mkd2YFsaD4GHGd+OV/hgUkRA06wkNwikHd3zuiKuQseoXwsATmD
9xmN1hP+LngX2Cn0f5nOEix/m6X+bhpN5JrO3tg9ppNNeWKN4vD690aqGD+YQzgC
kRgZ4+GOOVWCK5ce8U4Uel1G/qlqrCFX4+xRjkj1HTELwimsITCQCPTSBVacF93J
A6ayQRJH9qGpIu/lhU/mHpTFBSbB9I3t2a2+jUuw8s1YVZgYbGHzL9u9SScFUvrE
qc06W5WD3nUs0U/0zVGSbTvdZiqovLrohrXwCgPhAhnQPvvPx+yVZJ8ZnCF72l8y
U0SrQcT6r1OsN/mOHFk7I+2Wod5AlqP3QERps5/vLXUYh2Dw7YBGv4hkoqsknz1T
jDu8V3pXfCA1R8Zt0KoI1hPIKZLKRjgGKPTkJ6eGb+G7jfXj9+3+jU+TudWMbuqn
JzVEukYltNNU3hN/UNWJ0TiTp+Xb/tq5RnblbMTQQ7GeWcJ6ivBcZopY4Gtxwe1d
qgv/D/ztiA0fOzpQWIDFMoSf1VXF1opUAevT0sFDikQ=
`protect END_PROTECTED

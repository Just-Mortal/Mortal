`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zceVHpA727fAf0nyg0v9g2+6X9YWAORQ07TOD4gU431rhfdlvQP9P5hlxHeTnOhY
UrDUqTrxnvIC2oUz0fj0cjkl8ezjoKY5+8oRB7Tz0xOg4LHUE21oyvdYTOsMMzbe
iVv1CDT1Qckx5aSLsA56WGWcKAmuMnvoZs8oGPKzDfVaQNTE/tcMadAiJYpVEBsg
1EU9Xc61WhzbELJmaXu0jundY3BCx5DHrT3DPm5B/5Q22MznUAYRie3Qm7Ns2k/t
DzfW+nwJvYflgcEJI2WWxd6sgO3Vvg26ylat4gxFq7CTaVRrLkxkuniZhtx2gjsR
ltsbTbTbii93xll9cRimCyb3oSdcHcyY5r0JL59g6/HdjxejlbaqxSgGpVFKcHmq
dKHBF3M2PqaM8bb7d+4W2pNgauQ2swsXAyHfs+mhyg/l+oNchQcWPN/FkMv8ExVj
BRQPMvAzEvT4I4meqFmUKVrBFrOCMb1YHIrkERRN2lh8cwV8yMGLlaFmTuj00jCO
4ljOsy3j9fQWxWPIlK+h3L+s/xSHQxvIxcYmEuMqm3oR1yNoorWk+wRbMv/zPz71
cFf3+FL7jAg1NRymrw4mhNCX/Enj/ZzW7gQJHuyY+ini0ltHpD9tc5HfnJxDWiYA
VrqXCE9SpRd4s0ElV4/e0GLbfXs+WH7sTaQl8Tc1IFKubF9G9apa6uTiak4x0HNX
jpZO8soEOPTX/XbxNyQMmaNXLzb/4KdEFhazzpM6Z0/0u6KOaDoxTl+HQx8grXVf
1DchtEg8hB3MdNgAqMp8+R0Lj1HTagzwx2vO5jlXYe22/kzRhgkxovbT2MARloxh
dnvqVyPrUE86s/xZoRGrisgU+R6A2rwvaeIbzN3CaTwDlRicpBmwd0IiO8zIHdVO
q/6LllWnF4EdIFkP7tgApgw+TTiiC+BQjcd4jp3co5XEB2m8zo0dVZORgdkiuPLb
HEAxU/cIRNEpeZAQZCMHDGdq7ARcLXisjH3gHA8pDNR3/IW+gKtaeE7BOaRBrs6R
IkTo6nyh8RsWBp9thc3sBEz5H/ZGgpcwHadjqRIXJvn5bQd4kSwFabxHeMrmWkPQ
u7wlRtERO/qZqMcDcm2hSbaFk/54/R1zyrBP1TJiP10KbGjwziBi9d9hHfMnl4Wz
p9ZkkPpUqoBt/XRg+Km9SVpXfRAz3a234TbmplblSyE1ivDDjkXcZvFJzLC/7O7w
t5j3jif2FeqcdokOadm7Y+bpd6MVeXl6Ze835MQv2SlYnbbeVDgSvF/6Vt5cYzNG
9qE43YK8CeNf5VpY9ij1hM+49qW7tvcRJUaGZbQBu2IvSN/aCiUEqoFi3xxedxNF
27Zp7/CG/nU2aThE1lctTdkBt+P+6YeQ9mcDDCJ91MixZzkjpzFifO7R8zgf2Ih6
ZmMGAHuxjXamsVXa+Ae/XcJMtZa4Wm9Ta11Xi2FHH3+NP8LZh3M21mcyXql2EEhx
RuWxpjqMlHmAzPMLMtrD+tDPY1N1XqCzAUIyHwkAtqT1tID8WCXn187ItkTLay5V
DvZOk8EurFDWG4uc9DtPtqTsP9KT8RJz3aBAevJDMf4krGGd4udy/ANps8wbFHnO
JazNWONSVLXNQQnUXso18G9l2WpCTE9GEPbaJio2jam4S6Jz3tZ0botXhxl+vl2D
O8Jw6Z0atWKQQCztFTqe856PC7wk7vU94ZgRekwbw9BprF/DDLr6qZ2SEIbPef2S
rbcn4j2lql6ykiczCjwp5rDf+1AuXD/Vl0jYrUG1YuSvIXlO03oLvDGs/eJgurZN
npTwy0iIe5Frux2mlaE2euhbMOnQDvy9CBtGypCIByLnZXmAA0MfQR3CkTz46ddx
ZF+AZBotDbaxQ1LNNNEEYHp0kPvbJH+X5agFQJzH6aWCkHZCK8/1hwJ00y7DibpM
G9XF09SxLmQpSylCjyEVzhkQ7RuiAeaZX/wRcvw383QMESddEnugHd9v0K7Sw0NC
9/WZPsbTojPBaVVmOmMyIQjoyrV1BehMsNPxvPOSfVlZ/bohwEVJhdt2cKT4t7Nm
n82xzYwHbcYfZDl/uVEhSJOcCYRqMGpk0BEYHk7FvsGv/OQUVS2UzRfr4IPjwIjF
HlW1wT8fX05vKIHBGYbviF/H3KJRJylb0nrXUKk8dnCM2ixrQxazvbzs77lpdarM
9arEIDFnbGA7rWWZvKeK+/ASanuOcTNssLQUFpziJ2wFhbRqvtQH+ZUT2cEOCPSY
Tg7PYayYe3qB/ghWmau6kVZpSvZ6E8KGXOXtcs86/ERGjKusSFz0Ztmdxd+WSu6Q
jJy2VbTZPHDp51G/lRhqrtdAmFvYQkCVC96QoklCP/wcFCPjUDYjzpl44Ph1Qy+y
AMmEjJMczNTspXRJ8/XQfcAktAq9fSXYt1V+2ZKsW1dO59BOP9HTiAntHLlPTPs1
8fRBBlO9ceI4nxyAA20Hj4JU+RVSHstftdqa42ZiLIJkvOtXRhZpHDXdEaKKxTmL
QIV8ZNx0jqw+pFbWUASpod6/Sv67PXPmikkzzkLcqLOppRCTQhUU03lFbsIzYCRw
l/1AYrBrJniO/OLBMkJV9FTa3cuNT3Q6Eg9Hyretr3f5nrnQbE0C00DSw1GkJWLt
N/C75SY8Fss1f9kwYUXEkQG8oFR7yw6eHsuU+8yOzAOVYigCru9IxzqnUbyW3oI1
+pzeyhuIugqwEUPtuS2TBVjv6+Ev9sWyg2JuydthbLo3dXmaSEr+rOpkR0bGxVVH
OP4Mo21qmgLoeZsoY83QOGRHAMQ/08cEdpki9GDzVSq83piYSTQaihFNJPRbBi5Q
An28TCDOzzSYMszsdPqg08NSZgpaVUHTM5Y08yPYqO19nmM8kNFhOomO/bVasMlM
7lv1zOE0zMB5jECfbuXE7tnQgTZzkWVTnLIcRC3E1BpL+y7yBJGsWGNDSmwHQ1j/
PIdnRRSVGPlBJX45INFMg27/C4ITQX8IXOfAM+q5D2l6zNIZxXHbvo/RNjZFX9vs
oreV8PIsPs9ghPowddzuMsBU8fEoz8Da2DDQq+yrwFY52WgonKXJjwI2CH9N9tDQ
V47OByRzhwIdMFJmA7SB7tm0O/bz2V6rHfGdGXDDqWmUiofQF0Azb3VEsLBi1y84
aGM1AMwwm7z2gT2v1nCGAbR//ZP8NF1DgwtcYK4LNkzH0pFkg+68ZT1hJq6zcnBK
IqI4FlqlsAgv6mv3U863I2aofXHnx22wnGWiC31ybwbFr+1j2ff/2SeChnXCICMt
S5D2eCXmIRmz1x8nAjGL9nPcjUAkFGMVqCczS5yWtN6rqrulXAGS4bSX2gd8HGub
yakEqfYbyPeg1tgpT6U47MwxJ5HpRRb+l7XyA8rasEsjSfRCWTcYLkjgbAWw3hi5
CCdNSFj8UNDqu56Vv7Pq2lZIea7mkDEcr0eqRRM2o27w4f3bBTleNbtD9goi8qfn
/CW3GNsNEaYv3IEbLE7hsxI0GhxWy11MSSXkEG9wCmRDRhS481EaLj5lAqY2MvGc
oL+vb4q+BKRerIc1oWo/c4yZMC1R9npxgf8qkn9DEDBvtKdmDJurdYnaAuSQ7oH1
tzAOn2hNnGQHrPx5NvtRNGm2bhmJrs/RFysAr9ZBEG83oQ1GahrwiISNBxNMYEYo
OUd/7GlovL157yziU31j2JZLmY0jZs4Paz/eczH7b8ronSiIkysXcm6MNNv+upx2
VvfTkZiFeuBMSQXnM7GfGZXReABF7f132H+pg2Div7fVEqcyU65oAADvRmQBKRl1
euzhhb0ohhQq417ujqSFwxfLaM7uGKpD/KEmDJeqeWw3KXSc0J1MpS3u7i7RGeR+
jNA41BAX0dFbtG7abFLIXc7mBwh24vxptfzAAzTROKEXXpu/bKkum3nkP1HI7NJ3
KSWM5u7Jj5H3BLJfTWb9669hKJW9fSVwdS6RuVeLbfnwOhVj7SfT5Jkqei1Z6U9N
/xjNCx/7zfwh/8o4mUdAFrrENLbNVUf3+5LIPRDogvfVmkztQAJk9VlHA62eizeH
OGf9vLhqbxZBbaEXQ9lwIoEcP0y9zb/RaGuxKQw4UfWBvpZ2nqQOfT5+yJyjDC4H
w1m+enTkIx15qLjtQ7L9rWRBIval6Wh0Beahts8m1czKJ1VzJDvSBxVgCMLbcg38
ys53vOBZ/Sl5n30QIrNbjg6bZZNVygRLjP4sGR7S4A01XoElV3NktqE7Gi08zSEV
6hOjnC+9m/zcIH6U2OSiGL6Lg47DAWcriUTc/bkqFvkQdx8PAnPi6WS6cJed3+RA
f+p4dgrpdn98z02SC+LSsBkyKBd8OBbHqpPZt10/yE9oufbu0FM7ltcQS3oXDNpo
Acvmo42eSTMarYUIh+h/+qUqzkaUhIg+UmNbrIEaOoJ292aI7QrwGsYMXXM1sSOZ
XKSiDJt0BXc4+alMGcygZKDU2IGI2DoAPICD5KcJWSveU2qY91MLgRxDbwbtpo4K
RxjfHnttKzrUN4gtAM7ym2Fs4UqOvCqOzT7Dm+pOjOTjXOp9/F7wqAuHZzojiep3
4kbnaU6m89NGeHCHKaY3Rem2m6MeuYOCZzeyvdwuvI+EP+nPmy+hYZz+JERh51s+
Ygvbapv/M7AeRBXX1OnnLMbpyd1eUpMWeBwknCFqia31fym+UR/DLCw6o74g482O
xhSU6s3pAQp6C/80T90N/vKU78PPznJmCybCeFZRQkvxe8Sg+mNacR4DVhZXpfCl
9ark4T+4IlYNlDSL7OATjUpkjWGv55h09RxtwJxWKyuQ8bNTDT8JEx5QmMh83IzG
xSecF912sDgv6klC0oD8VSlcsbiIkxtbRGWqNNil7gvJ7c3lWMyCQq5uEuJd9GMd
vQ2EM2ojHnGVWBsxoVISUKZZIfiVYYfY/DIxoRXTolBTUERKw3Ew7rEIHXTaN2bg
`protect END_PROTECTED

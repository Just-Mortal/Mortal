`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWo4CTrE68dMVJ4q7JbFc27syxfQEa0USXbCAJ883e89+cdbM5j9C9tuoX+eCXNe
q43LTGHG4EDwf/2hsVI7vcU1pVqvEFPVHj+6DCs6FLU3ewZ1stpZZ5ZDBqNV/aN4
sMZkZsAfj5GB8UmgbKAd9FIp13SPesaPMqXRH58z0J4y9KwRsehl8VinOdYMJUih
B2Z5UcP/Dew26Der9veelYI18EkQ1hH6QqLW+X6jMLBGa74eve5dZwcnh7Pj+28H
0Zqu3xVF93Ee2UIkOlm64GI2n0RctUlOqlIQQpD3bAaVC0K8JDJM4h3mK9KjsqR5
AGMk8IPzdJjXf53PxilK5B9AVfzeZ/JDhas5Qy8anmAJ7tBJRNDvrEhEGOibytX5
f5ArF5YjUgd8TXejkpixSWbEV2GFlA1BVC8ry9QS0UPEBx2RbJjd0OIHeaCRg3by
6Fi3gG1MkXr+iy7LE6TsVtyo1VlSM3kgRCDMQSG3mKCA+460020DLZy87r8EgY22
MQzGKZDjDe4rCEQlQC5gqiRmiWHX4zvRw1+nmmxLY5EjmZB4XR0z3yW9BE7jiDjF
6B1nLFEYonbo2UOggl2+VLcrbkP/NpgZUy/s3RgXK0dVsCLvvojwA/hTHqjpuEPy
NPjiFS8uPUuXpYYFtLUnkryGoOxbxmdPaRwKCSYvzSdL8+E/Cf3SbBlBvgu3jvUC
LHgag1hII8CsBpn9fHNqTc4rFFtZvAaMg/VQx1GJIV6dwXmgCABRdK7UWEjIxDnj
siL4CqT6xOe6eScnPt6e0V66CEmSzlrwf5Wuev+ehLgPgqigKjbstDE2aVsBz0Dx
EIaM66XT0CdowzClPUmpRaXkvgNTGVFPkI4+8YXF+gRni34T1pxZMudTqV55Gd9A
Jo3dbUJNXpy9Z1LFvNyqcbG3AmeUoavdvBvYDCamn7fp6TnNA+HORmjWa9etWUSO
xxXDEtw7MdKiFwDdPOY/bNsX/D8rwJGWMSo1a0i17xp4X54+jgbZAX2L1Fuf0upa
fXc0fPrhhipotCxZYGE/DrsgozV7UH3lpcpHHC8OVTU=
`protect END_PROTECTED

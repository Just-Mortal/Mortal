`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDmTg6EbcSYALqytZ9evl38HgH6vao2fKSMgtHe6TbULUwz2cvl0dRGkFYFCRtAR
a+3kaFEnuZYGgM5Zk0hKnQZV8veOFi+cnVz/dps+Gcx/JhDzk0rIVg150DRuV3Vu
mhkrVufwz3+7gWo/sM3OWuoilbOjm4Rwshi4ZN+Tqci5xM7zqsU79Y+0VO7qsnbt
Vshp+u4Ax75QRwKurgmkbxP2xh5QYdj/gl8YXW/pp8GQGdGxern6A4k/EYQNR49j
V0ynPLHUUHddNnkVPGEuRZCbSiuHDZZP3Ypc5dF59mr2VMxP5V1YS9D1amOg4Kqh
2IawmcjMgYKyd0KA0pQwxzis/tS+Qwd7V093b1+fcnxAKGYtVCcilHDO8Zs+7OQ9
tJt5NvV18SSLYfg6OAnJ2RXkWUG0eNLzcemW3PdHwBptihBZBGW8z5AdrSYEv/l+
V9LL9zS+vxb/z9Z3UIRUl9NWG42b4AyR0LdW/c0/aIjL6FFT/IAuZP/YCfwOHDzw
pDxM2FqjJP0q11//1CIgNQEaTTXmqP/6/IAbdW37YMwhah3xRiJBH05w+SpVv2xc
levvgLTGxrrghEyi6V00BEffSOwyHezs8kyeBS2DmNa907qR2ztrW8+7mzpLAyPg
bnm/sbHE8ZPqPtqQZa0hbldOkN5ZSGq0NYUiLte7YvljCcz7F9MI66+LG3veBtdX
O74D8GgHyxxrYuCLxzFgKgyWZnP70JSV0AW+5mLWuzHTgfZPioLz1BGd4uR96uU2
1yDPCVW00Y371mxY2Sdwq9Efb/Wd4qQgVa3EnMCa38rC1VbwQwHJ79jXTLaK6EAn
z7SHATLpsfAwokiVkEdDFA==
`protect END_PROTECTED

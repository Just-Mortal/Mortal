`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BDfM4hp7XqOajPcjBvhAqXcNmWegK1ONjZYlcH+yzJmaaXgNatb5QxykW6LylUzF
e3KMy9dgT/Fk2NR3SM8ivLFRER2pLnYNi/n3eKrnEwJMaJphW+6qSt4ulov0R4MO
tNAAjcotS6Lm2JhhdvlEMmJ1q5NRRQbropo5uX53uBAtEg9Gr6VsDmY8FKomHGrM
Ayxm86KQj7GDhr7V6dtmysnGSwSgUHe7WHXiHoEvKQJJjI1cAdAStE0CyOFF83c9
2UP0KiF5vYSXzlqhYr73Jd4R4Xed5Kq1bjy7lG3NsdE8gfLFxPaFRjdvjDYWIgW+
YhHA86+Fyl5SlwN/LhqeNv+HISPyfh8OSGTLR2mmLeWL7bgWrrhZgOoTbgKvrb/U
SIZJ73rlQAZDazcFBWznyZhYH8PmaD5DeMMFHY5bTy0kR5WpRRwi+iqQttc+zLD6
GGqtQWHlji3I5rHmR+2s5IxkD1BERcf+ZoLjHIH2spQloB/ORvF7JVKJQySzXjaS
r5zn2MdqycRwZwryR6YBA9OY0vu8l62l/d0KAhHsjvZTOXz8equsZU5t9CPeldju
vasvogUBdUdNO6gPcU83AdA6pbApM7kmo0Qji9Z5nq4sU9Pwqzy5z3G6c18c98rF
z1GTt66PD8vKcHm5ze+Zyv3Uyunp2WLZCzh3Ym0suI6WzcWp97Vz5uJik1eTUxK4
hGjb9ZAbz4osed3HgRu8PqTxi9AdF1drGvPVEwZq78MJX/qC7XqPEig/LFQrVloo
pSI4oVF5S0/iFq0H1WoTqPImE5mTCzAHImrf9dIoVIR3tBTIwUzhoY2TaMZWK1zn
RQD28tS15O/JFU+LisbDs1ASPwBtpIS0vc8b4XRht8Eo6kGxsEFCNAEfmxOAavvc
1wDMKyp/NjcySDtOPwwXfaYQ3rbpL1NLQbBSyc3KwFKHC9CebdhKW5CKfrUw3xSR
fEm/o3UPdksuU3kWuNTLbiBK7d6A/XYxhqPL5EnrqRG3DndiOH7hx9CL7/nOaSCo
QfgdNK8j/+MAven5jOcvyGbfkJZTii1tYJAHLNX4/IIF0vu5WfEu91Xbun9qEZ2D
nAIXzgTkmtBulTF+gPkIu3x4GYzOlQPHaz312vQnUJ6FxRVeRdlvQ/2irarTaO2f
Knym171nFA/gNyknSgS/Czo43wGYG1NfImyM3HMVEDQ+hv2sL7wFYktw1TfFfUHJ
bIiGy55vn6KnJ55jsZCrXFcvau3+EOQ5Eyy+G1xJL2LT9Gj8RXaJKr8sMX7+mzj9
9KnZoNH77ZzTUhZSibGkC28U7n3sHf8lRe5Vi4onL1bOePRQShLGehzfWczyHyC7
i89PXPsbuymneD1EfkrPk6pxizuzjfOsUqVSeaWOZsY89D9Z7BNCXmhhAIcH8aBE
1JhTlx2fKMQ1XKGXvSzJclsM8s+u7+1PWRqyNAKjEXP+EahrgsFUZH5HDTsp2PbJ
xUY1ElDknbCNtwKpR9WqmXIg/BkMvSIUI05AtGs3UvqdydegI4kRRugxMIFrSYmS
sDWBdsv5lrX0MpGv2YIjxvhni722QaGiZf4togoUtwL3lOzAgdfizS4mjGVDr6mi
Ej6y+QtE+hsfqu3GOOW2MfGRpu2Ze0+Ra9cW+p/aezMZhfCPkoaI+/QQbBG1dwC1
43i0+uaPL02CCF4i0+EAl8zKv9TWAx736qtujPuVnm8Uboqs8Jmy+yf0/124Ck+V
Oyj/zs8vP3BqXsxPRN6dRqsX5O07QNNWVYGf9skMf3s/vHAQO/CwyPNLDmFlXeHL
0+u/q4/ehHO3veEUxnysr5AL6CxEQQRB5/UbMBnG0oCQ+K0gIuFXiQnHdzisc6il
+Cd5Ny94FhvvBw/TMZ9Bo5kW9tg6mX6IUor0p3LYE9TfGdADE4bKczCBbtwASirw
mWBncUNqxWAmlOv1P6aJ+iaM16L+v/MtzyVkZ64O6MVPtJ6C/rQ4jdLNsjDS2LRW
/0VRE1TEom9rpILDBprX8D6WOW4hc9OEN2/8B3m63hEdDVIQbRftjVy1drvpCcU7
hmILHADbb3NKVLDAwcYCMAfftDWcCqBgMjTeRhBEFOK2Y4nH0yUQedTwF+VWMeqE
MHUXrl7+ku1yOukPe/W4dIUc4nDI3pUhFgLrxWgwKCEfX7FqnWQJrOwJRNFP505O
JqionnrFCUXXzYhM9gsDDCoeLaI2CzUrlY2mEz18gLA93WEtaSoElHwPJQJ3vXbC
K/K/RlljHp4+eMjKBiWYCD8M2Y89eLYArjDPff6ej/HEgdM+8s6kdpsV6TfajrEG
LwSliE/ooLXccl6HnpqDbCRBZCySANhmUcvNb7fl3zM0Yyg+zvzJ67TWmwn3Wp0+
lKHbLjj7ShzfwjPn+1ahOKV47JzFVG3KbSmcObOIxtW0VgqpmIgp3Cr9vocMnp5V
6z+tzJ0uDbJU74nb43uNu4ZxZ6iedWmuMRUmtaRazdHcss8UIOZIZghtfR2d504C
h9ZuAvMXuolwYyqHeFllaRYkiicenLsJQWKEIAaOx2iugCw2Jl+rQ/RjLnvPA917
t/AJ049FAOMjXl37PRBJUclZqkm/zWBR+n6mpKiWjc1P/CTsa+qg6gE1Ob+c0olt
TqKr40u8bcyyYqO/DKxorsGVDbsraK6V9On9vpYUppvbjc+xxlsgvwSFFxOSZXFI
519nagWXy2ujhmnnS0QDLIN60umzwbGK7FBMCnVmeCIlmuaVgIoggO0vxmOETfyx
RKprteNpGqg+CpSWK96dkOnjTri7HhqfkLB3aFy1GQk1RncnVj97CBjQ1ENQXazv
Pdk64fVExM0xJEozlOzViTfAbegquinFzIZzDbqfQ72sbUx0LHyqPdfwkdRqe1c/
4ML4gwbxlg7peOSD+ZiT2SAh9bSI0/ls1y80M7r2Tts+CmXbp79fmVzfnweaQlCp
7bgvDDDCHM4C3r1k9PjjxSYR+Au6jcjYPn/G5ffQv727sj07rsuPptzsaZbr65I1
eraNmNDPmUlOkE2JTOOapQSkKxt8TQ/cVc3/LTkEv5d5u2Q6EnhLWkHVB3eq6u6M
YpCSyt3Xlm1KUa++PYdzmGJu9zh/5MGgs5C6NgCORlyXMKl1TqEyZYWIbFR5XLaL
GdrFlPuixFxnEwbk0KPqqgQHR3hgNbaDsX7Zcxbx6xGT964SQDI9yqfBCSiJLKmy
F8oXwaFu4XbxsLwgULeDOygZlnPxBSYUgra3JD6wwfIGWyH08lYimbc/dfzJ4ILq
e6IO4Reriku/g6FQuykgMxuC8O9DG8TxeJNLb5hoBmstSK07lSJPWD/jWvTAdjAU
vsVTOxW9ZKKFuNSATheS3K8qEwUuYNrNYxKlBQ7qwJIKWAeAkt8TWgeyGcrbyHt3
Z2b4xes9I5crw2GRiQYhli99PYMHv2oZQRymAgRTL948DigAVZfZ5SckgN1rq9Mz
GLGFgfB6CRETXnqp13IKr2o4YEEiLg0UPrb3l0xJovLrwgEj1GIMF9eUHwkUL2hD
nqx3OuSPp4QjUPFX+MQFWc8SBruhjDjCtBr68DQKYP+VYXOrFbaMDW9dNfUupWFz
W0EWuYsPP++bzECZYgaMjEWnqN1O3/v7XnP3BoTplLgla+QiW526gHlWjViMuQFF
MmqfqvtMiO9iCk1dVE6zZA+wDs8UyjkSGkKm5kNy0B150T4Hy6gF/Pb92MIbJuo8
+IeXXsXLf/TgZbi50QkXWbEiTiPqhfDLudxljp7KQlZkrugBeSrMS03NbDAy9wG5
eY6x5tM88Oq9UY/MU2yoslANYeVNcm6MFxJnVbbSdpx3bArU7IGVqsuWcfIEw/st
Gohaf4lUUqc1RpG4dSQ2tDvvb+ziHUwKkhO/Olej7eeT1K5w++h8N+vW627E87kU
8zrgs8Nv6zaLXv7jUYQG87TPq2UAJLNUzavNwg4gykpoLmfljngnNi+cPHj/Ucmc
RDw4SpsWxRUynozgpZYVxtWWmTWI6eZNkcO2LJk4Rhk/nyM1Iv6OmrROyZqRlDXj
X07LNMpfFc04gYldxth7eGKOUUZZQJASUlXBaf8lG3ETI0ubZGZZMYECSiberMsA
1tl/7arXDp1j5qf/xkpD3PMbXbr/Gf+urXCiM8UKkNEPcYzL7D83v2U6g2/U7CMs
ohqPAuEoLSpI9KtWabCPXaUaKrfmKC/mXl+b+NyprSpqihmv/h+51W1CtGCd4Gkw
SzHPuAlwBCSKdfidCZ7hcxe7lpOD+9Zq6UVCjXiFi+s0qAyA8HoPjPnYpnhHhBWk
lVOmaMTK1E/JNRshdUwc/O39D/7Hq0m8ozoq9vsBv+TSG2Mw9O8pKaharFP3lMds
CZm4grY33CX1vJywdNEfus7YbBT+sfNilchcl0WnDhM+EWhsEwtdh6uhcauE0+7f
HTW/qynSJjBBXhtC02F8hiA/E+p5EMqXuGFHDp0jzQr332BS8wB5Ga7+3BJgA9dB
RtLpnm0P3BfwH5RzIhvdC1iYc/ThTRYvHG0WhTrGwsQib/WQ/NitceZqKHvBNLcy
2K6nLl7wXr6+IhVdY494Q90RKJFGrGdSZoEaO99upzvB45oPAujqZYK/dnBu9vTc
S+H1haNl1HtalHank+oZF+JkUgqy+X40712vh8QWlvUuhdjbHgJmi+jFpyJv0JWz
jueEqCZCtUiEkghXldDOS83x8pL1iv6otSiZS8lZhguOhqAM0hJ7X4NfMZ+KCoVP
tWU6UlBkzJxZfEjxv4/KEIYwzndo4QsVE6J0wSg0AxCCIYdg6yKlW5QyhqqlWerh
caSHOOGF8sDXNYoOcDsJtSjiwXrQ2tYLFMQCz7Y3UUGTIdXPS2o+B215T6xbvfQc
2Ck6ZiDOdsqsoWYtXECso99vjr+fE9/x+UurZiuN5QfNLSN13lq5LNd+F0e17yPF
HjfT8PqTZ6FffKG+dBf4LVweSg9yGUdvwXuGkDhI3LPF9w/I0cR2utWJJdblcUIC
0o6iuiJyiEFhJSw17xxD5ifyJsF2FZyzbWXEZdLE+VXVUw6P7JHGqEu0n+zCmbLa
5ptmGPmVZ2hAPg+RHRmIKaDoHzyXM8UsWhIOI2g1vKqnHqxsUdHsCl4cpTWp8puY
6Y6NnXs6ZcXjPLNh2L5Rz0S1yNi+mEW8dA610uwMHR8tJ3OBz0rOaMxTqdys0KHp
kQrfxhmBiCRO8O5cqE9a9NHqFx5HkGsu6poxwM3Q55hCIWnQGhJdNFSbpGb4gqhv
vQ8HOgPm5zREDVrP9w/cc2G9Uw8auE2GY9lXNIKty1197gJcx9Ri+flYbldD4J/E
5RtkGIKZsv/yqEj1PrVt6GL2xrC3zUwrsZ6TWGKYIdEnI8uWbp2HlWLETk5x4zeb
+GlhruE1WuC6kNfe0DOvk01puZhfdo/ss507wSHRKth7cwYMmITOIsjOtivnm/iZ
6I/jlu3ob966fEGlipovLTm35HS/kWXs04pfexTC1mbHh+YCVRhxFFPJZIzVAvg1
kZqWL1T+zD3YOSecXXDIqn6lFmgJkKGZpLLpFFNm3uWj7Q7Pheg+vMIIJtJPOXHu
LS1zc7z1g05MYyTYRyF09cwJuYCBLXrAn+x9yck03fPOnwrlgESLxL3xA6sfqW3v
0Uz1qAdK5eGIkhynuvJdzXCKEbr6s4crtVKBwflfLom+UX6EHfghcq1OSqqnOSQV
T+aWQtYgnVWvAavQpMWfNXQ0xG9QHN+S+0+JK74iJRv+ieJTXklRR4Slfkez+9QL
7VNGcSJ+NZk6Gm5gN4Y1FLlpTTlJ1YtAWSjHP7Nwm76Qt4+W20pItaKTdZuE9BD2
vkOBubgCD5+M7aS0Xegusqc8iXchflS41lxOaquvcYm+mzWd8IdIoQcWgjhVrM/U
QLbIrDVH+A7fcX7LfykXGgPQgNTWYmXofdYcL3/ZeH3kIQzXMiwPIoLpR26Eke/h
CaZ8/OwuZZdHDeks3Qqakk7RQkjcxzNqYXGECWxZJT14IjaccLnlxekIq68TOJPn
Cy1rwzhYmZQlFYWDw/ld/htNFLzuQLbInLeFdku4inyyoTlnKt341JAyyhJ/82jp
PdzVQx6APlCbzEI0nDWb6f3+oEziEiOuCpopu2OK7MYtjw6r1QvN38tnzyxQH+/j
AAGiCugQTSFsfFssC/nVCZHTAi/oSGZOsVYe920DmlNjfoj1ktZikrAXiDkT4nkF
MQwHi6PBHPjX1FTojX99RlkvqFsL+cBACEZf9knHXG9jGvg/dfg3KJHeilyffK7N
M1RHWhCh+K+3JRn3IUDZArQBQ5VwY5JbkHdCAGmQkAeUasJlxD2YTv/q63gPXrVN
BO6FOlOSHzShOpRHnrAaIOr+XZgLBhlNQ3Ve+8clzmXMr07sAajQliBuRwyAX74n
LkTh+TRIRa5faRavIr2JIlg3aYa39eTrAQ/g04L56a3z9g5JNpZyyI1VAc0TzTSb
yqwLZW2cdLBEry8WnNiOjQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Z36XE/ouxVWWGF3e0oNo0uR52OThQPVU7QLrNkZxzG73ckGuXmCLkJgrYaT0KtF
vQ6ohlBG7ceSAZQjEn8xbvrszTheE+kMArpc3UC+HXRouzLcGrCG51fEY+XptQU5
rTlmR6aCj/tPsoCphDjXncEuY+sAidvUkrhaamvty4T0vJSgwjxBaUg0YOsDAKd7
W0WjGZilQ5k5zNSVSSETxK3ZFdSNRxmR74H8Axq7F6GOFJDbp0vO2KbK7+h4E1Q6
KrY/oJ9sG6AVBfiw+QnkPUuQm1DKf3lVtYF67gZzigPGGCXX4VkBEj48ylWIAOQB
nRe1SYuqFv//rO6NxJV0Cnw96VnBkOBhl6+bjAFzf9d8i3iXOIKarKby01KHFd74
`protect END_PROTECTED

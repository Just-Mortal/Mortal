`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0tyxjXvyPlYT8b+keX1wOR7FsZiJ5/ICO7rqneKS1IWkyxL2EfZcwbKpiO4cxita
0UjSU0qd/5ZNOiAdHpNwxe3lsztSNnAD365bzkZi1HE9bnOVc9RFE6MR7AoRIf8h
zf/j7c5lUmdVAQ92ZKmvCD3YB3Fs4BzwOEce+MM8LC1fw5DgKO3mXnsxTfcFGbRH
BIoFNPEBlHWe7UmsILWH1gzCNsE764FMhR+6Z+EUtBD507tzWC6dlaLgC1eOE8ML
mFKzx+pxqVu5LqowToM5CZdLYY4gv6m7wgDiOU9Fn1gE8UqP+VDV6c+H0dqvbOji
GbNVGnbCmWt3b/jBz5mHjsE82loNzCBwJTNlnsBz+7ipmVz9JToHcbRmL6scFR4x
fKhQwbAhLd8O/bTwW05zpQxnZWuU/+tMdcwv7q1e02LFI8RadAeqx7vXkXGuUAvj
Xmp8H401Wn0WUUMMDG3kw7hMC0snVvfwWZ/Q2iinGdiG43H75J5IVEAc5zbdca8X
BLcfaYBSXabxmybRGthFn68uKctKET91WdfVsalsBpdUeCG1k4UIR+6jYYGj5jST
+cF+Oiw9n9d2X+Z8sVvq8jcF1pmV55r6RQkljXmuxJN5eLjp0s6Qxwq1PM7WICe1
E6c2yUO7E76hlVeL8EAiYr8ba4lHCTrgbGi2N0Jy+GZnWH8QogzCKJmBB4gyyLbe
tdHCdmc2Alw/1lenRQLlgbunKmxPl5dLQyXVE7IWvmZ/RHTnBs7MkQybtfHryVfY
uFw2tpD0nviFcNY6liDnqn/pRUnYB1KyCEtW5Ft9EVyN+35PpyUQ81pCZ8bn2Js/
YUBuR7DNacjg1boAe/mlbPeuzzrohIaP5FKKAid//XxEmg4K/hgsFYCvUYNQgCOw
MIJe0K9yY090gt35Djk5J8mBgqy9XY5TIoylpKfH8UWOHRNonwNL8N1rJhMI6Cwh
I4gkwIk37satB2K7TUyhFv0XO0l0r7QopW6nmN8jxYmm1XwiuFH7ml9V27bGYBt+
WfHgPZyOR9vbtI9zDBlAWKHoUxMtZhaXmMQ0Mu7chPH4+3CaZNoLrq4JJ5DqwgCd
p2q51r+xa6l9CYMooxFG/tu7Igdb9WGpkwMi7lJq4gRoG4T8ukiIFOqgn5n5AsnA
V8TkC+kaNn9KAqz5e0eC1WCNbQUhTzzUwtMFgsoYs115O4WJfBTo7jwWLq1/GLjm
+hLI28NVYnlaobKbsZNgCS50OMKlDjlGgl7dBdhkk4EbwlcXMWSnZxWdjcz6LzkB
0LvY6nmjRJqA1ToJ5qDfpWzvR+VdISV433mJjjfeyye62JN3C+m5Txf2OFqWapin
1nbqFFNXdz+i+33YnxiG6n55rnIRHgboYIrY5cL+TcMnYLF9zeK6lm0xVkRFbD5j
y8Xkn1UZ8f1Vfhuaib/4RH0GGyV/AGsQ5DG8U/iOr5UA8hiH5Oz/SmRkl+pE66u3
RqW2fvFdiuDNlF7pY9dCVUqO57xR/aqmfZXAg2b14lWNmR65QE9wg6pQyTwvmWRw
UmcoYyxPrHZ4IxpgejPnWY0NsBlMQXI2OyyJXOiaTBmSiZ9FPjueFgHeB8dwpnQs
gzU5CMnbHvDDO/OJzccpdLPEpSHE4Rqeya+US4Y94RwPzh7qzq5iTgJW6fk+1pwq
0ZbBijHy6aEXq0sIbWCNk7ry7mK5Um3wzq+X3xW7eLwf/Dz3LWuy/8DQT6HyaUX6
NUvDGfULJo4VJBOPBNPa/Hy4Yf7AggDoZN0agUO2RGOB3qHpJLZbTmZPBoROS07/
bPMmVDbusSyVteLhBZ7MyuHOBzymZBzM/z53wFXq51vyYsh3aUMB0smxzCOJYkyR
/fiQWK9MBuA7KmfNJhpclGa4F+n9pE6v0ocntc2JKEzD8i62Ok6XqOupQ9UcpfN2
lxniBIIvC7duPB6lqXTzKGIxBuJCGvxRwkJunYLyw8caVzkSbTZI2NLxMqmcKqTA
YnXcdUE5HyufE2lrNyVIaXQbdJHPJpkl1lr9KLHHU8SV4rKFYDbCZqGJlP2GSXR7
qYbVVKtJzPA/cfsZBGYYL1RYpHP0AKBnIoylZQxe3dCqaPiuwEh5yvrFjLK3j8SF
0J1GmWTEhiH6cB1lPrLxYRI6qT/Ab1eVm533dg54zCuL4pcuset8dDN24+m+Iz/S
iY0c8GHkS4fr0S17OcGrQ01673VtGhZBSwha13eqBQHRy5THqYedIG7KE/Is66CN
QzGd5u4RLCYTy+n9NC9g7Xcp/nb1dW4fOvwMTN4WMzA13EOMfD069f6FPCCqVtfp
YMNOplXEe5uu8GpOW0bLwaNTPpC7lj32DOCqKjdALdWK/biNCEnLTRZRD5lZ1uOl
ECMayEp/A0/iuR3ZRfNK1C6HIB+djRWQyE4M+8XIadgfxee/WrBJ3Q/ECDMe5A7Q
TAu96mW4GtpC/qG0WpWxP0qkKdP52zd9RAKTZt77Ck5j3hrfflg6sfqMh0DTKgXF
NoQAfKnhNpGX3cA67vTKRAePzWJW90J+GKQvaibNMLfS5J982q7INBR2KMxwMOmV
AR7eFKueGzxfKUE0SxfsQ8JV2VHBmSj363/t9BEl/gmNbNYJAcLGaEYj3viFagsL
Q3kXKdB5KquK/o/0vV8C8WIa1lhdEgFKBIJcCFKnyV+WF+s2UM8qUFgh9OF9QfL3
VbFB8WJe7tZOfB4zDiHcRd7j9koahEUCmTyytqCuyQSLdcF8AYAOHqSgZhUtDy0T
sJLdMWjZAJ/a4grEpp3l8HKy1gzumIfA82ROmtyl7Nm031QWdhaOW42818I7vQVx
JafiQKhdqpUjJO7OxlyF0JQeHMQqz0h/UdWj+eGF1H2VK3UB+bhj+w6Ztj20JWEP
7AroAPpXs/yBeBUFE9KGLnFaOOC6iKlLDD6knxlzGUsP6ouy4qkkZ43LI7uxF7T3
/GR1aDT3g1DiDOIK9YPODrZHOCLA+6Sz+d88cR0EHxb69zD18glyKLqWDXlNqxXp
yAyeadIIjcHW/CzpItO7+zfZrou2N9ID3DY/eO7rqO1xa3UrHQtxKBi8HyoZSGrc
T1GTPnEVEh/fQLeSMeKnyU9PuTUBESnt3+WHD7SDb+MZvHReVUFEvXzcZI+R8Jpt
+bWDVp0liWjlsBKTE8wv0wVkJFlKMB1P8+Z1Uz8087GY81w6atQIVG47wIKEVd0Z
EdFFpSXXfTX3JC5cDmSCqsCPom8LnMq0oXdw3lfOZhhHoPWHs1lidMqvJKYylV10
WDzcH9p552THz592NZiGBk0IiH5aFryRG6kk1Q09RAU3Amtw/g038y+Ka6a1y9gx
w/WaKH7XOzPeicrg3DR5mmbOFs6STrftSxCHEu6xNHCfObzGKHbN2+aZVS/sgbz8
d92TOneG7aF8JQDqwR1UMleDDzuZPRPGQ5hdF8Li4bnjzdGOAmCJpANiUMJe+bM/
bX//AtH2RYZUS/j40d1Z7DZ0k9I5X2klanr1TIs0ZlyAEkO6q8kiOXLB0/QnVa2+
C2iqcNr7Du065Psv89xQ3lKR4axKfEvUvdh7CTxBy1CxqTVOaYUomvKXmTO8nw17
hvtRdJ08WyhW+/dfIpFQM9+Yp2U2w2/nfmIi+g0CcYr1T/iAaFVUEjvfE05OFKyo
nPEJVcCFjRQQAXoKCPEx3Oi6AQKzsPnBW/XOr+7ATfqMq6IyFJrPjHQ414KyA5gE
b1MckWaAbmbkdwfEgj31AA/BNi7lsVEbfwuRakgX0fiAtXBUMNDM4iOKxkyyCikr
s10AU0mFAjaRW+2IKI9Dkt2TKcJLST3cK70q9qLGVd8hM+KCJOCHfQcLw6Pw47Xj
zqnVfJbnaMjqAC46phlMNa06Rgyh3meXXG1ZttaVFd4=
`protect END_PROTECTED

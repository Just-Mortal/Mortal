`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JwvrMwEODqz3vC2q83JQ1BAOs9dHbvPcFBJI8OEIEu3FbvhbyXGTQzrw0TeoD2i2
Q5YJzzKQt47lpmIHhjnYqrdRb2U1SPmPg7X501/Goh0vN9zJpMCzU5EgGheJplhn
Vya26Oid2EuuxNPPH5qbEgB8fiENomIlj+/SwYE0leB5v0p8wps3eTjnEemeIGzF
2jP8RB61dJ1QJLXTjQl3U9kbFZx/SA6UmXqUGGylEE5NGgwvvE8Kuedds6f6nS+P
lTYsCqtIxM7Ml671fDRN/FuYt5JnshE+Khy1014PvJBEq6Ucskw1vhbvqPNXlkoN
UwcPp8bYL57/7Khqg7nvSkT/bTXkaJKuL4Bh1U2AXDtWnxwOOZ3djXSTD3G6XUTk
IU7+dQax8yACn5nDiBb93jvvM0hh9mzvyfXhgO60I9tOJiSCHEa7fc2a33YHtgOQ
vvrqV979/Z7S3enguvJ7tZZAbf7yizmHvbA/9wQL5rCD7nUnK2uHtf6ThuY1KOPh
Pcoatrw723zVNqUR5u8EbfHd2xxaXjihcPkqVYfx95Zvzm1RECrXDJMM5O/90W1U
vCCm2juScj22ubsOm4Vze64hbytfmLga9+tolkteLbhvYZjxpymueX55nFCOZxqV
Ino0sImqS+c4DiJel3PgA6KTdaqwrBzXkbNNO2c+EgoG82+ccyAdEl8B2h3o63hz
Wc68uGXv8G1mwLrKwjSZulRBOBxUDVRO0+1RwRLUdluBQ4PRp9TlHicSh4yLRl8o
YgpvyqeFZLgNDoykDsTqr6q6EhzyBayKp+2g67syf9zd7L1ASjO7RgWGb52hhb1z
HC/jE7Rw/g7okk078qFn25PJFPY55BOpWKOW4uvOOvUJ0C7clLUIYSqdagpyF/xK
arXP4LZtYbS6n8C6kgf5UCnNDXxjOYBIoY4+09byTbfbtDcJ1d4N/919DwqauLI6
iVLC3agVYDEgBaev9xkl3oRlQw9O7/aAOxsHhfmukZfgYNdaxMi0EKQUqpTGHwgj
7BGo7pz+Ht5FyiDvUSjgnYvoyZg9iLskM+wJxHnA0uATiLHnECQEamtEy5hs8Did
dOiD8L1tPDGhh5KbWC9xfS1+n/lC8obiR7V6q76cIAgMLy9nOLA5mvfMVPvZaWyy
vG9KksDisBKB6SOCHW+XL5KBFTUYsDlJjaXTldM+X3B4+MSR44ahghC7AyAjoCVH
ALW6uuLe9ZXgXZztvl/CvNUgM3B2Fh3ArFozPzdtsv7aXFMAZy+A/U6xanS322m/
ppTwDKr7HS6fNPOZGeOlGAgSrv6O1ZR9rpourcQ31xq6xfUH/J6ZpxLws0SLzZju
NBl0XY3bMNicehQjT+SZE9q1MW2Lgp1xDt9Q73kS/7I6zi4JUyoxRbNyUArcr7/g
IdWD+HDQ0FW3GfX7RA+bdjj8jMUmi6Jy/voIBM7fMhmA1wbVdFd7e0RW5iIbT/+s
vNNQUGg4Xq1VhUa/5eXp7oMG7hYWmAX8n60+eIuvWXcuaA75IYgonXhjjFD2QmIB
JjOHv4JYB/Kkal/c0VtMLAKR4umglHSBqq5vKQHuw5/7DlCPG1rq5p3I24IKisOu
HlnZ9lgbzBcg0kjWEcbi6XRF5KnA4McGVlWy/qBu5TW7TSWU0b4HfE3Aj2oGEs6v
N3aFndNBHRve0XYWLOkgKeWyVP+L1bCDO73e7ZRAqYSt+P0hWvuzzXzmfbFGoj2y
KPN9X/qSNSA9BQIqPe1njheysGvTjYA74kwOl3+pykFMa/Us+LIHaBkdYz3NknCM
FyRC5GLF5P2JOClFEFRq+SZVITlbBxFrGWBuICNdP+cLM9u0tR6E0oOGoCwbrDfz
xxun+TAthPrD8PwBVOtk9w4LmFrqrGGPyBHhyjhZZseGQbISOqy8cX52EjyyR+9R
+FqOTjGQ7wYMia++J1yNwXprbe2+MoKMJbOdFIJ4Vqw5qtAx/5lCn3zDDxj/c5lT
qWqcjtfxVqQOR+0kZFd+9H3o0lS/tX3Eh2EdQfMy/XqZcP7WL6DqFjlDHHMNOy0m
n0FV0p678buDsHEh7zOM9YinU2bc6qYORrMUYyIepjbGc/5d3DlSvI7q7PVR7iHi
3rkpZL7f0dSdTmhqmkU6iScmRWXSkKd5XuAJJIv3SULmSZAh2FHgacaWD4mT7PrP
pE8uCCAVYwaYbFH4Fm8D9o5HDqOsTR/z0XHzZnHQNXfG5bddVQfy9Eotc4TfF50O
W7IlP1S5/yjqOdpTMAseDKx0B3i5V2NeElFjGtFF6NOnI/zbO5xUXbfuhlk/jWf/
Q0UgMctfpdlS5m0mpieRxmsLo5y273p9E75SZ+eSJ/0=
`protect END_PROTECTED

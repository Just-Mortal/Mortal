`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpvbWNuho6DjXnQReri5Dj2PDSs1RP2DD4iaj4bgsg5wHxzza4Ton7a1iCCUO0hy
poH0priyz2wolRt2fqHJrVNzSUzbJMbA1RGEzx4Jr2dr/ZP7OCtNA7a3tgdUGPGT
EfGzMPuO8RBmZElV/8DnxHtGavhvHxFLeGEmBu9GtyfAVUSFaaBVXKgWt2DU/io2
RtvNbcQZabJzTD0boqP4l7ohvK5gAf+KEtdrOor/q5jbdBCXtbAGFblR5djNSrr0
DJ4TEZwDsUnIrsnmKmEsHLEvG+JynVB5tWq8GLKbFty/tB+X94Dqd2iy/9tRxeBZ
6gBX0Qmwdjb+i8RDlqMILv6fNyi9JNuN+FLXBI5R8tlxMF4kb0y28u9FQid6tCZs
06ccTbjXOThZq5BYsOx6zLmOj0O9Vcty8NWWPor/EpGEV5FcFxU+kvdEQewd9h9e
nSRBT023jagfOQ5tO53iqFlOk27wQghHjNIF91xv88esqCggsd+BRovWU0SB/Esx
IkgxXcvQmWCp1L135DllkYz3AJlS2QIFMdb58BJvKEF+EvcJUOcOcyHJzU0DiXs/
GOFt/Xbc0FK05k59SW8eO1GZa0H1pGwkz5zKNbXXzQzFgoFt3FFxijngBEfEW/5p
Bp6aO772dZZZYtiVyrPevls7RPwG3hW3xGjHW8eHPCycB0wKAsv6kwR3rYm98fiA
crpDr4xpmSZWYzsECvD7BtNnqL9si6UAN9UMbk0+peIxadvWFwN6FUYzfcVofn7+
AbtgfnlvXcYs/feZnZRO8AN57NBPdMU0uRGNLCtegXhl9ud/WmdZNWUegaEP1gYm
XklXtu34UlNzxyv7CC6tsEGjlQ7iBxDSPVOtliVUukIfTzPrbFRmpSF1TGmn0BAb
xihHMRA4vcWOf7qkDp55ktjEHOAD4/xHrGMwYwTaZQVkHhBl4fWd8/UOnJizPbdR
0z6dl6jFZE0Ujz2ZS9jFYg==
`protect END_PROTECTED

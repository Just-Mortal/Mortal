`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OQ+aGi6g8xOXIShGHEn1YGlHZCShjHtzCMq3FkOLXvb0WS1uI4glq8vNd2ZaXctR
Yoj0NrNDn9SosBz+uBcuKy1VWXjQjS85YHvuOHz/91LjlUVIAoz2ubMtFBztKx1Q
KvpQUnyYBIfsZ8XCHu/tYFp7mn7myXj0elqpDlGCqsmDvXc+V3LeYyTslSRic5dO
XFXlxtMVqFn13L9JFqWfOzWk3OpGEghCGdqw5Il4TuRnQSIIfDeDYgQtwa1eju86
vw3NbjnFQMtvFjaOzNdsQwy5ZGHGmNJlzLOE/OzwxSkOD3IDmd26HWCFWGA7wofE
OfRbSiJ88HGf+eOLnKIgnrUNbKZctlOKEaaRDAMCTS+iISou9qHi1+XWNyWhFCL0
cSv+Z2lJnIx6XkUjjn3TB56O6TmspTaOH79c6auGKBWTRM5IUWQS/fY5p3xhTMAO
ZkFZV5EE48qcPCGa9ks1CJdBz5eNrrDXKXhSl6nSJ5cQqJONJuHIZAx8ttlqwzJu
0xC79kyK8KgdkrpADZ2Hie5gKXoy4HELmmqFrWjddPphulFjTLnPX35mbVmtUVH7
IQyxl+gfMftLvPfsPJRzlfP+wiPo6/C1sr1ptPf+wQOTIObZPl6J2HKoUoxqrLNm
RwZNDJyWtIMvHNIOx9avsAYEy7LUtfq8ONGGy4hT9lVIFBA/J4KjuvAasDx+xcSF
D4myRn8fKwFknbRC9SdsImkGms/EUsEkyFDbaB++qp6vYUBtSRIMmwg1aW1uHXJp
HYsjJwOz+x95UbH2J2VRSQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ePMvgxffXlkmlVJpfBTrQOJNN/zynmD3WQGUYqojYcmUXLYT/5RGGo8iMFLaAPDC
+tBMmJobwoHgqP6O1BTA6XkNitI7FxMQo99v07wIrrEgbFGkaX2yvstm5K+mASKs
BlLq+yKfgl5TJu0gQZYBBfnmBSd7yUsoHizuD1EpSSPqWHvcUtWN//nsPaf7M1S1
eemKE6m76kaDxEHrjJxzFsGYrX5+mtHVLKTUOa6XyZJf560Nj1qDIgmXUY9QNre4
4b4s9LT84tXJQISjQHRvXNovIn0p98dFCNQFCeIS7JtklSwWrG4RvuRW4vDP9Zm7
BbuJI0JRhghkEVVH8t8icAoI3sVoOcFby1zSeCJjAJZeKKoEK+GsMvqwQ6mnejjg
aUXOuvjYZ9xW4vDrAO9C1gF7iYm0aa6fYvS/KGuVNM4SYORsXyaUGBgQgIUbHC69
7KEuISPNMYFB49QAdvGANS5/oF4GMXW5CkjAP6IkQyBMC2Kc+wHLc+A+rBtekRuh
CBhBlvKgMHJLOPmT0Uo+ASwO3jIxmKxkx9J6SiRt+1Q3GJfm47YsoBwom1+0Bbwg
uG9DqG7bkk40F5Y7/hvHjk1jgah7G5rRi9aPgQYn0NyFCNDERwI6M14Bbl4Ay6iQ
qDl5orVpkzVUcoMBGg/xd90SVQXmyJKl4oHHgkcmTSuL+0IcYGcylqu84zPHAK1u
V0H/vUbeQ23OdhxQ4UsnahzwqQ3ZVRFqtVVq/hQfY5hlGswwHwi1tLFkhgW1u4KV
e71AeqDz2ktUMsONaeQHjzdDjsSh7gvbU/tz3fsdqkI=
`protect END_PROTECTED

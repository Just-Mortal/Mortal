`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GJb3GNWgpoAS+lcT0I32BZ+v9usTzESl9hj3SHamXpjHUFOPf3FiM8c9qvDwzcGL
ZZm2O2mC6xXlba4Huzyjwwn5zaWuQSsXqCsWCrx1tdAcrUNndcePdr0XKAQZftWO
YbiLwG6lSTMgdlWQrgcSSM5k030qdUENfUsWRiNnmbgTy/85dFQnDGXLlwvc+3rY
Vgpj93pbVVXoi4kJwpdAkSsAb4LG/o7Mn7PbayVs7ZNBHqh++FriaUbdH7T5UoEU
sCLJjk/kLI4cuP5rbnh/+jJ1EyWXR/rb44iWYeTYENUzehMbE/ManPnxe7UUKbjy
FCGxFbigtxoxpVs90009ZePZbikFqdz1keEAkyCqWVtwzQHNxwAEvGMNLELMvSxT
qWTVY8ilmJfcEljJgvgcaUk/G7f0s0595I97wtdIPUXOAc+X0DkbIMPZrgaKAU+X
AJF5lWnuqUzDQxHDcD+6oAQATgzuxFwV7iuYbigv7TKWX66dkluQRBYGxZSJlIL4
cBQj8BK7OEVCb0XUZ+Nd9Y8TKCAm5WlKvGYPQ/RviuvRiXGf/4hEHPXOVLt0xWcn
k6+ZBM68uhUqT5hLY4LF54Rm8t3N6g5n8J7rsiCFYkwgarOGpfE4ZRsM42edZnhE
ghStiZDxcKFbddHhZOU2SvRstc8DGKduwwdF92zKbAfbxJ5pCOYFtNlDeYlx5PZT
t/kx/eWYruZqnbwhAJgdc2Rjmv5JxRwFwpvFxJ38pX5ZeJ+Q8yNovLUKD/J8zoWk
XGMW5AzC93icvlQmWhpVDhqcqtPpC1VztU6fZIQGO6sWFoF8/8vRPDQ/EKm+Oa7R
zH/xiZ1Ao2C6qwP+gpyA3dLY/TCGPil+XfSVsV41rOe/i+iFXqL527TZmHs/8PS2
/q+vq6wZ8bqugz6o3VkmpcYLtYgX+zugQm4cfbS4Pd5MWJD0gcIdm5fexhIlNYcV
3KKMFvgu1EvZiJEaQaxpGID7ZxCakbiouirB6h58UuD9hKzFERkeO5ls8u8FIf8r
7aS53ByQOKccRM0TxI9h5Ta45rWMYLPOqUCKq2xX3n+RbD0uFqQElZnR0dCE+rQv
2LYQglU/w8jRj3CJglP9IuJBBc6tS7jVfKji+17NnTubLZPZD+ctmRvC4b2HVNb7
e+R/WC6iGvhBiAetxxgdXLPoqdNobwDy+BckOveP01oAb7eq7wVUQQxh1D6Hp4PK
tbnMTc29tch5CWruS7QdX8j8ZT7DfAyzwdDNCoH0hN/dwsvEsi5Ub1aLBqJQ2KZ6
yolANjMB5lD8OSNKfrSmut83i9OGRRlC+Hj/dXhiolTUoFEKzBZgi56XjpozrRk3
5/qHxzwuW/u8sKShh/SMuAZNsgwm6RHG2YWyqbpwYRmPBUHKNNZG4dJV46lDFTgP
GRbA7vU39DuTC5S2nII9/x/4krEHyZiDd0zO/Lt1lsYqu8rz7Pfnm4IoGuFLkxhs
3RazuyedCpNvP8JHjjsQScx2brsxpSsydfXn3bLsSCkYBo8XfxfncAiqdnpP8Zwd
Lf/Ep+FJoZv//vt5unL5dsvjlOvv0zHSFJc3kn+LBI4riED0awmzA+rVGqXu6eJd
730Y1IqBlo12nzB8oUB2S1LtIdPOiDX6gzCBFkwkdJnyP1aYC3asji8DxcBfoQb4
OfF5qcv5Gysvs8VOFScOOl2zptGJt5gHXuYOmV7PzERwDBHgUBg1nRhhqyAiyG4R
8emaY+CrusHe85DZHDfSLhWLCdJKviUYSV9INFVqQpGd71xPbTdRxujHMR664/2V
vjl9f0rkQGgdV2vD82mBGB/qKTAuPGjvQ/acMes4xQ/GTT5nOyzbKAfGlyadOWHE
YtZQRnq7/864lFD7gEUZL82OVdGUqJJ6Vrr+WLbY7gmRCgEx0OhyMHEDPT+OtbtC
GGRo5l1SyiKKhIQIIOnayLaXNg0nKXO8vo8JxEAZecfS6/2xAAQhkR7LZqdz+9jH
yZ96KtJHds9Xo6n9HAmVJnUPBFT91LXDq/DL+0ngzrQ/jpIeo5D6lCpvlTZfpvp5
FkZQ7F2F2qJNao1xTzKQA3K3temUxIQlDMzKLkOMAbKRsc7185D/4Z4geztvMvpv
N8fDEkuW0MqxdgF1Ad3qvsrwC5oe1y4XPQPIeg+cv+RKQjRm0HNMoO8Ry+m9sLnD
hv7UCwuUdDLaOGwomgvCJkDSK1MYEy4w35oDaMYxpRXoTql5EGRJ2hrm5gvF/oe/
zumDb7u/hsFKCM6x+byWgm9cLkn4ragx6PVXpyBM+l/ErN/tLmP0654iw+XRkWAz
TTgN08NlnhsGLd+jiWL5hcinZC8aYFtgstuwgwJrS9gRpgLF3Lwj0WijFtKjhutc
b0Vdm7wvtrWue4qzotYldoWggbqk8/j9gifsneVjM6INYu4pMWezFrlecCwHUM/n
5vykO+Hpg7RGrV/VqEgbnFdN18/Mp68e8YAQuC+1y+9k+FEqh9Kjn4kjwuxl3PsZ
Ye8NDe7EpfDukfE/sllCoP37uYgjXfI+HeneFFI0MRpf3Byw23TelIlfUFkU2BD8
nkB8Rk18SH5tX4NUlYSiQhdvjHMWvkdI6Jfu30SZeyiQoYaGbifPAYSV1Y2T3QTB
6CG495y6+w+mE2Eon7MdPL2g+0x4ac5FujI77qjhe3G6B4fFAYqZK/TPTuJxHmam
bNsUJNTI9DuTGr4JpMfUqbxQZk5XzsooobIwIph6cTFIynpegYMNvpM6ngw90KSH
4slOFlVfKMsl2YXDCfOi6LycXDnFl1vPrTSrGd26P9fUz5aQjyVXSNi4Uzk30BQN
vNjr9IzygkBQLx8J7cV1tnyWZtnid/Vq68Nr8XpGmQZtmF/swyWhwxWZhGx6peR0
OSiSLuitxe49V/rvXDn+isbNMC8/1rVPZmywtxs1OvmcA4T6/YLx+Hl7sdz17k3G
GxsRCQgXXelkuVlP91OPNmqtHv0RX1a+ldB9EdpuSLHxyIOIAtPmY8DV5Jv3MvNv
UQTGbVbi7LMsdfhnZ8gACskdDdc3b4J5VZ/MNKfeengwmTifZrpJBqUgbfzJGaS2
xYkGjqMTgKr5REy8YTgZ1q5rvcu1XPivUYM5BNh/XEO+A+7GHK2T5I+JIN5X5rFM
SW6YSVSjt24eVxBggqS0DufYh6e7R474CTstFicivGUcWLXKL8JxUe5WalCc5m9Z
cV3wdhf9gesWCn+tW3BNDiLiicKT3BYz4x0z6gnQ2SodBArEV8O4nEuVOhZAR0sQ
hq0ISil3unmX8dmjpRywTDTOrUXQglYrdrlz0vorNugxkGVuz4S8ubKQiOw9KRPZ
oGWziPApr/qESl2PQnimysNUif/9CULLKD4UV3mCEi/I4eTKcDF68GSlVT30UB9N
VjA7X3+O9VXKzF8s+TzoSrKOwPms/9FNjnoe/4a3JMYoynDdvLmxbpyl0QlX2C+1
krbTVm+bWtO19G3YyneBWuWO9RvzCQY9eQF6HGYpKmvvtNa/na4Zd+KKoEBwZPF1
0Dszf3+1EZ0JBJtGTVrDD0DPaFJY9u4+g7MPV4VJTXDvFMtg/D+XkScU4CFRSmk8
fIUinZc5s3LO2qz4fGlu9Twg4hN+s8qaw4cs53e13lYinw/sXfSeWZg2IMg15HPw
rZBEP+BJbrbxw4x0xVY37SeUowOGlxdOlGYRpDz77nhIPPEieEsYHTXgn8jw2vjt
YtXjpb6zjd6zS6cJjM4/jLe9IvhwVl37wpyL1G9KymdMMyY5lr51ywsfNgDB5K88
RTvQLZtaaAx45sTmKz28dYGWPfQQpepR4/i22DMMCgx58tZYIyHaMMySHQ5JwAhK
ajFqjDBTD+sSaAJq8SPOFh8t77XVOGEwpufwUdSGhIOc3glQmgx3Ia/NFLDdFcwd
tsrj+K3jG1bpNSROJ4VnngPnuGfsuzAJ3E68Xy9yQQzotWARyVolXJenTKnxRHV3
bfQGa3Y8djUVm1ugEFZS0NOdL2ZLjaBQ+zrGpbP9aDspP2qGrzimqR5GknubOQ4J
QPFhUfR34ZIsgSxr7b7sJkqblGJ/mxn+F3KPNuuxcFK4avAY+9Dxeg0Cl7BFGpFL
JMYYInPMMz4wrDLk2wWGv8UTTf2Vf3skkYO9kGBTwUDW8kdIxxf9P/dOq1UZAbgg
Ysa02ZZQyx2J+ZRYDVNYxiusaUUqNTsutCxONOT/FsxWvir9ssQbt02bj2/69LaQ
Yp4q8kczVg6fl3jtU4dU+DhaIpPCxrFZFJKnCspwxw1UC596i8HVuYii/SAPgRWa
HqUOzaK1SNr0TKcwlX3UJ6/vIfKmLRrdF9q8+VxclMyoQ375VVO89D6qpZa3FTKA
ZyqcuRjK/fawLgo8Aj6Ja5Lk/cU7bxYowIB3iyUjh01klkZlwVJ4zlTcwRw2IizQ
2NUI87R09os0zfYO8MqCB31k4QD29cEW5Z+NskOOiLJy+B0E9hKFfXyJlPUJ000H
CafnYwJx8oNxOCrXgo2pjYDoYoVosrLu8pv5qlhuWUsr3U85aP6KyDS2hBIy7FrM
lHaU2EURUSblXHmVF7ghh9Ihv5i35KkO5RoK5/MdfADBysjNAfbyrjC6RWeQaE5G
6YsBpCZOzBaYiUoOSSw1mm+TnsXrzZKNx/SrkfWWlo6QtCCFzgzBT6GZy8nN0Rz4
tQqFYdaIqN80GdKXHu+DH4IL3ekcWS87pIYJSQjvbgeL3iJgB+o8Js+ZtiHyMgXO
meo7aQ6ehRipehs74sBUfwUxPNBXJaKdhi53349Twgc4/WdmMBVKJNOiSXV7+Lbq
GG5d9Nf5n8YgtainmXswLjgBahCvBzNizz7Ytw7xUbBAwLknlMqyZqi1u1778CTj
TTDIudOko9kA3cx4gyeMU/HiVKbyHK+e2sYPlxnPq/ZYtdrC4gnNXRrkqfoxznky
Psg3WslJzWDsn4QAN++TwYJwRDRd+cSnDhKYKnyXHtN+JxBpo68uo1VNbQmS578A
GjRi6ZvRylQ/4H1o0bMBIIy6BGUGExz6uiIM72l0tLxAJwh4dX4vrx+mW00M/ye4
FxUC66ITHXYLfr+J4U5X5p72w4bYZ1+aGsd2M+Py8vGtiLabXNsDmOfMuP1nPyew
rkXzCIG+XFqvGVK4H+0PenOckL2HCat4lzvvCwamAMcxMt/QFQhMkrOitrS1Vgic
WEG4WoGKYKQei0UIuqiAaW0V4Vp59nCqmaHnjdCarz6f0Mf1MMFQBMXPkn2dhM4j
GshZLOyg3uWDMD3HUQVoX+ycWZJXuFKsFV7jgA8dBYQCHG+L0HDhB7XEIkUzX/mZ
AYEs+Axlf9c90NHX1fdcUrFgAVPAjbiWoTn41Rtc/6JbDEIVyJ/NvTYshAyXXaMJ
q+SiKRLEQXViVrgBmQ4pkEtz7hFDC3PaGg3qIPpSc6PviRYTc7Q8NLXRZT7L9tzZ
2ZSDLoyXk6sIspkg9RhGW3cTR5PL48zwpRH8jkVW4hpW/Ba9tNyGDJSo0+IGmXGS
qxmxuR8AK3rQDhMqIx/j8rb6JQTDKZgtv5Y8NCniCAftOt/no9KmhXnVehw3TEbS
Nejt+Q4L7jGb2w1bPAQ0SK7lEtsrG3VmUXLDFPCxXBzIDxhIRTA3ZKHyHw214SSN
0R9rZoqGi2dH7AzZo4DBDN/fJze3hIeCutH0PqqugGYcSAesur8v7EIibowC4t18
+1WsjRTHLNMjS5nrLMOy76Y2hnmsp7brWPYP2vp2zis801Moj3SM+REnoJizhL3x
ZBPL1HDn4/ZUIp1ciPG2uQyeSU1yPsCF4SdimCmfN+RtqHnI4UPJTROe88VhMJEe
ubDJnsiHYDB35rjPp7P5wU3cQ4dV0YuZMGppOgV5zE9xNPoZXyqEBWtwpcXF7ijz
yiRsW1pEBeQFRckPmBzBLZNXr1TAnM+ppshfBHD83NLwEUy9z8zDimLAgPaoi+Mm
cqWI0gLmMkGVhzxGAr36IaWvm0OS6y2z2R4QIMOgFVPsRpqSylQjztvuyDGDYI0a
rbFxI7g1QfrndKbx4QPx9tYgE2bonD0CWhiwbAmeE+S5vVRnS4UPRxud8yHbxyLv
3PILcU8zn80h/GWAUcqKJj5SXErHZeTuBkOTL7ls1TwbBzmrHvXMwzDN+ZynFvP8
eUQQ+Liov8idcvfs9gpGm3bFqUosIXZD0aRR6Je6YyG91gLUXmP0icBvC5VPGcK5
CWDwVxRsJd6VGAWjpP0AnbIfAkQRqrmLyf7isRuGIofVBr6bGQUXwxow0VJO/pDa
MoxTHBG2Vvn3CiaFzTeOxL7+on0GDCpFRURxGamdOrqbAHuXZsabHiIYgIZ4qxef
wKhFIAsnr29PG3akrvUdGFKxvLOVcEBhkPX/HgG+B3gxB7ipodRYft71IOsHQRZ8
0lrxvoqSVhG6D4PijMfAwb8J7rDezvraLaEzIS5kB3mSVCDSbjPfzeayoF2qDpU/
SXcYK3Cdd83rih09T46d5FX6DwCnfeP7sB1FdgE9oGO3GIQ0zuVKID1ii0NNLlUP
SREClpVSDeaaL6OF2khIsF4JbZpViJMhvvIgMYneCuadnM/fOg/GCQW1d9W6z4yu
jlmFDSpqjJ3J8I61Ne1Ox52OA2DovIJep8vI8GbJmr8CT8Ye3SPYp1evTGeG+bQf
zvO2D/Plf7DFK+oYXZ/CO69IdvnZMOHDGSUUGkHe1vB8scJx0lDRLWVpfoCLRxJk
ifR+7S23UgB7zsBrx7GSMUj9pZ76jk8uTWr67ql/0E2ayJynadNyMOUhUwKtzPMA
+S/dOaEYlpGQmt+8p/qh5jMt60Rro8iEz2ilyXvFqRd3vy/Do5XA3bRkLDsfz0/C
ansY4KGTDUZe8Q3tj+Yr1wliDI5rM7XPSKJ+8yDOAKBEJ+VZMucBF0M10spam5V3
UWxDl5YkmTxR0k5kfLZn0NkEYK0PQ83Gm1hYhswC1GJZ0GyoTaIxhUa2qh5gzkTa
HwO1sBqreVYoJjIW3LiW4AtHLcNzhHcl1XtkTrcG1pFszE+tPh8dddausIUrDr3K
p+uA7psHkaDdrDmpORByyuRLx0E9xBlhIljuhYSmB3ANC/SA7++fRHgr4XEOOXas
2ad8lbihIsUByjsPECAQlGHWW+nOvM8NLSz2E08WBOIVks4fEwX3VFIhS0+aS+S0
2+HUu+oCn2k5TbPrOJBIry+G6cNztK1yu26I/0aoj9a6MOK+fXf58U4UpfjR78OX
hOiHus7RMFl3T7xZuHIVwH3E5Zri1kArbQyCJ07pK/53919MoEIR4OIocmQqRRzu
5vdJ3Ro1LFothBB07n6/pTPK/FY03op+0L/o/AGnhrdWOrwzR1H2uYxYi+xntTFR
GIJNKDRa8rGEAembdHm7XEGojEkubSkCwNzZSC5UeYk5OWXFr5g98uVAaQrV6Xu8
TMqegCaMsAokFIYJ2iJdFFantYxw6JgUCstzoeRyCMnoPAQrIW4eDOp7ZIGUvCZL
GwxBP7bAK0uLSNB8kAFjnUjYLDw67zCokdVqRikuyHFvn4jDONtHew1zgrne97dg
SNOXlnpM2gJP1MzKnAhBtx1MvElZS9NWZdVyH9T4MdB/2xcz/FJlfkOI1b9Vb5lp
KmWFP7MI+JnR/3OfzCCwskFbFQk7FtAwXmX27X6ed+JL09OXtAfMiVxDoI110+Aa
Dj7hoZCOIOslEzyjlm963v4hR5V6F+ul7ok+51rBFkMnKukgAw+Pzgzz34SvYTCz
4lxPeJDU0RpPWel5eYaagseXMzYnsyWSsI6+0rn8Cc4b5IWDSZMvR1ZI2e64LGDs
QN39XCgcKnt7MsRkqNY6TASjKdF5iYoXrC8D2K5X3JYkgHOjDrBlEfgaK1vjvO8T
YrQM2V/SOYBMf7A0FrMKhg2HMLzKSl+4rSKZE0+Hm3jgTJizCYFi+anK0gqWOuGV
+ZnPE20qXLPgymYEuR+evTu1DBaC/tNIWcya9EVRbxFhRy6I17AS9vQHdl6w6vgT
phmQR/OiHQbx191s2fpzxsNtjXl+OKmKbZhPJatSYIB0PTuGWND0ZRcvQ/LPGSFy
njpb1KF/SRS8am8PYCoMheLW5+sdfICkC3o+8NNEuyCgJt6nIiRTzJvYq2d3UK/u
AY1OtoqezHUJyOqN63+V4sfGUOAO+dW5rnxI94vMw8Er7E+DQjYxCcv7E8Ua3jGV
aZ381ntcBHCibHtfUhVP3cjshXTdW8Tct4Hgvl4uvwJHLO5gKuX8ve3FjwU1nAjX
w3YRcdErVToXvKGo8irU9nWd29zZ9lDzuQP89eMa3e3pj0OVHBm75vdJrk8xa4pI
zJ/heGq7LzwmkR9VYW7sYAY5EI0UykOw+4h+OJuxkjhor93p+WJUMCCP3is6DddE
o6mwjNvZUZGc7d8HdtM2ijXRfoRNWTEC7T/1GaXmEnIWZo1C45wzR40RTwrSeipf
8+Z0Q6zJtEHpQi29m0kGTQ511PjyB5dixc123O4NFwYq1FpfvaEInNUrWqY54Uqb
mjkTpx7EYmpv5z9Sa20FyD5jhyt5f2S5aZ4oaQCvHvOBRrw902OlrAlsrMQurVzP
fV5rJ26hfeI9Yn11yAmt+SPptXpU34erAUsSLvrOb3wYFjEw3vqr1P3vofKeYyHz
cGvFFsILPLqAn26dgOND5ynm4JKaBwemg4+jf3CzR9oxJh7RT7WkB4HaMQIu9iTo
JgWs9e6wOOIPptwbQNv/cK2C6eXDC2oERuXTXYOc7i+Oi8l84OxBsgvnPWHVY2rH
IbR5isyjDxHU/1U3o5CTR/Ely+4y9mKgju9nbDCwwXdLfxoGC2vz1y7Xj608uGPm
KPuvy49DD7wH6QTctH+7eFCkjUHgFvPmEMQ0qbaaQTfkTMivaGjZXgRv+DZBfX2n
toAkS6lTwunxgQGwEYsP8sTgyPgbZpDRGglbzfFIDY3yDNv5dMnARze70UZGATct
A00iC9XlJonjAAARbF4v0Kv3xUPlTZKIwS2w7djyCf177gtxmKIVuISfUgWWVgeT
R+mKWgTttZ6Sg0DCEKUeUgLFXFKEhu6trK26HUtkArO9JFBzI+i1Vg083zJcC4oO
kcC1Ac6aWjim/xb+nJSNwke2HqByKOZk1fkMmhDDsogledY5lsrgDYS18p7VGLcd
bzbb2oJwRGqlrnPiV8aDm4KU7XagFf5mKK9c+93K3IqZVm2LZMX2c0gE07c6c7/b
8ZXzdNXPGSs0wLzeEOPRx4N4natgzP+ngLCcI60CF5SOl2mqSEu2ynlHDqbDm/tc
XW9om6/Jc9dKI8y24PDZhMr9Q4vYtOIS4tNPockrKg1cY7Ebl9wd1DWevxPweok8
5WPfDu032mqzERulo5D3XeH0U/1123uNtV21wZEqb27Z0e2RUEF8FtoDGukm5c8p
8Bn4/MOUI7Gvqkkpgy10KztwKKCN1JZOlW0EHSkRScyJlLbhJqk8zjx2zp67vLBv
aGxUsmcphSwbhS5gqh69KD1D72EEjPBoajst+vAQn9slsKSxfZg1Y4nJ7LBabT1N
QW7JXpoyHEZTFjarIftEhUPivx+HrJxGtkXHF3fqBNZyGjmTrfFXFlXJ8eRVJxMt
+wWJ7qwxsM9771Z7XjQxRW++k8k+VwFU1+7BdbnViub9Jd4ucMEPz4cCVjjskM4V
WTTAdLqX3okQs6qIfjMHG8ilhvKLlEzojFK0ufF+difGax6sRn5109U7B/be1OgG
5D3W8iv24gEoIP2VRn34KBQK6iyASE5LunVM6dUzLpoFKk58Dt/ZTdCexYHdk+lH
bPAB8oSI5eH6pyduJRSlGonvwlk9ea/0lxcS/KTy5LHDqJZVjliMuGPwlga94Iag
ozr9nPgzipv6cf/pviDtRx7iMvPLLU+Vy+cJj93DckOWS8aF2bWVOhVtl3yr4QZe
G/FIid8gd947UtCh59GjBTWanh+uL8Zv4wlVszK4YEqX8UVWFURDKSyaeWvhsbLL
axpCHf+Fq76rtHz13nyqp8C2ExwRaSKfM3GsqxHHdh34yCEnUpUVQmBFqnak4I+L
R/Wt4Lavk+hzX4m5RiaxZYOR+P/cBgfj8dip0KTEmwbECYEjDP3ttzJ4UPvkJyGk
19ewymoiwfeoUUNWyF3rpX0xYistMswtZZxxde/dC2sIchMhMHjzTkMOJZLRcdwG
vygNEWd0hlB/ICRaSaa811ZRv1BJT7AHxEp1AjIni5MGTGvFk3/7gf51fNgTFVb3
+xVbALBm8pv91ZYcPgNPpTmLkFZ9zi6rx8vYF/OzQuAmldpLpcsLojE3lb1/ix/M
+R7Bg+ZcdPQLIFHtdiJz5DKJAIOi7u7TeNc3l0Bf8sQwJJUEPXJAT69UB5CP7Bqd
CJlEl23zt58oORAxJAhDsjt5xrMuHX5tfVIfOHk4BfhlFMlPOo6Ub26OZHG8GJBB
4rOqCUxP6L4e2/fd//xjHxrG5pzbvJD9N9xiPwI8z6VMigjZROkH1/XjftJbSHr7
OcirHnfTo3sasotUI9qdsG/RgZaAwsnJj7EC6uBSjHasW6HDo0dDqyPTZvPitTxf
izcRQdA9TPWrxxqfikjaHCM3xwZBnQPKhcHitTsKE65wfMsK0R2b96RN7U0z6/iS
6oGqcFhGRs9VrHxEU+Y8FGwM2/ZjIilhjp1ldT4n2OtRoyIzA2XcGiJHkqv4Bwe0
XcllesyKRL5ulh39heHgg9Tidth9OMangWvQCSGNdcWLWrs3dHlcp8IdQPJNsVop
+KztotsNi57y1+Z5ZuKcUkCkil7eNGpFGhwiQKx+vtiilZuRBL6I3IqP3qr5MRy+
8Yx0SWUAaym+95cjpTEtVcaN4dSRKb/13PcsYpkm3jjNHQ4gJukUutwFmwqz36V2
YNQ1pWUNsqdN560l1wmSwJj170h83pPWa+e7SxECmTu39FABJkdiWm44WXrsQDWS
aA39pfIohDlNokC9+dztJCDAeWAC75cCv+Z9InzOKBX/Aw2lHjtK68bKMnLLKI33
soZfDqt57VuYeu5qCwdcZyoz6MVkLTy3o5MayU1Eld8T3oibVTLXwZINq5wYOnEN
q3HqCPqVESunL2dw5uCnlMJ74ifEfSiqJhH3xg35gH+uJ8Oo9mXgSWt33mMxSZga
KcSToYXKrZEpr57fT/v2ICAeIAHvVuY6kgCMoHJyBUb9tyLwp2qm25g/iOQ/jyfw
uXWo69S98UPLHWG6XWIHNlZFn0P1izClhCoPbDFeWynjzdycu7eQuRrAXRDspIcH
WIrfBp4Cl5W6O9mH+b6qa753Lwmi3mUuUKt60oDkryWPFn0ZWt4zBC3Ua4/0cq86
vt5oX2Ld4/7gnOhNf39pLxhjp5AYmg0b/fpQ5dlIiGdWFZpagaQpwyXuXAJYNqJP
qXyPFxD/f/ZVh86CzhulrwIRgdy1w2PTvqWaUSup/ir2H7VQHqk5jFlfjAm88FEJ
/7hj1njGjIugx2F5eVpqNr2m79+ywDjqDSgiENJXw/vkBkncH0mx/a/rkzYsEU+G
skTSBLo04jEn1T9hp61slpoxzWwo1Qwma12FUEpeIXyDU5qfVgFUb1hA7TAi5LY3
LEUE83Q/VQ5VTkq/Aea9oSHx3+XuyqqLJk1wG3xDjHVLeaEUbXbGURjQZC/OEQGO
b+wI2/O/DDv3gpz5mD4UKe3chtLsljjNuIK+10lwXW0Fnwe/4usg5uxUzDU0fXZr
I+4QJDpwZh7gYifRCICMdXYZ0ZktK0NbNiFQFAfhglPhTpKdT4JFSRx1mnuzV1Pf
g8x9YF5/zw6Nto4MpdceU1q7uu2UqrFTDXokINX6NlYD5/j5MTZ7vNFQH7ILKfUt
PRYSar11XKwhYoX7HDpA6GBdvCWkijt78UEy8IsvcLBTFtE2NbTcjI+HC2sjwEw2
1ZkQGONnw+IlLsqOS5yQpjyznQBRurRQ7cNS4N8PqfQrSe7TXO6NET7jv7FRrj6O
N39mXDi/w4AOB8WM9vVOaJx4roJq0PP06QmamQ2BxuhSzJ+AJd78avurB/RLZQDC
ohfvyVV5zxBNAglKibmE8o9TwL4aOsrRqiZdMtdXiuC+pg2BhfX2pRm4qaeI3d0/
NtvMl6h3JNxsv2c68kxjJQvW1rd6+e7fI0osIHpSmDGUr+5uMI/sFShTGihhmkL0
Pq9whG3yKTrtMoxY/xTKa6se7uKrTBDPqk361kBOZCYGFlrIfcjVrsekXeaIZafJ
bwtuuzGQrHM5Q4sRaooU1mbdAzYpS44roI4+I6Y0D0AUegeXu8+bO9yII0+Jk0RA
znB09nibX9T3h83KvnHGWf/zGbcmQntGXxNbKDIVzL67I/bg8nI5vQ/ddt5Jreyk
GGKTzw+cQooOTZxc4yoghAdrkcOa+9qv2T3MLiE0TYEKopoFmI9UQZ1tZGWITleR
LB3A+11PZnrpM6oor/wbJGCSIZuRtjADorhDDpppN9ghFcmOPe4ZSSuQie6HhGQs
GsSyMKCk5mBhVwEkpMCOrTgDbSUx1NxkRx1HAAq+PCapvMvUQOPVPZGTPlBDhtH5
tn4VS96euzXC0sucHoSdcVsE7RVXsr/1fsuJWlnPcTdSrHE/iNmiAw1LUwkrtnEU
U+tEeCrFFA1kAGR4al9yP3Pxrpl/FwfeUSLpauUqEFw4x1zblsjIvTc3RM6hYlQM
wjADrj4bnHEXTkyGqJtKB27MnrEoVH3UEivP4D+3xBgOSUzcpx6YnYe1DvIbO49q
QNqYWuzxFLAeK3eFsDwHzuACEwM0Kn4MN1v46YxqLoxGR70NhYqDCBDyny+IhUde
axtzOrElFzH0Vi9PgH+Lg17V2KtjGuxm0OSbVuWNUkDXY6+rTgaQz+zEb+J71Pvu
wmAWtc1nzo357dOrOvck5n5KipzFEaGKOsyt6Jjjvq4OIouR1BNxFcUyet247lXK
OaWOxbXU2/uSFNepfl3adWrTnMq44HbIBFDSXJsbqUpIY7V7PXniM3xKNP3PIIvf
GvO+U96O77shaOsHb4bPK5FPBZUR3wABXeVjYBWYN0ugzPj/2/HOdm6zAbJ9+g7o
UI1lSjF+r77wtrBHDnzz0ub2m7Tgao9Ck0n4lSlYA+uRlS+DqhKtNGtmVgEPcrzt
kHKLtfI86lPDJjDoZlazAjkqziKvSnAIF7JcW/JWQHT9PMpZQBMOSHttfWZGbnqQ
fq35M+vssjhG26Ui8uYNQ+KwjTKqhyjFz54mDXgH9KOda/XPhz7l1I6geHEL0qsG
Wjk9Q/SKthi8/467J9DS4TeIkAPsn39Hxhqx5idQH9jYqX3SbDWme0r3SYwi37yk
R+UGcmdqcYUv3zE8PbKq+xBqyDDjYO5f/wrRmvY4JmzE97HK/btTiqi4ndp5Tdfu
a/UW1UJNvU/C4XyPyEtNfsXPqN+A/uOAxDeRqNZKJ4KyQKB/7bBej/dOS+j3KALI
qRhJdfi+coJSulIyyfalUyjELJaXFq3usiJAd46nijrwPj0ArV16O+neHA4cnhQr
4fGzJg3ttjgVP+KWk78UM4dmBMysYJVR6zQh3TW7kHWwHc5cR6LiL4VaRit1in+9
HK3n2UJcE5MgIhACFzDHSBLrRLfMNbWn2RLlXSp7apzBNpbXp2IgK9mIjzIVCanw
z/M2ADqWN8Tz6rWcyVOW3hMwuBTW0WaAb/VFCXWpGkUfTzIrHJ4YXBG5weCNLf78
C3fUr5pYsk5q592vY7DcHN+zFDVFx3Vt3tEf734JI0vcVjOTYAPbBjlZ8HHfSylx
5eIOX6kOKJIOMIcrz8NKN4JDXtIkdMkBAZVyDyYXFUU+QN9MPkF2PfhowRjyEdG4
qY4foTQVt0h72foSCCFp9kDlGGyU6iz4kV+4dwiTxEOzYSspyZgRH3U6QbolDmq5
wipJCNew2LNjcQ1963Q2OmI+MNgOAm2vW4DZPPVpAyudZQFuE2PQf89bh9dqAOkh
rEXPx/4QbQ72spj+qQhoueKI3hdaNMUK7oKsk4xkJUyeTmnWeoO7IkxikftYfue3
JhKJfdd/vCb8j216O/LxmSm2qSLiBCsGEcRfoducN+SKUjhDmhKj4nRnsyIiRWxZ
WkOChrgqC0LReQUk2mTjvQVvy7m+pcFz0BC4+mWkGoQIrwuk4xLfvT8RLzU5nefn
IUodf0Zr7OeOlG1Kf7i1cX/m1CunKe+qrWjNYcLEg/CpElZnzbPmXq7/Yi3bX/3F
gDWrz0a8ebHZDO0Wl2MBgrXXMDgboezU7WeBGDIrEqCTqlL2hq3W3kFLs3VjWFrF
4qsEByeS9Ivjlsq+h39JAmHhVq2i8oO12UDV73GppCuYgOktad5H+Zu+8JjSTKO1
gAs+r2qkeeDgqjM8Aoh/fXoDfHtWe8m5gWmkYt5YubHI67BK/Cfpw24rq9cdoLWc
Gdjzv46zic0ohMeDeJxDHgEA3qP+/gWVxvBjlk5nCNAQHx2thEF/zIc8SQshJDW5
rnY6GQYnd+3xiMCmpY6NPLoSczqO4EaKhNOGzvU0c+MP/5wfT32gb+ZO0kUx13FJ
Yf7lV2IaeMElYUOORNYQBeVq4+0g7EvYMZAGc9UysvlD6PxL+TBpBfQy8I8CO35R
1BJnknGkOmgknDNWVs8A/PKT9E4KUOWmBelaOcckZOUHiU4a/xXuqnoxmzCHfggI
an7/Q54lHRWmSpI2rNk6734Tfr5I+s9ab3mjZPGckbkgeHiJNW6+vteOYmxHeA0D
m5ZKEvoOqUuFspDowAI34UMaN/DkT8TsdoWD3m+5MvSXEDvY2YccXV/XLMm8B5Iw
VyXuK126iSeP9SwAi2iiQF8Vdm2GweBIb/tm4c+rQZeGk6mUoHTk+fPBv+8Dir+X
t6hVDKfqrr64LP+dO0YwRa+qsIn4/6taflt2cNZRfPGxu1vP+GurXEhJrx4F38ey
QHzUNwC5pnc3XfNG3R0SkALw6MY3XefytCuEnOT96nbWYRDKcgX1+4gNwX9fdKKe
xSPYvkxvW+L5IoaC60meZ51Y+6Fzlu7J93zyeRKap0ddPX6KMx5OVAK4ee8slkPE
dFpuqFQAGAKCbbeNwaf2taPd/yNagdu3dH28SMBrmob/MalT3uZK6Dz3IHSKisOK
ueNmrDwwbby78OEhVothKsI8v48g16xP5JiunJq/b/RxoZQ9YWYqenRpglUbRiBU
LfGketODzxPTEqtZ0HP0W5RIM5v/tsBM4bjQP/WsboBiBEh6GetSxp8M6QnybCcQ
zIkoAwAODb9kLrI494QeMFl46PJl7W5DEHc/440bfW3o+BTCQbarcG/1pXFatXIV
T2UmtHlFJWySH2Lbl/ELha9tLIFc22bro7aUpC13xRnmtP3maMTsq+WqVRKZGxh7
M/5p4isgOTvYDsrwMMc3yWatucRGvI0WJ1jAnQ2UWQr12ojnfHz0sYUkfRjaEbku
tSMIEXKY3gDuleuFR2CaILYGDv2XPM5m1m/C0vBPJrqkVNWUaCM+8Qq6BTmFzqtH
NWHrqnOyOSuflRrlr5ubZqOLX6NCw47QQqgfHPNUSEBTlLahXJcBTlGc3DxYhvGe
Spd6R6smHE8VTxfbgLrntiUYzpMv9zaUsy6v82yPA5yyc9dsHZbQ0VMeegFykV1Y
ur/HuvglwBuuXh+UHVu4ttT2WMdCp1odUUrR1U3HnG+bUFEEokPJ+VnZR5G/eQoW
qvzlsPPT/sn6jOdk3mtbZnsKIueYbo7p+4dSZU5DTAWK8TyzrKHwIcr3ctUGe+i2
+wbCF0BIl4RaKCyxr6rQYFikQ23RIuIa8+1b9PfZ9pHDBaOjepMLdNuxy1DtTBMf
bvOXYzKuqpFaTakeJ2P55uJJIv0zCqj5El+U9fiFBhqaflNQX+vwCvzeaL0qEK48
7/7JzJgcJgLnrq7fyhhxGImy9uNgphp7U2kvCr9cB/zJgsBj8HhOJXdZ+Bah1Dw3
Z6WjvdIu9c8PGTFxUMOER/KGOot+EFk3wZY10BTuGf3eHZ4neTR2j02iO5dsNjxe
r264bBl+pXWSoyTuOk3k0wa6b6mifGW3QEAcm27W2LSzKcwE5VhNGzSuFg3OYIm/
GB2D1/U9w1N/ZPUP60Bk5y36AqM+yxJ3pDM4B9ZSn08L+XHimEFb0NipZWp7T6AC
z9HePIV2GQOgnn0RzVOYVkt+oWgUmhBXLQtz6V4TQ6RTeSC9FSNa/sCouIl5ZnA1
yAQJXc9Y25BfJG6k6lVmA0TS1HY1RulnFUjVj8qo+Kb3cWl5xaSt04DgwH8cEHtC
4E3KMP8Uu1INGWe8RFczmwtUskMwRdmboKdc3xmYnNaw2QEksAFpv0nNTT4nBmBE
AEhqPpnPjBhB8++Ti1SeRQuCDRZ0Lc3s0sWnJQfPm4ptlrGH4LQTRUW8U8zvEaVq
7DrVv3KaReMy/2A4K+LmvQ7hOwvjKFOnbATvJqHxZLnd6P/Vt2Jgqh4Q6t31MRJ0
TTyQXjgCpjK4ZngwKe0yN6d/xBnTjmtdLYmck9ncMDTRBF/FUlNkTuC0xXO+w0Jz
pLibY+4SMbBuWZeCpumdRYNX6TYvc58wikBSgrNq3Xo=
`protect END_PROTECTED

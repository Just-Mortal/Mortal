`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNYljRUsyKd5Vc4+zmt40PybG6ZUOgObnVjCOKs7OUMp/bLELA28Kdb5HUcb5eJl
+GElpCyZDbcDrg8RjT/RIMeNX8uA6gcCLeVpnuN2mJ5LQZZVLXX+Zh6YuYdesyJ8
azFkCyYuaJtx5UvTrweCRYPBEs2SN0372HEWNsCablV+toSxQzGDfcuNkZ35yokD
0KamShi+RGrjLe4JFtXHfBLsVXUHb7KnlgDuryKP0Iq+HCnpiS2gZWsxmxRPT5Cd
XPUfMXQMBezSHXnOBpriFGbUpY5PZCllDetvTxagjsuEVq7wCk9FQWMf0aFGMIyh
oWGUKAnH8o8RDTVmy52ZvQ+bUdHu3vZlySK2n3CIUnbn2ZWFTaQE7hpXkDS1Fu6r
9SH3HbqRGgFwaZ2tKLpCQY0ZXwMZalKyeXgBEayjP6W35y1HoknfFhqe1P639wIS
S+rVyBKqh+BgHayjBfJIXB6VUrRSD3RhNXzIUmul+aUhfbFNScHJ3LVdjCSIBwId
BhUi9hVNtD6ASApO/H5EbaVdc3vxb9/jV5uK1xOdrlLV8+l4ng77TnyLp6UAnkqB
kVshRxFe/UrkGGHmGBXhK/KV6M1h3y1yaocCXJWkZ45WDVw8HhFoavh66dJLAwVf
FeS/oxP+nObKFk5tvv+ZPagkm7KexE1tlJ/GBrzL+Egns8HSFrqn4xMLOuYDNvgk
SvAk+fjHdeopd6nsbW49qgxZxemSurx6D3/efqN+GTasZPZPZ2A6/XENAC7JAnCW
2acRgl9A2w6agOvCtAAIBQ0Wp3eA8jZ/sWpCzymGpSim1sFfWkOFzCZ6MN8BtjrG
GLaPQzU36mA0M0mOlt74Hga9uIbGZPMZAQABBb2WegQ9TA+HYjtbrrOt0YwhWFRC
YuXJO0o0T1WdHNCEtODcz+9dqDsJHWr8GG0rYA3aMmag+YOgUNB5b/cCB95thM7t
LY8p+08lGgp+GVuKpztr/qj+Gift+EGxWKNDfIq9oBygZvrwQehl7QMu1YFmf6Or
aBst4Y2oQc33FMLx8OHTFRP/yKC74Kzt/oZxI24DGn3/L/9pwsNHsX4ilTp9XkEX
tkJtubWChtbKnD3Y7yvEGJU8SOTPjqcZ90hEg1fJHDePLM23s7IHZ4rNLNWdzDA4
0QUxBHWgT1fngKCxAEEJVwzUFxG3N2EU58aDy6g3eWvp8oR4+fUMccx0AcfN7L0x
fUi64Lp3bUi0VC8Jr7ulIju/HkE1NCmHXFE/T3rGKb4sDEyZeEJXnU/LKYW6jnc7
U2bcOBZrt8hT5Og2dno3JTwmW11Pt8FEHnhgukuqhodgCinbLW56ZqIeVOoQNeJF
oJicwwmE0RicW2oTFygVHzkSejPX6LZPyWQXhIPlPNlpsxpoedJA9o3iAnn1OLkg
DbvLNItQg8fpFVaPgYiqzYT4la5BLPD1RSrtISVuy1vho3HiB0A7W7Tl93JHpGMi
QG6VsZeykInxoQxJ/kIyhRGbQrYGNTR4/NXrrccg5x1oNhEGaOk/Fql6HRWXt5CU
QUZnZMV8bYkUXgE2zx5teLlYJbfTLasQPmY27XDDvTNplfOWIf0thrmw4s6Beh0E
JLZqmR3JwTTdpIS66qV5SXXAuwrmaHk9Pjk8y9aHZIMjSR/2bYSNsuXAF+Zqzrd0
f6RTD44ckxvB8Jc6JU/orrEhjVbKM8mrTscff0oL3gFSs6HJQ9nROqyiwcmTip7f
lqLF9fb2iTth7M+aP1gTGcSVA35Nvr07VQpRDetAmct5vgY/l8GJxeA0x0to0nrd
0WGFMnYMRZOO8AeiF3dbsrhhLxDnmjzGn+xQyLJHZjm4MFPpHDdF9GP9tI4CTg9W
B7Ty7F9ar3St+EoIV4mJ2NYMNKHmKh4nUp1tfIpWCpEzN/h6rGJFKN+FQBcbe5j1
zP/Zm960Rtm4Hn9kiaoWaQ8P62z9mmuQOc06KWJ1indK5DMYl0E7c4lhNonjAz4P
CrMcjMIFhP7bLVWd9cTrX8LUk+biDvwZRBWUB8d2uSdCmTHAC0yqjZoyVzatrPwk
nl+PjcHz/uErf/yn4yLpVmksQrY9VymEmX9j1YsiWUFE7yJoyz78dvou6RrmmuMZ
4G9scn5rPgm+mym+n2px7hw7nyGHixgRxy+WjbnG4hDIfIfr6MkMfGAWjw61a8FE
aZJpLIHujB04cxun+fC/0LIV9AMf5DWQn0x2SkevapEGS0v8oEMN2idkNJQfVz/C
5frry3GmZaU09muB7g9MBvZF6b84gEFO+CT/+4CSVAhn9bzwYtv6aBNg2/HGYcWD
p1Dh2EPU8NC+szXB36JgFK79evtcLEjxVhFouU1fHfdAp9MEr55q+UDA4kgqyw5T
DHxIPr4vzzNUc7C/hMFbtQaUIX0ETGj6mftoMP+nDh9Ljw92XOWLFahMfQ+R15Zk
N+QGeeGRvgP3g8ITASlhxuBOFQJxsyGxbjXWG+rVzymTokwq/Jlgsbff8rTkLscW
8CI5QPBQ/FMQBvE0gmPEmb0tsLGOauL3tloZood27BPNxaHAKnZAco1SE1W7xyya
IWwwBLebI1wSDh5Jck/f5HkHMk2Dbxq1kkDJzKwl+WXzIFSJXfZv4dKkpE1JtlTH
v8N2tKqC2joiMvwuu0X7CYxmxe3XxoB5Imso3zk53xdIbCSq2DgEi6FxMEu3hzsY
RYPvh4xyQqGmzukfEMzAxNFU9y1Kjv1o2Kg1Wud+2cLHoeG6Gf9Wua4R94vUYRNp
wuaFj+3NAdNRFFiA9YE+CkOEu1m8djXWWP4j7+Hdm5g9dgO4ATdKZGxnIiO2t6Tf
rQY7TJS2gjRkttqBNbeC/YlM7Mp36uVKqnuBaE+SxO+vl9hPZyHqMEPaK3R9fPMi
l0YLygDkaZ4rywMBoClNvtGchyE/EaTKxxVt4SvyVygGADo1E0xb6GL/5nuuRMXG
YVQ/+Zyht4yOa5m+oU+R/pOVFaE/tphTtle18Cv+vWG86flOKyM77RqwD2kmfQ1q
P4u/TBJwY9j1Vp+tuq3bjxiJOfoJPk9B42u0sEBeGia0sy1xgsAr7ft05+ZYA96p
SBbr2I8ImD/GEkTFKpHz/e48xpfDG7gCTbLIrB8Dkt0JLquhreXP5bLyIR2edfnr
duR4qwzLQbRkhQIZ8U+OolfYlJ6LncKvZb6xqoxhhBGOVxi4t/0YDOXLeY4O76Mm
/KNhS6OqqkC0pKzAFZDJtqCe+YtYRXsHRomSNvaMXAL45Owval1eBRP5kttxgxs9
zpH3CZi0xdtwP1i7wuGRiRI2J4gqcdM5PtTvShMt1P07BObk8RparIKl7saoEgS1
Bs84485F2ltXWqmKAqFdUidGOV+fzCb+rT6BzwEfCBDdrejd/5Sv3q9wYQwK56zH
A/DO8bv1QVqEJay+glz9XSYsFiBZkS9/PRsu7CnD0AhiCn03/PV/ujwT2yrAIszS
lSqe/73QdN+lbIQYBoa45GeTK+Rky0kX3lIIfXS3t63s5/Vh+iL8PIhjtbhWME52
6VkVholRYRbmLzH1XAB+Jr8XQ3FiiprAACd5v+OCn5C86cMK2WF1JZKkLonEnjnm
Q4EkhxItfa2fy+7y/B6syDvW+0Sv0K9zjsSmHOc4KCUnTsoAtSjezhhrwuiuxqQA
wTyi4AHeM9IXyXJdT5cfSrQqjdV55jHJMAgj2+bqSxE3E8IchcwVYEFdUU4cJz3E
d8xqa5ks9OajWy59eZumrBpkyhkpXPrAW7e0yDm7OuUwD+syAtB/MH+5DEEkIbfa
GdKiC8+500gaThlxnHZDq4tLbeSrivBX9RB0HqesCpb6ac9Y/9L4TMvUqZRmB0H5
gE6mkGL86bfb7fl4bTivzKdQD6RTrWa6JY12zImr9BY9kk6A8sh7GEEsQI3JoB3a
3b+XUSlLTJAOEhdFtxfur3pWdyUpCHPH1XR5M4sbHRLmkA1EOUusinIFonH3SiAx
l9OzeDc0fwN70Q4vbsMRRvPwNNi1LL7ZPMKDMo6B2XZOdydr2+Uw1cgRY06+XNu/
o4N8XAazCkjp6NStE7GsGOaRmjVRXDrHEbsp35s89EsgFqqbbLEyam7b/T2+0fdc
Fr5W3YMgKq/sru/DrwwYMfvpz0Grc/QtlGAn7e0kmG2x4alefy+Afdj3I3C18FN4
8mAupTWR4phIheIL5CeP2DLxeF+NujMveeCHKbcIRrqj9lMzcqEq40Z0H0Mv0xMy
5Xyb9HcAoMqnHzJyni2dFy2vZQ9GxhCMymbAcGHIQvxOSTaACZJKacRJXZeq2E/n
Mf/0jrN3pT4bLGznKxfYAjBhuL+TFe9KnxBuzbeyqmc30V3ATQsMHJrfwXLcMMv1
oYifWw4CxRCBrp2g1QlNTYgwmzTtsuMQCaL//Y6GaV8U05dWG0z7UHJUqCKsOrVL
Ts+cjXDs1PircU42nzF58zjfCLaKCt/jdtYROW1SBE8WlmfRNbPSnBTnaEz/ObDl
9jCI16nZNhqEcgRP3r33vIoqpFLI1Kz9IJNOWycZa0apwLpvpcwj6rjn/im2SqOq
3qRqcnygiUIM/7qLbpJ6r3Tp3XkK3DoEzUoG2x+QniYIom1Lkv/9OLjLqo2iHsXW
dIJr32TlF66m256etld3l2wsdotArVSQbQqeO3oOrFrYf0ig9yuZ3ZMSsgf1lWdy
lNSWEKwWSlkYyg/Sfo14xTlyYHHUlqvIFz0IDyYHptksFBKBWHU7ORYKW8/J3qTs
vI1VVituBrd2leHvr39NXZpcfjypXCCrtrqMEfRWDD77Ar+omPzhEfUa70Sk69Yp
zryBTehwzCistY7EKqmPhRHm7J9Z7ytMVEwuxt/RuDP9fKR4zpeMddRko4up1FoK
EahqULdRoypNbSj6M3oUetieOW0KecMTPal173iwa6x08jeJVLYs9Imc/3sfjlSi
KBLN8txxg8KMESqZ5hMVDQ+YftHvruicEKSJ3r3wlCg2j8iUC02HXD+l8x9R3DYr
rhG/cx96dA9MIJ3wCE2oZkShXA5IZ6Jvr8X7n9pk3KoUmoCmpDvjGNU58k/jYFnR
33tjGh/HnZTrES6Mk+8imd0MGN/KCgkyDiasQAQwJbSBTkjMQr+ytt7/6UWYe6Dw
EGyW15ysWhsKHtmBmr0Q85uTjqx1J+TkcspUCmFtbBNHbh/pbatRY23bm7h/lHbl
GRJR/k1yEggjqXSLrDtNmWTuCLUVTw13bQyKuxEK3OpxUKBTHsJoce1UoKcYUYc0
ix86gDKCKbUh8sufKhnj9lU7QH5BX9KpFxa/YC8Ucj9AzB1H5IPD2qBliWd/r9xv
QoecOgxsqCkmiCgeUy+kRnKgJalsjlDVfgFZ0Odj8+GJQbZQ3XnMlNWyoXWjBAGa
J6v7Rwm4cOf0ZgfdJg32djolQPk8ioM6G1a5agp61dOLjAuex7Q/L9Rw5j/zu/e3
UV+gvemxsKu/+7L1JyG0KGqe6+17J8xeSr5rWMFPxRietPThr58uhJM9s9DTRhpi
FwBZ9+zaImaCYUVYS9Y8Lyg785zRXkgE3FfKo5lTKpSFj0DRtgDHpyd/n2TiHLsw
kuD/O/pOJFvKFVAIBiLYSbW+CF2DA/wjJWVyuAawj89onUDe8mIiIkEfsrP8veUk
jU50gFOw45QpL+EJLqCIw0whHr7NXi1yJzmacb7v8ZXD5xZKqRaeXpGa2InYFxMf
Wx0CIcX3ePKVV7tJf3CVTnNWIknnsBJLR939m6EHS6c9LG6KG7EK+6jZFSXu64KQ
D7CKNqgDchaOiw1+kMdVKn273LWD5D2Cc3fedmP1T4fE6PO3gq02+bACcFSK+kRz
Yk0OZfRnVKwgX9qgA6DBlDBkkyLDhxcsgUtOAfxP5++U8I2TmBAQlnAl/62/4Ejy
+cAK6KCEire1j3Q0J8IbmTFC7D6LslKxB9gQ2s4q9qj9OYtTsEE3cUKLL323T4Dt
X09sdqIw86sWo9kZKrHfj1YjTVn4dsox0BBtKEXdRTvimi2Yi8aVu5lJg/7AL+dU
`protect END_PROTECTED

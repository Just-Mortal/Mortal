`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hlqRGAaJgzlBoOj25hquwZswyBs2mRwo+sE5GkdaVx0N3PE3SIXy+B91/5y8cEPg
MQTwKJFHUeGkN8O99T09L7BmTH8DTCybLsX+m3PYY9Te74Q9R3e1TkvEwR0E825C
nspO3kllOmSts7X6rDd93Ls7HuCCSKjbXDlrkY1AzNx6vG+RQ9kB6WkSNvUtx29f
5fqyeYDp0nI2y8BL2lS/MhnGWtywMsOKC9bUEUzNvFZxci+oWzsKy0xfw/eV2FhD
XJ3r6e82AgxgRmOe/ZmnjVe0r2drkpsG8j3RzK72GFj1U3I9GucoJX6OHFbD51L2
45B1sBfijyVv5KIJSquf84nfNMk0+ss/KrZMQv4Y/esSxxtgCrPFCCiNstiZux9/
R4fLdcW+Pyrx2c49ZNjo6wQDODzgNp4OL8hBTmmXt14kcuqvySB0UPZRiqSohwk3
eI9cFHiA7E1/AaS7V6a43aFxZ3aqn1m8bmYAvIsE05r0k0BwQdAeADeaH1QRgHep
lNnhm2VrBYgiQ8dv4+CNL5QRuW8kFwdB/PWP+7Sucw3ZCIU4eN/3xuH4tuN3RDZn
6QIkCjBGz+wjPV27kf+MwadvCmB4zIcMAt74fsnI7lsVk9ZMxHqjNVbbD+oUwhvn
J+ucxK6J0ZTSIERtV0fEwBGtBPdLmtVEqT+nEcTP44i1rW5wRr7hVbwgsWaiLKIp
3TgwXf4VqCl93pfnsYoZ5mztme9Hp/XrQG9TA4ZcvNDkUZwmeXqs0aGjEaaYULiW
L37vB9uBetdIbiiXlTp1I/bTZj58cA8JbdAAFvqU03RtU2f1f5qwsMRW3kF9+FpO
aqA9GCvkIvVCJzJ7nun89mcqXdZ5MTQJ0rU2s8k5YLUtlvkkrh8w4WNUmdy12imq
5zsFL5lhzte5vOTnfDYbxAnj9v/NkzumRZsrZIKJPcz0vSKE9VOb4hIQywWS5Wcm
o5XuIKOKm4BwlRqdtLnvlyuZFFXR8yQDzpavKNhSHavS3DA+b9NSwdV2nDIpswUm
11fcEKR6FSTl7OFPjvw77HTDhy7uffVsIuFsuO4jMs3pfxgwmYXb0g488D0mtKig
qxusinDQ7Edw+OTlYLvCHe+ub9GreAyf0lbG8pfQ/j8YsdPMJj0iv9Zp1NQTtdmg
8uguJsr200f2A4tmE1BI1AUHL7Ylku48gtK0c5vW4F+RCFnq49j+PZv9fXeuoXbm
S6G6qr/H7kzk5zJtFhVUwKth9rlwFqQCPOn/7e64InIkGGx594MjvVKBQpYlZQIN
yBcc0IGlyo3xNgi0R5RgR4rSshB7bRfUU7hinGKQ6n6/2cZXV6yihmznM8Lx93aR
kug1nfnl9E3EBp2hZc0ytaT7bbZKat4R//au0QXBg+HBsBaPSeHReP+P46DGH17j
JJUGlZMit6eQOqdh5Mvl+KEiQDuL/XnZCbY2WwseHSHmKFONX+85yPUDX/U0Sd77
9RpQaELn77WIv8DkXdpntVVN8GKK61jrQBYSwcu7L4YTVGBkdjSjzlwda19V5qsG
tBdcb1YkvOXOl7+1C3HxGCIwtv0Q5x0O8qBeT37w6MR8DEi80+mhRV0fw2Zx5NPf
IBkqRIpDGYdhVSigRYzMdcGlR4r6P6oR9iy90ueYYQqnwHTCnDTVl/aeDOjbzkH1
uHgewMMKXJRkQtOFn9sBWkzRfwGfTGnxswzKfkO9TztfQqDNbLWT8cRisRhgirIr
zQU/pdqRlECnQ1F8+fetav65h+q7WryFgMwV+ZbEG0xUdP/Cp+ehsx76p5WBteQz
F6MIbwe3tfTP0clEP2uLgjkz76kXnqdlwUs2n0UZTdfwIy6kROhUKqa0KMnNsGJP
mfDrVDiTG6HV7VF+kMCoYiahtkKBtx0vLYKN6ki5M5oc5kUqMuKD5unlqcJabWzn
G4CfnirQRp60c9h5+B1JaXvmgwbTiQmi1mLf5MTrKcTSVOqvAGUqybH1oBlbaTwe
OOTd+R8Z1MQbgRd4IAWXP2oN46pZKByQDdlYZmTDOzfJggepX/T/jElZ8nChEK5e
hSY6aP6jGbrZh9d5wSP2cnG8cwbriQwrJlR2z5HURrWPFe/86rXaR+lLkeEl2HyD
cizdZ3CXjrSWhn5kd4PRpb4IMmU8c15lizG0XEjb5YcFQAfDJeDigXNlFyo5s6Pl
tKwaeNicPpRCM0xJiNzOHEHz4FlLb7sF2fBsRhalM72ebxlN00UtBtNtzJYfBLTa
RDrvk59Rsu6lI8X+vKSZMMNnWBXJMzDuSoCb7F3wNC2vBBIbSayrAXGgvWBW1dE2
0asAjMVf4lYAAypUf0nYiR/MZedsc43MH6lsoLLvwm5P2GK4Q5FpJMH+ntrzqnH3
hP2Pa5rakqiXdVkjjoGe4NXwzBDQ7JdFNzduk8yPbghG0PG3wJ+07158juD6bfkK
h0FOH/tzylYAsr6zQNay6oM82Qs+P0ohcOdg/7gZCqc6luCzYaNNY8me5M3cXlA3
djRYlG+Q6vq0Ti3RV+69e6bXKiC+8qPQd2np2QxGzE22AjwgKTb4RfLT+vZZ93XP
8mMe3MjvCrzZ5l3jG03c1l/l7ZiLYEk9482lOSu4jXWHSWomnIihXcv9gB94Dogt
gZdBMQeJ7RBdfSQZlO6tgL5TPf8Wvh2nKPXtyheCUUZhldL1pQhZDsReNrXDnYCC
38wCz86/Xfop5/zT28CVNZE8yoT4mQhXg1P2v1sJ80PLw4SGpcKcw4ulP7Vu06A1
AuW7ClbQg+2Davg64D5IEi3vADYB7Akg8HdtZqbPNoyJuPFhbbTRjiD4cxrzftja
wxBjIMbmdjV2tPD9N1bc6Da9k6ThmUmg/dzf3+L/dyIPbAvWJUpmYTRp6MHfUHcX
qTWcCvt1bRr16+hAplAUW01Vi1STDkJ4wTGoN01PjrCNvkllc+yIokAngYXRIEUz
DTpSY5MGoSqlPCoOjvnJVVxku5yEP3rd2376ZifjTETiB+pmT3dmQPw9jNu6HQqJ
XE7Enizv4eMwUmg3u0GR0xBf9g3mFE1tRI+kLWhw3eEdXO5vQgAfxDHKfWWBJPd7
0V60GAoQJsyFuMUQVnSKF+X1NpKpCUVZqE8ZLSptlVaV+SbWYOcaMK7+8ARfePLR
w7jzvr9eVrY82v07tBXJt2u0n4mH+I0d5FCO9dAuD2tIcCPhj3YsXDutmjAtjGZz
8VBJOyV0YmgFDqxPv9gsDjcq3y/nTkfPUbIS/XQhiyv86NxCB8arPHz6GuhZaC20
Qm/ZHJPZeTy3F+VcGqPSAdjHnDa9SYZa7MsC+mcV4nlNrAIqRYDdjK/+IkreiLAE
7Wt0M6tmAC4buI0Tm8oWGVVhKe4yKlNaCBBVXLS8UhQxhUa2czMCfJjUFxBBNplK
J2IqFFQZH/OOZ5zoS5LLqdRDZBUxfLSJUN4JdHpHARScWKG8ybz6mnqh1GItk4aO
eAMwYFd9kvuqhFXTGsk6aP0KiqWq61GEEYTIdClpJmCxKoodE1/6ppzamKPSGx1Z
gggqv3JXwSmjvOpKS61D4JDRcu1Q+WMyBC6ATjS/5vD+mmAoaS1shooWMysY49tO
1gEdsIlHBn4yXxqvHPCGpul8kmN5/s1K5ZY4rqv8v+UwPEkAnx16YKZPgkfelvEA
BoU4qGy7K33kJbwzZexEc7H8V26oyKuKLfrpQ3LVamdTCXHEyxIaeSjIXVHuq8uR
f4Wpq0dBuYwKE2pDTUkDl8TPjOSen3rHw55ppPpROGURzL4g9C4sHiFH3t2TP2oS
z7Tt1QU1A3CgpLwjo6sXKNw0DOXPTBSU8SOd6EZIcXDzHJuED0b16z5uY2JxbIZ6
qS4vnG9M4sdBJBPESEm0P5TVK3miq2KDT29siAp6lEt3jqx8qlN9yG/T80IvLCSy
Ky+o19n6k1biM5zF0VT1xznUO45+c0QqymAnJqgd8/9zo+CthiAINfjaJY2MC4Pu
Ze/g7pCV180IME8zk9kYQZz/45XkUHGM705bre6nEt1lViNhmThUh3ISv9uNRDhQ
rSTIU8gZGc6s6hWOZ0IBsU39LzyYW/qe1onxBz4q+oRfzvsljwK6leB+1rqQJ/P3
TH45R50OJFP6PMr0Mh8GAq54OvMgqOKoC7o+2SzxuJPEzwOULdLfq1jKXWwWBzvg
qhN4ZYhmJ7vQOtPB+C+aISxdZYPWe4k/E8h/FhphaP0Fiv/kbhCNP8XsNmvpSaUq
rFAq/9mn7tcKaOtRFUeUOG6WrSQoC8upDyG2h91mAgopST247BJNBYfyz83v5tHX
aL06IzzOKi5leFR8f1TqQlT9WGrXpPjfwkXHKlmE/d6JYTaRCkn2n6rav6T5PqPl
Yrh1e7yZe4cSQOiCVDp1txVgFrcAWWoyy1sfMvEYVowJ+xlfJBByeJGJegb7w+TT
08rs3x/YflZWZnqYZP5BomgvuZ4NlFHVNW6y27DrB+Jwy2HmNACzKJQHyACuwhSl
qxPdNQQsJE9RKAiaqnzN0XCPgUP+JOVT+iWBPl8x5LrXkpIT3JcxlJq7Z4XKSSdm
PI8k9bGrYvZssh5H8ohpO2maDY1OIWg6pI4pak40Na4kKi7xARv5DhkIRDL8iYCN
arJZXlzf3wT8qHBZhPBlCck7gMq4AOrI4WdgNhDDEEUzqLOUvGlKxwOixXO0SS1q
oxvDe+KV7DEXzdie1oq47I9MVt6yIGjI3rRluVFIm3/F8N3FWz4PlQJw+64gpkEv
ZXsHaySc7Gqjr1CVdK9qbgTvT2PiyWSzoTN/Prog2ueE2aEhSO0iGO49IW958LOt
UXCdhJcNBCNGNQSlWxJN4lE+1CYSxj6QnsuzOKM0uwNwPqy7qK+TjXzu0ediEWuU
uoudNYoixTvH6gUZSnWcmJpueVu4GMnzFkAmwzEmHxp4E6LeW9xqwY2HLXxAMCkK
W+olUqWkZSwClEav4+oJKScdOUhXt74ki8FlPOCUUmQaLhwQQ9wiqCGa8kYlM2t2
rNMFV2p/nwp5A699m/l6Dxy3NzSp19J3t+8aZkhaOldTqJZxvA7Rm7DuBZ/p4Zkx
qcDhPEbv3KPE09Tlw5FtBFDRHMASqv6MurmwXp6rqntA6xCGuNvft9PPaIt81Erj
5IgzCtjQoHfiQkjVgMlSk70O3KAv2HVMxsEgzBVhR1I97VIByX7SwPgF1aBlfMx2
LPxyZABEqZknuPMd0Hdxz89Awm61bzqwxC2UfUaMLGa+FcUeABY44KrWhpvBC+L1
YmXN09RwtVmH6NQcKLmnNH/FM/7Uii2asZ5fd8Y+L9vYTYhAyo9uxsLFehuF6DLP
PXa/a40U40nkMpCTCTgQAeRYJh5lleesT/0wS3X3qYvgje/xPNEQ6TLDeFxmg4IC
CiCdzQwTX2SOgZmMYlqjr0GXxHZvsc+fiMvSUOLQvB0jZC6+19NJtE9IsHCmZHgS
1bgpK8fSzE3r9fAJvCi+3jCnWFh3Ycf0ji9x+FCkN8s8HemyQRkQubmUNZr77TxX
PrvA+z5jJ143MfYCcMxm9PLmw6Ws2+MHKV4pWMLlcUWUBlVjL9znfZok3XI445hh
nInAPpnCpoVDmcV5THfVGfuz3FyOcp856RslHU5uXB3g+fbf8xv7QIZbnWcpMVx6
SHUBvhEkM84wkdNozBNmuaWqzNeibd3YdQabzz68RA/Og0sHxTpwaKghT0tWW440
LKZLi8NokWjXhOfNF+Qy2LZAodHWhP18Wtq+B4KIzxdbIRlXqdniHL9CcJnxBWJs
HPAUupT4XJcJtBdl8UNrj+hRbNsBnrwgaybDnMc4TIQdG+DiQ9SFaXvq+/EVq3KS
NiufI3BYiIObwzm951P9Me7Jmv0eWQYzT80Pbqk3dUO0bFlUauEqB+w8LfeY9dZZ
0AIcNIBLChkulyT6TX+KYkrzlRyhxTnyNcEtCI/J7V1KAw1Ww1mL17vNkQnJ3UvS
rl8NTeQ/tKR+U7MFRzxk92qSNQ2BC5xBtVH/t67zCueXz0PJnoW/Fuos/sCNG0Ha
w+POpZm9J5pxnSDnWQi8GszS9xKinTZLOv1EF5HnYswAcUdq02eiXjel4AcfjmJA
O0hupvvrenMDUsOmlZfc7kcucVeqi8+xMDPwQ2ecBnr59rZ8mCPP8cQ+Kvgbmv8V
MEBHW+hm64x9pZmBma7ZDHnLQxB5BnpFBxxWNlU2KmmIsXiMxS/PoxEQzAD9yFty
1a0/dH682KDJYBffhkbp0ZqYBBdo8YSIE29mQ21tyINj3rwmMTlEqckOo/85VFvX
VLJpsfDxw4vgRZl7TKTBSXc+KHDztqgcB6pfDQrZVy/9l+Zm2nI2MTsrOX8Ak3X7
o6HuftZCmTt1LSh8lxGDQ8/sAKEKGBWWaW7Z6nJAsJiNuWH8iLvWYFOIfkP4ohhb
s33NolOrA/gTYaYao46pHHStkfk9Uet7ni7ObO+/O3VMSKZ3mTj9PWIDns/h1Jx3
asr/tj44tngWolU4eOkhhZ78MlX8IYoRt0atGt3XRj8B6glFF0F+ljvWFdFuhZXt
xL90uXOcDbf31fNA1Ba7d6/sTyKEbv7wjW2J3jLLAUgucGePAJlfOFosvL4hGLX1
4NbEYeH70ri+9QODy+6zedJd8zu8bnw2e8kXpwBPbFCb5UOOPEP3HCqBzJ/Y/Qwx
JRDRiN7H4v3CWnraY7f5FH+vrYydHjsU/bXdS/nRjqoVrenXonJ48qinYvoXkjjr
jP05UnCJZvue23/GFCaSzWOM+iwTuLCnXGzYVZSFG3f0DMNfPaAkMh+wZTSsiJIA
So9waOuFgUFC8oQGrAYUfb9EugdikOTijyBWQTZF+WT/iimnZJry54nhpJTVLNYk
wzru7EYbDHmPg+9Z7uHAPdqw+FYR/sXSiN5MKKblEDj4eSyv/0nGD8wwMLkYVxR5
IuO5G7Fj80xH0qdgSSIqlcG8fGZkOyE/iE9dJfPP6YE6Bq3+05dk3HYHrx4nGhZ9
SazE2y4XYGpbqDKZumHrGzPhnU51oZHpnfTJVXMpBOVZTSo3F/7wAffC+osj9l+/
FElQr0jw3CUWyNEMJS5r15QjkLCA2iTOjgLOLGvlwEQ4BrNyd/5QXryLJG2vNrgR
+k+hwvnECI1jEtRbBO3DJS8wTejNdof5Hcb3sxLBMv9SKrTh8pFD3CbQX4xZmYjQ
WOgHrAqRdnQ1JazhmjBMN1dEOW8UL3GrrloiMPSxw4vE10z+9Lxc/qlMdPgsag+F
nAbqlx5DOWOy6mZIHKYY8TSM1rD0xXf9+eBKT4w0HdJwgGHGskvVJOOAyluJKBr9
xtgxOabI7OvuJb3Cwqln2mwKYZDwIvZWLn5MvABN7DVu/6TK3zcckWTO/o6zoW1o
MGq4ebvuThfZ+IDHdv5jECu73oBjl7SYDvJ+evrJx5tx/ukMYp2sMfTt39dT/zsS
xgxT2zyI8cyyL6PNIzXtYHxSnPhs1DOsKcyktr0AXBo9fSALDiP28djoPBorZNgb
rz4CyJPE6mu+4oxUegyKMt8aYk9fpu/s5val6+ZGE/Z/Tgj65zTPfFecDQnfaIlT
m0z5ZgiQAgm24wRHTFeWYz+xoJIpWo9wZrJ3yhUQtZhnebiF3XbKHTulbpYvu1vK
6yzLknmPxXkgaeCu9T+pzgW1ChOECkzl0KaU9rHOwAvbnQBu88uRTz8pRh/usUH/
OuGxZqeXSlbd6XGMvETgHkw+F21sZO1//GFg3M451sLmXayUGUrsYx6jkG6Atpjo
yAjYwd0/ACc2A93cA3Npb0XOY5UFLS64kd1g1z4zOCvPudvcGv499GVGPumNWf0S
VxtYSKjsNwAOIgP427RTLygr9ySXmGPgK7cm6y5Rs9iVky3BsxVGoqZRHiZqPgnZ
6cenVEPG4mlRPjm7LaHCPLlWn+GMVlpeyCLdqw7J1Hh8aNWxdA8LwncrDYqUXO9w
pa7lKJYWu7/UKcOw/Sb7PgwUNlxLRkenAmdIu3vDrt70YTspYr8amSxt2MI932cw
WVbaqeLz0NekpmMNw6Sklr91fMYZUYrWWfUZlvwWnIx+aAktijlOvsrGBeoM73Nw
e+hB9H5sVdkKQcCXeuUd5H/IO6Iz8tEkMT7qCt300ww+Ez1efRVRutvV9uQXi/Dn
AzPOFmORTN/NdbEulUCcjmokQbSDXWcg5kEdDs9P/er/q88S8E5eYqGlpsnMlBvL
12ot0RP337dhOxgk8CSrXjR16+Hj17cZNbCNzccRtPimrYpAFukS5G8wuwI9gOi3
0HJ/RbL099uNHxyUYqx1kib4EWUPP7dSRgIRnhS7hkLrxRJEVXcMiLrSw7pvHN5p
9odElcN+JAJnYfifkz3EdxT1TJSaGdfzrCr0t7p9HRnM4d6U7E1J8y19E5R9Ay18
x27IvbDFN4qLRlepRDSrL54Pj92EGmHeCDYp1YXFd66hVWpCbVtvsOs2i46TadQZ
OcRLdZI4YhsahbVcdvGbygEdC89z1isJn9F/m/R3j7Z2j1N/gVP8E5VBvXueqgks
E+7whVSNKp5AmEpvowaPbclBTe0ceFjoYOJlh3SgPM5pfGJsr1gKCt9TsdSPWKgG
XdYcOnUM6Hhho69Xo8Znk6nP/9sjxPkMBZd+ePF0p4Ltzk555KYPyb+6HIZVxMsI
Ial4f4/CPRHsdLLAhtlyDdh75AefBlKeJSJBVgfVRGevKJARNDFLf2r0WGUVVKhI
tPE/X9dSVg/oxpIASS9O1pGnq4Vxx9vmhDDJymlX5waIfO8VwNLpdqx1Pcb93pUB
Jns7I75wmMcp9LLT/wD/tw1Y8Djyn1lOw1e3kjas4OpawHxjUN1799ksUdrD8rrQ
hj8yjSlEhpLBW6CEJEwBzSn5FCyukSM3dbA03eqJIh6bo5bIF5pkaw6oraa9ULgn
sMwJrvTnxgr/Gv7DaiZw+6icb2yNBIPHhoTH2qsR3zfUfaddgZG2Q2Z0y8ALlpmy
BnQkHsiUuamstXDhjfxaMRV1X/l/Z9IIZj8LGOzzb8R6+V4xT4+T6B7odiWnhh+4
+y6LLseQR8EfDWAvFpKehcPcWYihdSm/OwW/ferTfB8LLLKqu63u3UaIUeEticNC
iOWiudo4hADLv3NPXn1oIKfDvMkb40duASV8g9MvhEpI2/izXTzPjSH1yzPfrXuR
WyGhFmQAE2EgbmMpFp1l1w/ncXgxZ+LJGxP83o04GGETwwhQ0b0fjGpECpcGLzin
peIQw/Qlepf/tG0aS1RUKE++1DUq1eS3c35eN6oWzAStMpjpfYTD1qrbj1sqybks
8KP1SqPW6/wZBRim0m86FK6tTBSuqCTiDpRHXUEvhkDuyR1vsLmM1MeVpQ7CC3TK
3v9fYsgGavnNfHIO5nO3LXT3D4e++wDNInpeeFDqDPyUTY+xE0p3GqiGv0Fn0uDp
O6L9/Sm/73r/+D+V4DcaLNF2BLOfEMtquGYru6RjMdHPrZiLo3K3QKpCpL+kvexj
GD7kC9FOX6Nd+G4mBf08PxENTcbbIbZJ1JF+4PXzpvWtbTqr6oPddMb58f0GcZNp
/rpuAwq617/DzF5McEGEtYrcekUb4Xznf3enf5VmV9sQh8MIqvGidRlCMhh45Xo2
4TDP9FVzFZlrgY+Xt9Dm1svMAvtI6HbDGY9yL+MIhiWs21dedu4YacNzXmpNhJV8
5vp0auQHsrVlFSHWZWvdmwvMB3DUI0DWgR+eZWNAcjbHZmqSQNRqtWpIjXPMmIv5
JhCqZbP9MLJ/C/BNs4FXkahfrltG8O9BrtvMPmMJtVbMHv3+/MDQ8s+Y9XNGm+YQ
TWY8NrvK2DWOzLQI2fjqCqhixdpTjnKgQs+Em64hv2vJuqgegFP0xpOoeY2lbNcF
aokSnFbTCo1c51ZOX9y1gjixlucO/A8Pdsks2JV53nqSVv4ax++FgUfW9/G8nN5j
rXJGTHmgWIl6MmEd+HmKxGS8fHFgpHhh2dJFe8L21SYORKo7Pi7GE4+r91NNzARV
HLqLvlVqSBYfx0QpR7qxFpL5SZuVY7JK2r+IUC/YXsdYZ37ipZ7+e4IAqC7/6AnA
BK+ImvOn0zfh+QO3eqwsFBrIGYWiyboD8WWYlvE7tr3GRftwF1wHDxrfT+yYwv6O
UMfobAm3ZbkAY6+48JlgIhhIXhDflC9+jGM6e7KU3tXshD3Y0N5s9OGqKirtaQMF
X9g2Wj7+9IkV/dkcM4RwwYGap2iSvD5RopexV4BOgS2pp6qSiUGbvvfxcnpQWcSv
AetzH0xJpv5Fn5UbYrKFYjQyCeVlOZ+CFnOeh2QDZ9f20JCGQauMk3nZ/t/EnP7P
Ap3FsVOjEEjjW+BEOwXM7ANmrTi5i6PPP3gT0eaFQMQv/VOjVTAosMTdR15iMHZp
EMxNuFJ/J9BdNZJWL2CEvIITAHmFSxp6fCVP8pjpc74wXK4fxN2FAuWCp+qD78py
g80+jLyEwtFGgWtcIkj733a6KI3FMj0y8ylHvWgwj1eF2p9xoKLHjtJ0ab1W8pMY
IvgdmOloDP46Qpuhqr2/5BO1ypnLkRJDmXgCr42/Kj1Lab4S+rIzadWDCK3k8t4I
9Z6gsuEJg1FXK8mWjdV97B2YbXJ4aIQHrnlGDo5iAl79bC3LCDCtGVRgJoWofhIC
WROB0IvraKqwIWFsQsXMyJnBn3+4YGXWSwWYH9+SeuGT5K69oLgI7tKnFiH/b5ho
rB7hGUE5FbcYSDAZwxEFlEe8ru+jlWzdZRYRzYLV4msuq2RFowDDhxIBOP5GaTAN
OTJgXbo23QtxEg3JSR/iKZKaaLGLPLTV2oA0VoOrNF4X6uHsvpICCRMHvpx0mxDW
QL7llK7reqiB477Hj70ZoRdjBUAOB4pB2mk/cWkiMFJhtRuRBa7AQZOVRo69g3g3
xE8nCKPvx6AcTvUX49JrY/CRvAccnNoAaKrQq2EwK9zh57snN/Y+n67x9u4z16of
d1ZQ+LRzgN8hGeWjZTB/AOqZr6WSp2vrugv1hUsadWxyoKFkTuDrRAA/kBUadh3J
LuFb7+s55b9QLDWNpjVPA+0q079NExg58X8WHf8cClaNB58r/0Xntb2kAfMFoqFo
jS8SuHpRkrRcYlhc6sZE1lzYYTLDaGTBaY1SRgJaRMU6aeNXwCLZZiV4G+TMxm9R
GW5gG4QVSmckLJsbKIOuZZownT0dK4C03PJVppNn2T6zSFjVGiKDB0H4v2FuFoyD
v6X4yyNLvrg8UIbnSLkYZv3qaQqHw2SssocN5I0/iC4ZQClsrQfs7RRmAB3ry5na
YbmvJqAZV7YipXMLaLyfNLgBz5eER/OyBaP49J3dYQd0qcMjCISXR/O6nf1E5MGX
t9LcSztHj6vIpWFamw2ZWYQnvOmztnPYIjUkCgPVM/V4X0EXr8Ik8MMJA3kbDza+
+cvL6dsMYTBQtAZUKTL/Fx5vu0FFaS1T8M3UyPNxvLe0xgcl2zxhQguf4ggtHIrZ
uonWCv8uvR8A+L31pLRkiySepIR9kVZUflqSuZENSpaOGIpzaNzo1afvDMYVgntx
561jHbS0YMM7ngutT2nBZCc/aS0YuxPiX02c5fir7/rSAF6rGyGfDD8FIc9mc3l8
qycluB2esUsE9DA6549VrbiRUB1c/vZpOWc9SBGPTAij9kO5C4lY02SdtoV9Vnmm
yJNklxjCiUFxtLmIHTvTT/Vhi9feI8g9CVoLqD6VnkxHR0GdYaaQw00r1YLxqAi5
4aZ+WNBAO9tD20UclsUzkHZFUw0sjV1KHn3Sc3VAukWstOPY63xZnBDIOQRz+Hcn
0HkG8exoCV/xxYihcdhGzG5jBHr3f7nd3P8KBLYuvGs+jtjF/4MWNYS/BQwlXj+b
7mUJyS2k3TNA/xTwCQwVWg2HEbW+vC9IKDiKE5Ganfy1WSo/mnjWdqgoHmYyiKM6
Wh3gKpQ9gB8t570n6dPs0Y10Q1WArolSU8rsFuBSlbs+k90ED3I262qtcIMAACBi
siNAJh6G2KbkJj5XlbJ9LUV2mVXdvTM7htlGc/rb7w22RhV8oiokumsVg4jH3VRn
Ne3DEqbjQmba1CYjFJ62fKHZ0I419oMA8rligYjpDQ3m1PetE+Xb+NWncIyChww7
etrfgilkVaRomrMrjSl36/1cxcR91nnExYt5aLKtS/an//u3yqS7Lpe3YBSABh15
bjOEN/diaH7ewobULS4JxUAuXxTTVAmZgx+dFFyXQHH9BVJNM3AWZMFwMM0+Conb
epAu57UoL8L9mq8QkCPGqkBeuDyF2mmlqgA/TI9oVDwDKpkWyE2rfq5NZGEr3gPP
Bf1xhJO9/eST/Kxy9nERCNM/2lnRO9eMqb7qJPISd3s3kcK6pn+6JXo8nnKWhC9p
Ez8QBCcJNNkW9veHdviza/xeVkXd3LgMq7nk7C/4zyA8a0CH7/pEl8eKa7Kx0ZjZ
CRqLDuGGSO6lJEZl3CL+XQduHSz9oAEMe3bdJi+dx1YVdCABSlx98gzBgXuWZ+Ll
zNet7q8wk5PVMOebAaIKOG36YJscwnh/jTCmYL8rdu9Q/vuixjOteyD4+JrTO4Vu
rPWzQ3E3u9+ZJ8xqFURIOjIzHmbXbonHN4zYdy+D5XchNPPjL8thJB+m5TzVov9R
J8b9vv39HN7th34W8/lcdl20GxS/rqu3hQ7yQ3c4m7Y3KmNqdIPKBfJw2nfiV6XV
ZFTYBgqESvatvq9/WVgGTFDg8BCixs3LPvxfGfZv6Qc/trvwUJe168lWGDONGW/j
h7Jr6zEKaeIw3cEtaOP+z3kB2NDJcDWl62vcFve5/qKZ5pvHGFRaroW6ZWSfvPCO
h3Lp09xx91DOzUq0XGujbVoRFIDmCr/hbxWuevuzQ8USb1KYQCYyv4ZiI6murk9H
EJBkPPfdc8rR3R2b/AUoU8ySNX+9wJvxAQ0aNMckdXWrzqCbY5DiKL2zyx1Gbmch
`protect END_PROTECTED

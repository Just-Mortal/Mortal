`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FmviMAK8ZkQEir9ZYSr5SVKiZ1NRHgUzvqDsW9PGOnVazQfQhXbePZCrx9cJBzo
XJq9SXD9D7+KZ7QlDzY3I4ZzeBjNPb18aw1KeEzDpYfL91x1yqNc7aJdHFeyaLj0
hDwUDWgd6eKGr+oJ+fYf9npQnjE5bUnuVYTmbh01TRww1eNZWQEXjBSY87L0keYl
DJBiR0fyrkq3Ucv+80mFEEYC01Y17FA2uhaFpFp1FD9RhlnxwCGhCJ1Nimsoybu4
ZAx69QlPZ015Gf1kYsF+GnSjeqB3eIZnj0/KP/hBDH39qypOGDnTMZrVqxbw8GyY
QaAqgSPZL/8P3VaXJq2ygZQOAED5dD61M0cvapEwGeDiAeTiKyAZxmPQ+yBJ6frV
N4qXsJViRvEzzMtUDVaVyowTyasMYn++oEHTmUfu321l1PPcJ+uqO58LYeFK3561
yRHuCJtcNmNzrwrTv4xiqWvMpjMTYnTHHx+Bq3mmbH1fqV9lHbPxO2nbesPRfzXq
WMFPp8c5yAQoisCqPzPMRqXa3ula7zPxWIV2gkkJRMu49lfrsCpzX2tVeD07zLpo
8otPVK4DxVYVXbdoDIvKZ44JS5I5L/TA/EWNS9fSqI2RxSKoMDfs3QBAhNuTq09s
uQD5aflwk0bBjP1KjMFtUrj164tLPD1Glcax0+X43PeZSsaO09+5GB2pqIuJh71L
eoa2ARjr/vkY3WlPYBJSbeCsLSol609B9g0CCcMDmhhMeZ+1a6RBxqwYhUAIb1AX
/Jqm44IDFoya2jKN+Km/WFH4N/ShncJxLBXbPsJaFvFeWl2H+n0Bysr8ZTBiLj2X
HUHoM+7F1Um7DJVNV/rgng==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
soCGSrZxjCKDieS7uBNoeCRc+XXcn/KyNF/mRFp9VJrMw/dYwgXYOyUbsOyUs64B
BNZHs21lLcHDEg5cLEJJiC7Dt0CzK8lilAHH+Hh6mqMF59WLkWNfpjWRyq/+8vtq
YEKhbrwjzBtaTMOpAF2gJ6Vg/1UCrr43RF+cBOiCYXK7Y9eflbhScQOlFlm62u1R
b8R6FxsY6gzz2Csml5AQ1Oo+Kjhp0kTHPxXgI/WZ4vvb+R60WnpnfXPjO1uiPxyG
6YJb0484MkXK4nKJbMbE5ruivaNP8SSmgO29fzDRMe92Q8FtM3hJlZnEaKqnKnfB
n4wnvn96SJPItLamPtAJDHk9lCK6Wkuqu2hUaWSDyqISdR82Mg3oKdGDm1PDb13x
vfRHB/yIR6u2IJbnPmHkEEGVnA/K7oOtpCYo6zGmtHF1ke5mS0+szAUzTa08K0NB
YHaPC7fLZobm3ioUu3lmi1ugXGjNV4B8/rYvVftyuHc4S7F1EzUem5uzYY16dw5t
eb9wcRcmQEYMV8fdQROIerNAPIrJYxihjf5IYhtSdKmxT08Hp6ytV4V+d2BLuGeh
OQLi1llQGRBJeg6/h2XevmwzXIM0/7oI81xVU9bN9REO56Mctki6RCQDqK9xueVP
uK0Dz7PpSznu5SSg1Q/bOa/aQSDSy+nwy4olsC/bCxNnaX3Q8yojNIihkNbbpFkQ
YR4t7RfsMRHY3SBM4ATmCr7Few1gQXG+QiNZQMTNh0tC4PMCVDj3N9eTuLgVmnmK
M6HLjJy2a+684F2Ur9H+J0Jg2SjkmOaWIGIOspghxwz/SUlS/1UdcaRyNomD+FFO
NpuqDONgbxq3xtGOZTiO5ux3TtA9cNhfZtXhaTtilLBAhIZbF2P4/J16Ci/uvJpd
ArJ+zVDSTrQ4Iu9/c0KYe4fje/1RpJ025s2oPSCj/oIISP7Q/CwaT0MPpUruiBTb
NfS3SlAriL/tkBVEdTdq6EolxzieWpz4PY9Se72UWMMoWhkyETKfFfVyIpi8nSyg
HyQ1Mt8y/ThxvblJlKF2lXtwVSKXKzhwstbZc80qeGy6omHHBHJts/4yUojjhnyR
b5giawEN4n1t+CREj3xKr+a/KpMKC9wq2H5X/zhr/HgKwkSXCBp7/rXJ4/7oYHh9
w/MZuTJYB7M4S+WTdqgaQo0RG5exo2eMZ4qo7KHSjkJpnuCahz1l/qXLVcKxDzCw
7QSXQUgEvgUbZlE5TJXvyO3dwgEDNNb4FNW/3iXn/qSctOZl2QEIBrpEz/H7sjx9
SBfvLodKA8LuwJI0bEyFuvT4oq8hDe+f4cQSg8th3vWLYufA2RFs7ncxET+0Z0Cm
ij6WGvXwt/HsBYpjh6GeeAviprRMOqId2GtDEqjIgOCXUzzCJyTm1mRKAGQBgN9f
PUuPYyAxd1txviTkQASSA/8Jru6Wyc/esndjE122Eq+y2ROKOVORb9XccryZ+H4D
6zNQl4qYBeAnqLhoQr6g6m1Zv90Q+QI4VFpXTuDqgbnL10oGQyzejLdMX3l9XfmH
/AvRHcLSHn08ies4MOCtYS11loPYbh5fjCj0FuxYqY6j2J7qiupGy4iRW6EYaP72
+N0T8mjTWLvQZls0ajrYHqMJkVC9JXSLuWDT8u3fbvQ0kD1/aY4Ny1b3Wo+FflTI
2q/iR6xU1Xo6H81QO0bzCbSuB5pGKKT/+1KyJfTiuVmPwa8CzJm12ymkjzbW/iAS
P5B8UVz9GwkUIWsBIOtGQ4PLiDjI/M8zPtTopXmi9QzoOnNSAjbCCG9RhBNDu80h
ykx1tbHSNPUWmEhMtnK/NsYLuGXN60xFuipRujWhGbV02kFTnf8+6yecEE22sw4x
qMWEwVHJpsBJ+s9EMChhdqXVJ7lrFJm4zpacCiONGqUGZ+H7gaiLXOIATTz7WMcU
LTAa2B7X3DwtUPKBy5CXKkQd4t4FIs7DF/t8NZO0AohocjhjHI1KmQKlk1vLiWHS
/Xz3xm7TFFEIgOGd+Z+GGXb/qE+zKg1hFxSunl70stzCiwOtfJb8NMw8+6uTogGx
mXhPuaoTpeENClHUwe1F8AWxtlM7dxbLDlO66C5tCCwCRcU2XAfSspRN/1T8QmXz
Ax83t0wg7DAVOZyEpyHkDLZJbJaBL95nuNUGhnNrcrlEXzqUpq4mfzJSeXiPUpV9
pn1Wlj7oFgRWfzST++GD0Q3Uow77owZ19aKGAs/OMo/tryYL7dowRSYOhVypbJxb
rNq/rGmmerKKQ7CwnaBgUcx9zn2TSH8AkunbWr+fxlxuvZ8b1K1xJdcrPkgHgMaX
XoucRphMzBCtPbi2f4uqsbID36c8U4hlLyGSiFj293oPC6lXb3FhlkzWy9Gfe2QN
iJN048uqofqqcUNJlKMXHixHu1pj3GzRqGZAMW8ilCdiAfNN0BSU99TuAF75T83U
sF8IWpvf8jyLWpSezApbH1pip78y1wdKraJmR2ABEzs2IWF6bkyBE8MLkO/o4vLS
MB8Ub2IEF64mSpRdZZzJq9/2kfAe43bfn3uizgPTB3bPeSII+LDT98+UmtpWdwVP
gS5P2SPYCqOzyFKDxdknK9V3giHXsyu4WH7Rc/c4ECMeI/qmKIApMLm9k9pw90OY
HrLpvBkiSB+KjeFOJXxzVRCe9MzQDr+ZGmNLqE/SJT9Or1Zr0ZOvy3gDiUVnLiNx
sqiF/KNjOWMFFajwFlsg0alSyjOBTjOe2yJvtMlzzYrnofDGyZ3o62KE5cRwoVhz
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ooNxgDYPsj6J3y2ssOH2ClA/rP4ffTbeAqMKIuHgoTD/H12Y9cJGvPEmBJdbcqiH
KVF568i/CuwqrEJho+UAtkWTSy64+8gtWbCmacbQ0rHZ/LWjYQ4ee1NExqxQUcPf
LhWg2ZCacNHd7kTO48GDOtgwRNrgKLZ9Xwi/xiAZPfdUIpn00Uae27Kk5WVA2MPR
l9LoVJLZhzDgzgN4VCfgL731aICIvi9qQh8eV8Ru1JhE006qIS9/q8mTIfh4AYVa
Pt9NzgF/wgIhKJfKB/fEQAmE2Con4PX3QX4ajDHAQzFwzoUlYI0yHf4u0Yx5kHi0
C938IBigVS6QAsCejZ+TZTXxnlzjYH6QbH/lZIMo6BRf/HX/FGHNF8corVinUfIT
W2UXiQT6aj8lCxo59ykt5CHDUS3YsdARnafa4ydG4Pv6nTJVUsw0vtt/XW5+x+EQ
dtzYMvJKZHEmnd351OBN8IShavkx7rexWWpU6Y23GRKlyWs5kMfCbsN8leuRDblm
v8bZkl0JlZ95G+3h8FEIS6uCBACMuBo6Jod18PzD/u49+Gg1lftjbj0cTmjPj695
MOQ5fmIpHYjDfK4XfWTTwiRA+Yz/y5A32JIfW3WnSGlITNleFWYOPUtKnEkyiCJL
8Tnp6FiOxL/2m8sIyBtMccDYrDbBBsQjxSS+tCpVZ5erk5tEOtnNQhY1QfDBIR2A
hl0iRvZDdbNhAZcft4nIA3L8mPH925rd6aXRgO0oZyx0DDSIyfp6EekmJjUCGsiO
g8+yUSTAovLomWIhD1w/oCSra7qtriC0DsruXN8IM5ohhyup78t2iWin1BlfZTv9
hYyxb9APKnxFJQV0LM2bCC0FNl7JscKP73AHzhiik1+9rF260m/ybZRv+z/qz6WT
OX93OFQofUrPa4PjSBfiLsbMH60Sz+mcouoaZwH57MTBLnBZfbKxtIi96zz55T7q
Q+IYUuEOIUmwOmyUnWr4CbfEq5i2+pEjb2U27LaS4dveCKynE/9lrHqE9uHgM7rL
T6sq2lNh4XL2oW2AQKxbFfr0DSwlttr9hfnhAUDHmpNUxzqAiRBCN3OgIhpv9aMr
y3XEW6emr0vInw5z6lR8Ew33djgWYqx8Y7+37+BjOQjez1WMV2BOkIycqPE5zIWj
47zaAvYez+/bdlV4kkvMafQGj3+EF5gY8aM6oopJMG8nfX4dynhqwD5hRaLf4zp7
v51Du6Au23o4xOavocwlnjo3Y1t0c7teBun1rivyxU99OpOeS153zI3iRTIsyvGB
mjaLi+eS0da93sFfiiiiT24aRYY+lU+WvcyYV9HeY7L59fAiEUB+iF22VjdU8oKk
HY9ATM55galseAgqbNzUQx4LB+2V/vECHi7AVKrGSyxNwqUr+phHWa+Z1krPBChE
htWnL21ZW5LTibwmnmKZ1pyX4wN7en2Rcz5R77aunB26D8OycZN+NeapU01LiTrz
0NwdsVbkOjenHg8dD/aEBwLWSEhxDUWXnLD8qMSkAVMF+qlgr552o+NjeqVJMEZV
PsBphBXrJz+TIziOBZ756837fw3DGyA7LEX0a0IabVorSM0gEtmxCsK8FBhrqCUU
iwuOQZwgkjVSzuTlgy7EUgCcW5MTzp8gG4C/m26PfmuF9JLybX3tG3ZZoxYGBz8V
9B4ND2vaI4mIgxtc7yLB5GPmseaQfN0IU75pIzIzP+49uMXFSB4RMaPmbUfFBkS6
utqnJ7uTAcXAMuKjzwLwp8Pa/YmyAIBWqzmg/60naFWgGKwDHNYRQ53XCmkO5vT5
yXN3IradpOUX1mbVC5Wjq4Jgd3fWq0frmRyeOBR8uWd7UKBXr1PdKBS/AtpbJ77b
JdpJdpDpiyGI0fB/quk95A90gUTYI38nqeIj8pQFcwH7FqvEgc53DET/LDRnpipi
l6AbiqyeSMth9QCZcnhwYJbLZE1VBLhoQHMrFNWQmEl1lUujGv9/aXe9pKAE5DFo
BncQDYP58LIk71YOefsqp+axoEPi+95K0udCTGHj9bFK6Ulndrjxit1Eru0KpX35
A1LS8shkDE6DqNxLphk77puJfX+GTBJ6KSbM9hK8aGpjpxZkcIosbPNNGy468AD/
D7q6iijCOcPN3dleNDP0wwOl75G5awp4/9LQQMzHebTLg+LwCUgxpOWPB0rXzCPI
ZIQOr/yAVPIi4/M1iB9z46NEKfiRmdvPHzOJCIly5bDPs+rItjETUmlgb45EsGWu
YcFWm6d43nOnfTZ2FmfPLwpyXUd+IEG+NpFmtQQpeaVuBYl4gkn8LHkXBz8zq+EK
l/2DsotD4FSYSGpEazDiQ8lh3XpT5kXRjS4/IjaAj1g0Zuky2yQKHNwCnfxouFWM
KpKy1DnZwtm5QOAkcltZFzFrbOqsnTIfHef604cS54HIeqk8G61ChoB8P6DMaxe3
P3S1y3Q/SevShKNfbPDhFO8DdtPu+OsgH1uLiVuwIBQqpfHR5s2k03hdCD3U5R6U
5Lh7qTtm4NMX3JDKcc/3rWvWo5mtqpmJiAw14IHS6jU=
`protect END_PROTECTED

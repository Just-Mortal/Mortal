`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W5tfXdV1E6lR7wTjQu97yqMb58MNoPZyaAD5a3vgACq19DteadCcUStoKh4pgdKb
NpnrRm1BRPMTlt6s89WHv13ek8jC0okkoCPC/PYTs3K/7ZG0YOkhMX80Mqu5e7ER
ZI1ZD4zvUc4GMVYK9iq3SY0SvALzaAS3644b0ceVVwoWKknXVWNPQgXCleUw7XsI
6Mw5zazE3xFWZHc8gn+nwTnY87GlFhSZRwmjy06Gdx2U9wmq4yWuPDUJ9VGUNaPA
YiKq72VuHgmFZjiavdySkC4W066xW1poOlBRp6cs3eBZwxABeQ8MXU5Qu0kuT27R
pguLOwYx8Gnk0FNaXnZ2Y2ZK1hUW6+diEjLsHHB4bmCdXWHIPKl9re0RD70wq4OP
/UXd+PEsB/Bbl7/FlCkpYOClUEZUoTnqAlLgtrPLZE2ph4LryTS6zq+wpxpTIfy4
U/p40TCwysLzbYYBTb3wSFds/dxF6ahICYR9RRNGna8ss/W3HbVSbjDo3C1rvbDk
uLeg0hugK5YAvfknab9qC2aXZpgrl1fIavvhh9UbdggGJUjj8v41vnemlUvXhyqD
59cpoXnCHlzq25o7zLaK/paZdTAIcQvemgqFWwTDLlDGRmw8ZSS75iZVV4GOsm8v
BoVeSoB+T9ph3MGmUPZnM0tFWfCqjLcVefDQ5+uU0dGmR+oxbQ+mTmbOBCPwnlBd
r9TSoEv2NI5VEzlG5IPP4Y+HNv8/VUMY608McrClWlgZKXTAl5SgVEKIMO6hNwd3
TcX1A5iLDX5MYjzjl7iwHTEfJE+W7v/hyL3iPhehmIXRxnYZZXch9ZfFdjaNx7Is
v8zuO5MxcIybw9JQt6OiUJVYTIz7KtuYlsal+AoxIwMGNQgfPmZZbGJzUJGsmWOw
0CD6lOJJNgIhnDlEm/wQWle+CixlpZpKIOMWhE95gfzZQ7GD5utKS1nDvEQjXtH8
mOMXs2RvUcxrw/N8yw2GSQma3Z4jL9gazZGuDcYoTEWPc++huupwe6JWRW4dP/IW
/1DXcPgMVz6zbIrRgcQPbdsL0rvYGyGq6IOvRkd9gFxfHKXQ9tKjpBe8pbecMriB
rbxZ5qAlOO9fPt1LgeY+uhF4B1G3Cy1fms38gBbXhQDLmxHESwQ/GebKxUfOEOxe
91o/qeWlA1/e9KVKMJio7ANAgMTp1M2f2qL8DiibbhCh0AtpoTwf/EZQFmePDLJF
vTWeS5e1RcXR3NMKlSwJZEk25wfQh1q391SwiNzCe9t0E4ftYsAKDgH7u9Upbu/7
6WoK84IMhR/W07tutncQlc6u2IjqhAKGPGzFPfqyc+DNISIrF7W6Ocoz0fMmhLMq
L/G2HbDRYGVB0yg8phdHEajHM2abVcst3lzGccO164BQCfmKMNyvZBK1KxN4cA5k
0E/+NjxMHlhcMpQMLOwNHU7228WduhKq6de7RWH9kHyEVH5RdwaGyXhp7HdYCnvJ
8MF8dKIJHNDxqzGrSVejwH42k0Oi4dT4CeIa8iLn696zUzQaBP2biYGOWtuV85Rq
jIxkND9sGLfb3xSwBRTnB9KAcySm4hRJe7v4iNJ5IWiEtUv5hAumtWaAa8ax6IaC
lvulygY3pePWILcETCb0A1nwkE5L+3/ckiy7bSc2Jf9+0ArbVKZcrSc+taUJKLsh
+srLqrA7GnIKwsE01qcbiD+djypTkB0SZsK0LIMTTifZ+P2a6smJdxMgH/yvMErY
MbrT8vFaAB+XLosqd+3Nu7uYricraZaSPVbwPU1swyJzpPhf6oIlfOuhEq1541md
G//x9HXOLwuYusOg6EBd05kRvDq44e8WF9MiDId0kG1beB/aTTTFnOF60OvxtzAS
l9qZP5WVgNGuZ9BxOZuYAEJNu+szcu+/dn1htoxup+FtXEBKtXspy0opG17abQ/u
aUA2fHKGulVuiNXt4X4h7Xz/u9WPjLvg44Az6Yda3b1IZTf6VDhjvKRyAxRa2hCb
+YwQxTBAQB7j+mOxxjn0aptb4lYhSMWY1RdCI5VPGpv1dUp5gvaM2Jxj6c5vB6CA
6Nn/18XpusMk4WwJyevo4xyRGppsV+FtrqTjKrLPt8F3RfBwWWRA7A3Wz6ZJ2RtK
fY5O0r0b9+WNQUm493gH52od6PcFsUEkEftuAsv6IzDP1oPy6ZR6RE4NenEzNxWC
71OJQula9LGvYWGUYAO03OZ3XAlmPsjQZ7zU+4kRxBDng5cUeCsB5d/spSRq0xsO
XD3BOMlnPb1nwzH0uRn8GyxE1TMI8BIfgbxPkjGP7pXAMLNDDpGdOqPI4+dhLcUG
GIHZep62UXzxsQYeTw+x4pPdzsgrqOUUTanbTgr9UO4x0KHD6Iq1QlBy+lCQghQA
ikR3pN1tuWqGH39xvPPWVNOUvpXPz/LMsONYVB+PkDBJxE7IFMGnFthrQK0Rs0H3
Fl0D9vg7HgnDZooWodZkBFtsXN5Yi2dGjENsTs2CR9Ezfq63HsRpGRiluIsFKGo6
obnfRpOig5B2MbUdz5qEWU6bAmbBblsVAmZy2KTQe3chv2qlN5mcbNndqF1nwQH7
aqQ1VZXF9Yuu8xwqGFLX7xtAromlr4sPkFAN5CbHOYCQ6Jy+jNdW+TBaMZugHU72
H2HrdU8axsjaIeKZeYn5I6yEhYetgtlDZZG7H0HwwH96ZWNvom1K1j9OOJxkxXwh
GqsUblpZAZhsDQNYtQXdogein1QUvVnQwCk7jV7UoOKunnljZb5Yy1d2rtCE+YmL
6KBX4MzbCNGGJjAJmISvdk308qr0Qbd7qYFncJntz9WSi8o+oGBDt2YzSpcE1EI1
rzGWbsCtKYe+lXaO/SKeIloymKFWU5vCI+rVTef7ZCNGewlZLqKe4A94K1DL/7ju
kexXUlI05a8D1vGcHDvZZ8zzXlIXiZSj69+rNSSHy0qBNaZxfI72sxlFCoaeRD56
BuqnNjfKPHl9KbOTCzbBQ6e9tnBf3I3bI1BpuE3BnsQ6EwgChkQaoaec1PCjzt2R
4JCeNN/3WvXH63xDRTSjxCPpmjVLsh193TZFkaH1UMGqLEtyli5piIyjRFcpMTew
ELEjN+/6ZYo7DFhqiwfnAXQ4983e1allDZnmlu6bie8I61k1AT3fTxFtJgfkqQUG
tT64T1cGHq0GfEwhQW96eMLcRtK+NuK8NSmkExV5mnRuNiGppNwzGhQCrmP5OxEL
hDgHXqazNh7bmRRz0fYMqtDnzwuYQzqLl1fHOxSUtocl464x3McceZNhXqjEJY3c
XszTiAALjYHz1ZLM2eBsb2RcKuY30f2d2613I4ZvpjYzk0FLf++3GUsA7iWnswV+
rJ3NXXEkbR8ApMXrt2jSnYNoLKaAs6iseyhpSr0SyRIkw/7HxzVpT9ZZvf72ei1L
NmWmxDSS3lKSgMGX73ps3yC4+d4CGsKKY9z6YfsTXLkIfMBo8QA5TppaWUepWTvx
DeXSmEtvcr1RSNyLS2lX58jrMHrAfznxpMyti9twdm//8qC81Znw3CF0UhFfc6uL
WhQ8t7xJj2WyNECNJw25UleiWFNDEWjY9Ar5p74fMzqrFK4vY1byljKwzRXekvX8
csqi3FRjWpOv21gBOzihDTYMIjPFVDDfccbwJqq+naVTqNjUSfFOUVsxPJXtyMRu
4Vaqwkf8l8Zcc+27d/Lewn/9nHZuM7R8JsiXeN1MNGkXh2Mbs7zDQmMOYiC98B4H
1rwlB/GxAcLuCu6s7eVfuHJ5T7mnPnMyT8gp66Klog8YuhadNNV/DZR2aACPRkL8
Ab94GxRakeVR6xmH1KfaHYTTcZ6SpgMIg3B8XEoJRw3VWBVS5pZbOHYsKQoBkZ7X
l25V/rLrx7hraLCzvEWW4AwvLhyuywRNVJOnkLhytIttTR89MiH2Cg3OTyrGLmCT
dHiy1qx4iDjCcLiAFkOkxtYSXGCdCX9H7IQmYbg9cwKgZ8Hx/XEENaS7Q8a3Bd5I
JjNGUCHppBb8AH58JyoovSh/BJKRKO8pFqDFEmnZ80xG43EK3OT2dbC9eg/m/axR
sOhlUq4ZUnNr7J7B5A2pBxtl2+lVFVBDDW5P7t5xZJLGPLJlHt6RIsa2rFoa7OBe
O6+ixLNTfJJhvz+J1Ucen05QjHjfsHP34J7ta9MfZJCdGI6HbeVwf+CBk63sEpUo
D/3GcrXU4ZpQe3scOD3+78PyNxDXVuSmnv09zeF9KM+ARnk/y9Zr1ah5+fgImyqH
lKQxag7ivpglX0dzYrDIC3eKydz6InPasScOGfGDj3dFW3Qmpq75Ey2Oan3C/2XW
W9Ra16JTEJR6+uRlg72rM8z0fojNSTj1qn6gWd/JTkdFTdz61ZC+ISfvFW9yN5ne
7GVn+eqDAyX5hEYC9uM6WhbIMbWtqiTQbHP7CWMHr+44aC3JskJ/Z+wS3Ow1GjTi
0KV7SgjxornJSWlDVnR76vcVY+sIxgfXvZQfTD6UzQ6ZKUbl5VwtW2hyuPmqTbsK
2B2B2s5hpDMOS7exZzfCJcWKGqagGmGHaI+1barXVln7qYv1zeoSvcTbEcmA613c
Ah6n6JDmBqpgTH54smm1HTB3pkweEV8yhaLY4wpO80SIfYWelbLDck+Dj0Zj43bF
sI1PfQ3bSYmY5EboxCDxTD4OqlG9qU3u1RksZFNN4sXYEd1hRdhsxPQyboL8hgek
l4SLHbkJnCe9rPBqtGVOwB8a7AGb/baFeASQmFy2XzPW7K/D43sv4Dkhe6/c2sx3
NdNXLAkuiXn7wwbGdGrVhKGNfpAFbk+VKP29ZwUD8HqazE7p1oZY1StX4LHe38wM
hCWvKjeldqMMWWQ7+HcIsRU/8zmqun3m+A2j/+ZynBb+YcA6FmkPTg1noc/jetfL
2CBE5s12LiWmQZ76oYhW7M4vp53duOPnOOZUyFQ5C95DGX0FNgez8DY8CSfjgcvB
zz7dPbpfCy3WHLo4phQGZwa2dtJ1RxMeYMETd5xfH7wNNG1AQBGX8R6REXuGi3wU
5//n9rOC4uymgZEMIEsAaHimvoBx5FrsshIHZOymeWfLXH3MWzyLXnGuhtmN0hmF
Q3899mJjJAii5UgvUXutmwaWIJ+0JjTq9vgYjZQQ2jokHRqBnof3Rm4aGpP6lIJf
oDbXyemUjBDVq/Mt13QNbKSf54E5nm8ARDVr/BYZgeufztVdQFhsjI5jeDKgYFsP
2rpIy+VqKfEHj2gZpq9BLnWar5VfbEivR8cfXD2Nv3mWhCU6fF55kreFCHSGKdoC
NWPt1Hu5IMpbz9/+Bzcx9bE6VFVtY7Xu7AftqbtG/YBWuGke/cHLnz+/vJ4+eSri
3zU6pXwWO8MBEAm6/eXPf+0Op2+5n4e1XMEkoeYK7sJn6PXGlreg2e2qumzf3g+w
mU2yCaVE0Xoub1blYt0iJn/PkOyTsHHM3qbFWWfGOnefeM6L4gz0nsw7GS5TgmTZ
LrB6i1HP5oLV/yqzQsroZep3DxQFUvhtpWj0E+/rTWSvqmq7rLwemBAbmvXyDKPq
mX9qLaMuxzAGeR9HF9TVCjrdQpDREAqI6hzubLHwa87nJMfCY29VobT6wx0HCEGt
W+XylPaiTUsC0S2JbJJFy7lfLF0/oB9y39Xu9bYu7B2ZFRJYYVjoduS42Lj5R7C8
zFjvuqs4HShjt7CYINlM7bxNievOPS4vKFJeCMj3iL6PmhJqPG+h8iTpJ5oU12wh
rW1HIcvI/kswtsArVnyGZhLG0xcQcc6LISfng4Lb3JSDYs4v4ATMVg173fo3Ng6T
C/Ke1AJ3VBY0roCJKHnek7p0iGOqWQAiLqQtQSz6xwlboZ3QB+bXeEB0KwFHhlZt
8SAxiiQj7Qvpx84NaSdBtl2mgbbh5Bs2GfBSZs2/d08h80g/AKEgbRSkWo/rdjGT
mQn860GqqPzGESqNqAiaoWyD1rDo6Col8ZKFOux/BculuVsDx7StErj4S+7UMlIt
Ez8Xp6YNKEQfFz6spug5uKFQEdgI5bd4HmtMpoHcCHA=
`protect END_PROTECTED

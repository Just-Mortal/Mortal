`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9btUfe65KSTmh3W9VerwNVn5UX/O+SkPjKqVqV9mInEHYTNxWtM/wJh52/NZNya
IIrrlU4IwRnQ++v5yf94XOtObEcQZoEyXzlzo47069PnxTS3lQeGXTMe1t+aF7vk
ucfLdH11TALOYQdiQNdEZ5KW/PYkUFvEFRxMb7me1m2SLO5fSXnyahuBqi0xeZEu
5WxWZYUokMiu62WxLmsDljSaxRX2SSxMhLu6yKHaERfkeQg0mc5Sx4qloYUcwt0F
ktMeMRmaqnO6LO5y2CVhRXTehvdEmsAD6JgJ6zTcSbpY5ua1q92KDz6PLySIv+8j
3HY1wiuA1l2ZsOQxfOMvJBTS+GdSNavtk6oQ3R+G38QQl00OmjMeERlFrzoFrTue
SrcQ/Vpbe6b6JRJUSk40Nd/R7WYiuR7KYlBjjHPFCR+dySo/aYrziqjEhxeQXoxw
KftiJ0cspE/iMWY+Ro6tontaD9t/zdLLfePlwqZQ+B19B/wsIL3iWZdUS/EprHex
lHHZzBIfgac3YMBe95rA+m/CPdm01QYlNP2ld2Olr00BMmMENPWF97hShBKcdt3c
twG4ln6cNtINfYIfoszKdfPUAoX5OO1B7WM3gH0kYnqLBNNTgiiBMLeY4pWC28LW
XJ/zfufgph59iYQm4ohHxtgGG/Fdwl1BT2da2aNbb6SuD/g3F/+15vPDzfcifAzC
+1pj+00WAeHxYjteMka7GAHENBar2pA5NdeGaVvRzDLcfhqLMc5bGm69HqzsjiTN
Is48Yc32kM/IOkV53U1g9ozttn/VUldueSTFqxwHPmJzxDOr9H4576oXTETnSJhB
mDVagDfJhliHjKHalTGKuaMO8BDto1YiMkXT8VR/k3SMbjm7crLAmhVb3FTDMr0g
OoYtBA7m7fHm7t+jB716YbifyXEHhyDbtHZjHa/F+8sMmSPdY60r2HEJvkGe7xXW
i8ib+5EqNbnYGrw25hwcROK5CEVG6ZwtUMGTGchC87o9OxvOF7aQRXF+x++cJc4s
dVIXh/u64lJXrAKQaSOyBDww1zUoNVWCuhWelid4sm7t5bfC3c9Zc8NSaW/RmQxG
7IVN6/Ma+JAQWvgZESLgfd0fS3n6R/yP1KdMYg8oRUZJsDUn+L6ohvT4x+yZMDWf
T5KQnw8zaGgaBuji9D3ShQn8JCRb8A/c72VyMCqOQP+Mbtdfzdg5Wng0Bh1EQzif
tvTNiXrXwUv1FS4V92ss/HCLxxunp9pKXxDSjzO3QqVrY7Av9M+6u/ez3O5HDcMZ
uy99sEfTXxWSppNt63XellM9STkRNwzk5lBqwRlElgh1pmZjjAnhb6hty32OAcME
3kTRw9jaamwpdjUI9nAK8Eqlna0RYsWNz2wKdLmbp1Hm7XxxRYIHu4EbOvnKbuxq
kgg9gpxyqABLw2iJ7NkBAdQ0VDk475+oCHqyBm1eOLOBpfHIJYP8FpcU8lXZt/Vp
hSYBKSZQAzwF+m2TJVqqKS+KVDo0SohG9TlACSc2/hqJlNR2yQBI4w/W2J/dqUlA
agaYe9KNUGESjVe3PmerlF1WRY1XH2iXW92zFzWr+7IeiIwz4U0FWx2YFF6PIu5k
kijsw1VoPhnraAUH2TPd73BlHZrtmGL2+GtsRc1f8Hz8u6Q3jtLXtlFO4JaWc1U0
Rrt/x4S4FmDVLpynTHFa6dKquAHSKZyvhqQoXvOOF6QRsR10n90GZ8bReUWHDm70
lQUQhpf+iXN64RHTX73e3JniVCuNZCJP1VN0T76Q4r4F/4pv8U/d0M/vjBYjISZU
yI4WgBZ0u5CdL+NRNTmlZs7TwgC9IHIH7unJNWyTMJUp3G0SS44HfE/XcofxgyKl
grCONVtPjwFwfeWWvx7EmTtD6RjGpced8rlNLVyTQ5IqE3uIofMOtzold7P/femT
tusyaPsF/Sj3b5iOx7vijG65wDjxiV9EALZm4/RHKQuK84ep34iGjbRVJAEcJ9j3
bdZul7nb5iIs7+4yVvxMBdQ7h41zgoMGbVkCsZj6OBXWAHk8RANNnD14ydbLv5Au
w4FUi8neKxLolssXG98FN7LpT9Psdr2bfidoZHA4InqPRHCNOGDX4krMPsaOW5d5
Xyiskva19ngFZ+JhSCzzcw+X9yow6mVdDmAwb8N7ozTh0LwD1w86t5IeED6wMXBz
k2NA6FwM0cdBb5valfJQUGX28EZreIGgQUm7ayGDflHAd5yUOl47MiU8DhtCTt5k
LvI9ZD5wSkJrqd/tXY+mUptEc2xwTjAobXw4XJxklwMeNmO3IIIaU0HW/XFOtmyF
joka11rpVHD84OhA0e8/gnd7tBPNRRp8hAV9E9WqlPF3OyksvKty2xwAOTreDXE5
70F3iTABSgxLX0Zc0/frIT+/QnGC4QDAuZrNlBWgUItPg7knsu0kcmgGzX5WDAr8
VPfeFA9OXdpgrKES6DeOqG6GbmdK6uU6Ul1NgE5tiS+6dE5nyER045oZQ1YKFrn3
MofYu9x8h5xXVhqVEWF+bYr7Qj4M/KVUdv3ROe439X/T50scm8gG1MdZTvKamliJ
`protect END_PROTECTED

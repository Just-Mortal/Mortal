`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/O3c5UPVYj1yELfQ34OqwhIZFHIp9odhAXmR+yIGmJSEUUYggsOkG3jkir3zr6K
KOJJTmrliW4P75zVD+FZ/v5nGiy0Sbmw2AiSiB5I0KcQSquPjHnfyY4efoG69BFF
2DyK3+iA7AzlXILp3m6F3Ph8DpfAbnY1WI1d9Es5hf+EqQ4M+s5beLQjAqhEWoxL
J+Oc/dox3fwLShpWGakb028lfXYGZMdjU2LXjOc6jabHRq3NNZ28KdIXCo03bltR
W7DkDMEZ8KyAmW6MxRJrm6nnYv3dJiEzAENvnWPRGtVF7eh714IznWrmHDpVLbi0
frEzpgdMkV0lXmJAKJpoh2gt7IRzjNHPGfWbS/n8SwktfANFwGMKWSU5RJxajNHr
WjsKXlN+2V7LOWj9wM8w3oHfL+LoXD7yXF8Qew8f/VaB+LfjSKqbOv+CUzH1NGix
RUWX9duyvggNf5bQGM3hsiKTFkN5MorL6+IR4RQO1NjrTu4nUnSUWMuoDp5H9tWP
uxJXojCmraPaHsoKDydyk/t2SrQlIKX6EcUmnHbQRbGYk0NiN0qMffiriknlHVFv
Y40mH2vVRuz1l94vRskIOjhYEP96uVuKUa5/CXZIiN6E/LNamF+e0cUEgLA/QjPT
tBp1XulAx7qNO8LtrEiCGoQeSQ43q3YWglChALCpSWsG4fURRS7EVNSEuVBOqoFq
x0Xy8pplEDEMkoXXmr62KuPX9eo3MAm5Z1u/IxvijMcL7zT6gnCOo2W8fCuO52VU
fZX12D1G0F9LqbwFUvGR+V9MWSGy1vDwjnU9HE1idoduBlOQMri6/LmHzB/CMuo1
Yjy27Sb252jAiyVuSSaBho6IBVN+1lCxfMXnT4TkFygb/9S8DpTlNGjpwIkox7wZ
Txny9a+Kw+8nQ0Qof5dZ7BqcbCnOcPPxkxA2Dw8J4f9E8eo+qOADmPoJ1eMzVGlw
s28KjNTDmdaddrF77XXgfno/7hDo5fvfoLqL928tpt0M1uuq34uggzfIasOUwIms
b9XmEuXyiTgq+IP0t+iq/24aZlu6I2rQ1VjkA4QqmRcqJU8S9OEYFmzvygHZmJq8
j/dV7byQ34azzuoljpVrTdwVb3wIczX6YHE8CnZnaXX0ENi1+3Cw4Ym2GsWnoN5z
UHyyJoKzac2AoMWKawst1EgJkenhb2IcCrZ/BVqi3K7/ZxWsPEeSwZCvHqAbsXF5
ti9Pq/rWlpGHpVA9b0f202V0XlGbOcjQwwtg8FBgtQlmAHiGMr/QlrpFlaVBClqo
jbcKx1CvG2/fRizOn/MKfGwx0j8gS6B5xOApqvB+Fdh2RRbqAy9qN1WasVICjrY+
Xp42QpoIR49FZyjv3Tw2l8/XtW6btx2PUBHfU5wE8k9S6gHAPb3Wyhe8sOXfm/zr
gtQiJXb1DlK076rWxmDuJEeWF0LiLVGtZFSfuJfEp2YgJ8kBP73aalB1kU5bQsSB
yAh0Vc4cvgLRUTN8CEBRYFAE95qYaYfWg9NN56a3ocTd9IfQaXVvr5qmu5V/wucw
MCComP2U0ePtTkq70WauwryPlH3CQ//zm6Zvu7iktthqQ76KKQaIxZhvS6wTAHvp
9k/mKCqLB8cbHe9J+KUg9iAO9RBU8lVAUrCCHj1B60Ndx//8b2KdKhob8o/259ay
SfZDMFBC9RQ/py+wxPMbDVHulqTnQeb4eiTbXUbBIAidBMoWfC0AuSgjwy2CBL58
QjtD5/AGyXvZeWtD+JWc6OszsY1pdF34QA+ZjSgrXRsAtshfOoZRagFr80Xnt0qO
sTcPT9UYzmmML48qBHdWFoxJaUD/kZNn9E+JDe/l1kusrVU9sxWvSwQcxtloKiaX
pQjZGpGUGc6VhUInoRdMS1o5sGd8JRLyvzFBvtvK1nFMe+RNagN71qEwh6Mg4TPl
/Utk1SIVGhbvaik6TTIkCIuTDp7XeBNJTvz+QTZbKYw9TPQH/mVwWSL1JLvhv+WE
x1yQpwYfFSrn+XOT4nB163FwW6dem6XPINrJZFhCg5ylKYeBwO+iOANS3kLFaxZt
wBJH8w11MyqILGimFlCCfBCJwalkyjqk8ZKTKcI/vjox4OwCsarqcJoNnPRz/cj6
O3svNGG1KQle7tynO/CxvWpaVfkI6GlVPZZGoJc/a555lT0jTp5pLjt8ahfxeoBq
WqfV5VHF1tU371BswjzZBnmlS8tpjFE7LR7u7DKDpjulnfeyJ5O3FqyDHxpzH1ia
F6M/ZxKIGClKUZJHe6inUMPzjSg611LmYI3Aoi3gjdbeXbMF3x0qCu5HIcAkcNaU
llqmCGrsSklA0z8phaOKlju9laL2X0vnGcB10ZiSJY4D9ZWGlMXtowsA6FaSMcMs
3qNDwP2svf/+KVMtOpDA2R3mTUuG7QwApUmJOvoqIAaenGpiw+gyCk0uyC2nzkEa
zYbwszmGwTrbo07q1q8zCg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FznYKicEdRls3qqkAtz7y7gAPvhp6r9dxosZ6IBIicH4E5Cn38MW11aX+bPffGPD
2kSIuX3S/NYJV0vDDXoIg9U7HplDBoUE+sCOzRs4RBY6PuGPLfvFvm6UukR1m7Lj
VdkiRLJfIbSaY1A8OUTkTXoLE/abYJtYQa9owsu/E6Pb7hJm/9XPMJ7hgXX36LJ+
JgiisKXqIuETMIRX5FMNWRsOVhFYtyNE2euqROmFCHaGG8SzAQ+6fjDJ7EflzoZt
MfHn7etmtV8zPfKGQoR4ckMzW4C8OpJ0orw2cs/H5IgCEU/NZM9GtfMU9mDdWHqC
N+tIIAn99+R9ARwdLhQr5Bkmq5FuOVX7LwcbKjocdk+C4sCoEvEGMK7c0WwgpaXk
i4UkYGChCBY97ThqX8D/Bjm0KYtgaW1qoa+8JUM0/MKLLrMGjnAsWcPlYq/1lzfv
TRBtiLsJnmBz+fEP8+XecLURlru5ClO8h7S+AyudvFzv8mcZXnynl6m9ibH3EAFu
soaILWqAsjAF1bG+RdvNMbv4Artp/cG4fBaAcXBP9B66rFGsmU5N/OQREJ4NTdXl
9pvmJowg1fO50A3Yjh/YyKD/5htOeIU9g/IE2Ky4ugBRksv1e2Adjw3J+An/KdSg
NEa/63Lde7TXePcPX6j3eao0G2rYxOjgIwU4WEMYi08cc72VaIwttZcu6rw1C9yi
P3SPuLQ8sOKakBjGXZvDVWNWigW6RAiZD4yl6ssAa7JE4eqWtpU8042OKWgkKfeD
Epxj/SJ1rM4ui34fq60x2LO5SKmPanuAPn0QjXa2smBF+L62VqSvSbdvaLO96bNB
j1mvRKNUdZSdWaIxZmGXbQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5GAgd8ROBXfRS2AeDlBW7EjzC6jEX5jQtLmkc0FbfzcN2mN2IcrLGUW8dMkzzjPV
4fjhNjVHd3l/AdSVUgrq76t5PiMR268rMFHRUBpoe2fhzcPVKlFdXtogWF56vs+/
5HICfQnMN6XD+yvyuh6+KlbCqwN2kxkT4r7ttOz1KbxYSfjD2EL4Bt7XpNGmwqpd
ntcebxpDwejs2jn0GQXiZfQs7PmgADDkCHam6bJ5lKJbutNnX2+mnJIbZg8QABr9
elMJ0+8t3m9zHGH20y0Gv8DCrd98YbGZxwrGPj4KLxJBf3yPZXzljkTjnr7NPAkl
3u1yJRV6F+5BQcEGlCO1ZOgcHuGGP5r5M0P4Rti1bPMwbEp7LZlZWSkeU59Qvol1
0rr9MNQzQ+H9D+ai41mzR8C7UFgj0I+yZJjt9QQsdS1o4NU/1ZtQjewsi6sduFe2
JOlEFm/GB2NIo83DwwsYgJyabjQSh7BF58G7Uk7Zj7iIabZvESl/uipcTPnW91xm
mTo0BKdBlluicIkHCZEEdISMZAwcb+WDQ9j6oDJsLgGewUd2XGqokncL+XI2omdj
0bWBdQ8X1EgNAFbWKuuc7PcMkEa7QwFkkgASEHCwbSEKXyQS61AAfhI41k7WIZOt
60VYTWSbDOlqlZNvjHr0ai+m1bkdlICu6P42WdbBh2oORcIpSeKOoWCOTZsi56nd
sB4UfBU+vblK36fFaf2BGoH1lUDEebZAcGq/9Gw1SjqNCZpEK1M88PwGA5NJT3S5
RYPr3O7H2qsVqNyx6mY575PR3kVbmKyf+OO9INrEYg36v2XJFAifwiQG1sizLfsY
FTKAeJb1tDia1vlAGj3AYpw3706lCl9b7Hb6EZoM6IMKMse9MbIx+2Aeao5uA8kl
9ehdyGyfwAeq286og6Jjxhn8nv7vDcjnIMG6xsoHPH308Q2mecL4rh2vYzvG1ev6
ns0gSVf3er7ffqav2PXAp6e9wlH2vqfmyplNwn9+nHH4dzEyMu6T4xQKq349Jp5+
ey627FCz6gW1YnXaLfXpshSeWn5ZDkVCY8nhyYHqeW7cqTmZS3laAxzz73PqP9yO
mb4O9zHQaxpoKZZJdqw3mHhgO5FXxaIKIByIh1HMlQnQ86vTMMeAfAdt5lq5uqGf
Zpbvu7EXiCj3mFvbBNvRCtdpfVWkTBibF2F7NjQEKuA3zcPC1EUHtM350/0ozr2u
7D5Dy6HSYZrXZ7y4o0DDI9uu1z/tZo4MjsbhVL+aDXJBWfcCySvQ70INUT6Br1wL
IOMxy3m6TFLKv8Z+SG6lXvy3p184JXuInSJdd4B9xpmmrTtZGknyw9Ni2R+mu1mT
Rh9lERZEeniVlZ35afh9mHFPSFWcQLjBQhE1YNApWyAp+oOUQ8G+S+ujt/O6ljb4
OVB3zRnZ2noOdt2qJ5eit1QT0KR9gO9z8aikkkP18ytLj7VUexF/ERXrPbQZzchW
blERsg4vx8auQJLKNTb3sYkShi5gzD3fsBxDQAdeEFUwl2x9MG+8xBfRZFtfL1OV
yXwJEB82qrFLykWkcxX1c3eFwhUapOJzWykM+xpDIFU/epwfftvoVjoKnGrOsfgN
mqh8NFLqcLGf3u2sW9+Vztq105LY09yAtAO0Tz6b3YljIv7X9YUXa61W/01FSQzB
MADKlxBH2g3yhIDsx5qNX+KBjwoNGJXRgJWkqNjltgXMKAgbHspnjKjJoxe495Ow
NCZ1v+i7cC4TBttUb9zbI1jL5FX4gm3G2nmAlmnvNR8mD0rfX7W3q6woG6SSwnlf
Xizaw1NIQzo+TnX1BToVrTrgBPt2hK38tAA7u9NhBKCqWOp7Hqz7fOots6gFuS20
+C1YcplNpFJSmOO4Sfj7TYh6iF9Dttqxkb7Zz9RpOvF7PSSs+MTusePGWyhBoEKL
iuDp4TDPm6mENxhlnlGZjncbDhJCKLHJ2uNB/dgiEgIhHEGOT/QvCJ4NS65qoIVn
L36RXvmmxv5AiGM5iMFSHWc9LcoV1ylK3weFmeW4CXqugPNlx4ETkNjRm6DpiVz+
AZe5Nn6fxJ+sHimsfiDTA6CB6hiYS8u9ygV+3ZqZyYfAbrLdk08LzaC+03m1pWrR
fIl/A3wg2lkAdOvnnMnZ3/aXZE5WPz2osmUAe8Kd2nSzGH1OqDCOlB8sofnw+lA5
8ijhNN9aQjJb7IwguI0f1KMaNVNjQJwPhrKdj4r5vbP66cWQZmEwWpZ1tlOj0EZg
RJg4w9Rq+8xuM/eVPrCRitvf0ItedAECSMhrlhridL87fHu0gYmllqNP1aWFZ2tU
7PnmqlqYMKGLu1PFft7HkIEmT5K3k8pyADLJZBJvMhomJA5HT4E0XJR6q/b3uWFh
upAeYc6+Xn+3cybytUQAg5o3OnuRhyIZmjY4HJ8xGs04J99olegPja26bKNrkCVz
2EcM91oj/ymzhObGQRB/54gefY6ZhJPs46FLMFKGD8R5tgjUCKP7bPwyyaWRUATC
gjN+2t1su3Hd0KLmCzuK6wQHzcByGHlvbZq+ok4kT9lJee2yH3oakZox58JYfXcy
T6xAlUHp4XMDOyIYhMmrl5nC0/9LGp86DTY0t0JnOgQeKzoa0FE3OW5iU5qKDODQ
c7Tn+j8YzGvgBAZzQ8vu/dQSYTMrLeECiM1ilfRjRE5Wkn4Hv33ZbJ3nFBH+31UJ
2VnCzfdrP0TV7XmbK/DBOADGenT9/J33Vag2UI+wrvST5BeXP3R6sVcwy0cvKyeb
iDyi4Sd9HeqErRhJ1H2iJ8gmJ4S8w8JNW6lzsv15hmrshs7A+eRQGnyBkgS1W97S
XLze4FeScrGfpDyGJPWwjFxdu1GgqJ+SDnl5zLywCR5Bd/yEnPUgYeVFeEP3lzL2
Do7bV6dLLU2oaRSosHwxZA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sv3WHvetygzdAworkikIZXXBh5vAl3BSR1oKdoTdvCpY0rh5Xp5VKWSI6yp+oDUF
DSv04VapzsS+vei8O9kS+7zT68Gw+5+Rw1NVcoVf6X2EPMp1UZSi8O0V7ruwmgn5
g60klC65m6bqo6T4WDLVd82cBQnFDI00bz18VYVb7qZbolz2UZuV7z4M5vATSdvO
id8JlvrKEu7k4APU0ZqIn/TS5VVGaXiWFApZigPQ3grRRT3s1nF/GCpKDg0T9PEN
/8bdGLdTQ/2e98/SSqYqrhtOMZseo/blOg+Q6gjrMP106eiPkLQrwbgvharp2f8o
ZTTC+NWg14v2VB6d3L4pOugGFxYKISaEK0AaajslKUSPblK+FPTgvew3DIJvVVRk
ddx6FG7+nK/rmx4BkNfniPbMilSbQjqqGT9a+j7MDgTAwqjU2ryaTbZBhecuUu44
QxryQk1/cg5g5cr7r8PnwRGQKcVlDVT9Qb9SPuMERiB7W6HbMRjvobnlAc2SPGmL
vNi+Cy1rCE85K87dE8tC/EGXtz9X5EVqsaccmPcRgSHz2SdM26rClHnNPiR/TkBU
z8abQqkRrhnyvs+FfoToJLBsxJb0X2ALrdbG5yA32IphJKK8Er6SIWZp4UYRONIi
1EgZyXdLVwolTZD7P+5yWC2JiLIizc7GQLio5/MTzL1hmHZg4/DKy4QNP83WO4U9
8aGmqtXrWl5BkYNndeWxyuI8XAdFcze7CR8p46fx3uOWpJVHe1cteceyJMNtva/L
wIrmisTPoOXJRZ1OV+nZP5U/5EZ69hZoyUYrHH+7gxT04sNkUEOnDGV9tXuMJkPu
wWoKnIRCU64WpJV6O3ZPvD8Z3G6Z0orXscR4ywf7LGFnmfRmrpehErEGmEvjXNpu
3JhXNd6/GMHHzyasEYF1GGcAs7gBpsVzb4iSo30PGEQviAwPXlFqic/coWOAMrct
Z9jNXq4N/IfeeLSS91IgxEyLZJrbLnH1M2074vrMqOCOXxixqBWC4iE/FH18o8+x
4FliA62I0fxVRE5nUR5bnI4pzpKFfmA6eOLyvFhEBCbOlvwwJsOvER5lGAGGNwVH
E+R/SbIWOO4xO/3CpC5h5upjMrYsKPkMuyy8Faced8Ms8WWKO7YORUhFRdv6pi9A
YAN/CO+LZkDw8174CYo/hAQ3ElFfCj9v1ahzrI+iUK0Xmz/peJYFooc9J4YLz/SC
LMt6aEpEez2l6JA1wNwSPVw9xEXEzc4OyXS5ehgz81QtcbWYzlrmC+aX2cbDU/8P
xe3xZ5DjEa4NpYUjkMosJ7uWxoyvFsjde3Vc7mdvC1HrqLa0t51hVY00Uqof3KHK
IGY/U0NmgwOAUt8stYJPiQ3VYfnQtAydzenCLJ8ljhz+PltIOozH3hYjQsgtTBby
pENHB4Xcf+T5yN59woXmQpAO+0KITqrSD306WXNxlwfKl/XbtH0APAZ2ooeQ6spv
tKJX5Iv67PHPg4J0vSfktLsPYPc2M1twDFuEEt0D7Rq1kU08pOw20QenQK9O3N1T
uW8Yuakjv36gf2AboPC75ADVU7w88mmNSfO8YIuoz03w3xfrVcXySpqirY4LURE+
JQCn2koIMC4Z31xzZmWKR3N1hwlAxgko2OIYPY/SgobgUHfJDBqoK0EPyzLu4+5Q
StlA4nsBsorvoa9X4tYjXEoIibI01BeyxAJFD+mBvQ3r+VBZuP+vVPJVhyf6qiTt
1W3iI6Mik3gG73+LZLYg+NYEYM1NVh5bD7o1kvsvoEUaJzXBdDJ6ToQ/YovCeVv2
SFaREOuObk3ZYJb0YM78ZqHbKnjFJwqyrwmSeT+yayXCcLPym0CfOhlMf8cYbgml
YHgaTtZzq3yoGnuknQjxeC2k1bJtPEO1OcUUUxdJog/Y/hk2sYkEFytSKcc46QCT
V0XVqNuP4JzqAkjnmfP5q2c/XV6+T7/6vIw3xrT/owmq/3Pfex4+oTwWBrRNIy48
LFIPaXhyc+FR7AruOip8c7z+hOf4HO1JWr1A1AN8O2PRiSdhAuRcIVj1U1qGK/fY
IymaWCC/7ENtznFmFCuFCHvtf4LTmpwkcanTQ3Cs51t+P99M7komRBZm8ni7qtr7
TpKBLG4rbV8YOE7x2oP+gDMstvAFFMkk6gX/DoyjEaWtDuYPTZokJwxk2XP5pIn6
+y8j/jwsP6EzJVBTS1IIV6Gx9JaBFS5Y5x89ijQWi9YkgXiQ8VYXTxRUercw6zAa
QpuuNjHRzXVZ+Ku3gooX7LTqdGg93gtODhUN04oipbLaRH+5iblZ2lUMIXmR3IwI
EQt4KZr0KsNeAhFn+BgOwpq5u5r58PmlhQpvxwSB+6AEsq1ckILvnG1lhPcPLKHh
/t99NZxLC2OhM5X0/8dbLQoVMqTPOJlocJpFt6ItYKfi5HNeHr/5UcTNAcDQCQhm
wSA4x+Y1jOXKWz2OHxPMk5sQ0ccTg/HYed26Cdlo0LBIqC74nONS01xxoc3VXoiR
nRE5IRABNbRxofAbfP80opIwDRO2uATqy6FJ9f8Xv6/dJsE2kMw5ntbuRb/Prx49
FUXVK1rZWqMiR9r8pn5QVq97fGfHqFC/NFHSBvAlZwuC7IWP7AZuMeQcUFPKvWJc
OxTjeDtSn+U4UDzFxxDSD6lfEHq/vZ4lX44/RVoLXCpkZva7JQXJWR9qcIjcTuyn
xFNwE8WB8OvQoeiMM9E97JE1JH7zskrYQUaCI9dzEAyAWoYb+WrKGCvoNq4skv47
sn3QR6qjszmcoynqIFKFM0zdN+HBkKKLjTL/wMW7wlMF1Za2Vy7kDc+pteO+KpC4
pd6Bl+l6wHZBxJEHm9uUD7ttvPoLuo6s6PLdVSvfS2bX3DA4FX9VN96eIRkTIqSn
7z+/f72aEVnAEYUY3DWbbfXHpQAogrzNv22DpbllGIYR3ykMWO2ERhor1YMfIsC2
JXZnT2dj6VsGeg/Lq0ikg3Kdhw83HrslZFpXbwmy5kt2eIIfVGldFJjtS8w1rLjc
o03lGkgLiXifNsCCdH6queb3TvEy0eDbmKvRDv552fM+7WIoU6sIxcxWraDdpITk
WTC+NOECMoabPpwKCRx6OyIxiPX2EZB5IDMA5h/sm1+o7ZSRtdNHwKeNODwvaNlF
+V6xUgosTxqRY61ChlDlvWdsAcVNg6gXPm+VpLTygX2g94E8zutxocTpW+atUYgD
NqmQB38cWE+DSCQEhhpan9BnGt53xcFNLgvYY9DyHDRbU4HKsqb+7p1rD1FT2uV7
je5PuY8L1jZNWKd4h1cwmMp8H+V+h76F9x450EwIurprwNtTNQmRaXiZzUn6Ngl/
pOLPYbjQ2a9650UWDNAysL1b4CwBDwrgcZTA3kM+pE1c86VZsdZXtQDrdfvfGOEc
clCOaFzzX76ZlzUmRPICMrulxWaShFMbZq7Z2FclByQkKXaKWs4mLNw/yemY0sGL
79xQtK9mWfi4b06Gddkm5vcRUn4GhfNJTniSF+5aUPXcQnXGHhTY7pO58/SjjErX
E2VfwZ6AwIiptmO05ysLVYb9vt2RDRsK/IWQELE5Eu4jhw/7u5b4sIaKp+o/yvyQ
MlR+nz2J96OG2AZ0czLQRy5RygOsJ8Rrk1KHQAXO39cZ3M4yiSNXWjwvMa3Fw3Qv
8O7W6E17579puJyxpRehfWEz9E+htlreLS64NriavDQjEnDjpItug+OpCpRzZfKe
PAxlJpPt5hjpm1Rce6MTXR29tt93x+ph+tPSkogbVEmKQ8F9H9h659D2m2tRBTmf
vavgBmUsQ6bYjHnve4G1exIwI6eorotmOmsfViHBoTtFF+9wsg5GzdNv/tjjmR06
w6Dqzd47DMRa443iczq+EUyIeeTFKcZkelIbqDz1N0r3O1ZZd4jmxtz1UTXp/7mA
Kf6KbnPb8K5OY72Pk/N51+yvSq1PQbqOFioYEnqpvDrMzwd1AT1amhYabTJUOXbe
EPntztOz8umt0RFDC/Yp162WMdonL4QmIjyIXLCJhahYId+/F2wNCApV6EZ5VhUq
ozWCIjbEqK0o9MkZYeqIyvx69cFWkxg+8LfDr62Lq2TXt5sIrJRXj4hg9fUlzYvA
xzhN2h1NER/1Qxm7GD0W+o5a+geTuA7LX51Ky6+XghmgHkmbH7/GfRNqX/6VL0Jh
L2GIL2/ifiSvpbm2kIRRd4MoieTpouAnn+RXNLLWShywR2bFVxqozBNDPaSNpFdw
G7/YFEvtdPJNSRBw/eQLLrb7ZFNmHjQoKLU41mnpwdU2k2Mf7k2kBGC45tFOp2jg
sI96xYClcgAkt3uGuTopOEzYt+3tto/BlXNnPcA6h3PrqXqMQ/lphccHr7DA0SBL
IVBM3G0GULwDGdNZXmPTKNpVz+MKGsi4Ql6Q8Z8ODH0UsotghJ6EnclMPE8M/dx+
7+Zrj3UtAbdMgtdDB04IY4v7sB7J1Xiw13OKExZcw/0vYDYA3kiGjnUFG8tjvO9t
tfsb2M+v5qNwVNsQMXatfTaka/PabUzPpM2YriAdbV8YwRva+IFNTvROVUUZFilv
UL2pKGfx5+tE+bt2S6oClZhjoFASq9TqXnVnTKSojUeDlJEuO6e+NNAfUHWMgRNu
O4iN49GyVZwxl3eye5Uvn+TiGdfbJ5jtZs40L8NHYM4gOeMzKRpK/ufjFPty92nT
GGoDubpWCyS1GvINqt+giphrSvp8819MFrT0O1EG+sMytGMLmuVlMa/XkxXMzHbb
L5vh023O4t6cE29nUt5MS3fcFSUTcnL7CQ7B/rhlwwwIW6DxONwQjtb4BokNk2pz
rI3Y0psAGKL+ZJ+g4ptZ25QnFytlL0d/deAtOBFXXrT2ED1/cCRoTUwCosT2iwEG
xhX6o7aTlsGKGj20/dRppWA/rRCYTyHcS1kZ6kupvGrPy/CVeQX5rrNvGsq2Woqr
Q1lRoP0hBtZ8WQbvQrXut3pvN8WTe1gGf/7t/YqFsl91ETcrmRz3RKPBEifFwBDB
A6qb4pVbgDgmn5lBM0yPT2Ha4LLtrD6QidcQkeoqB+B/S5FJjjCDU91esHueCSgU
TGNsuw0cfayvcnEVpYZcRwd4AWBDEfHpDkJCbuMDBmvfwhBW08BFgzBPhToVjp4J
CrcRVNfcL9z5WbUoQrKeq4qrPzYspR9lsCxOYy6+fzzTFSfkgny8yyZcCHScq8nQ
Ep+Cx5tCoJsyrbGWjE4F3J5JsWv5gZ4PmQ5bSD0WguVtIPEPFRiy0D6WzA6bRu7h
BF8mKtvJJtPpTr4CauPzQUYpfH+93UfOAG4xgEx/z+MMVwKNKMkAa05QZphhysgG
b509Yc83LW2fQM7rZz3nu+UNWZLT4CPbmEm4NU6dk7bSicOik9yuBNO8TXbY2dol
3sj/9hKwLjMw6Bf+9tEntAOfwwJ+WUhhQ+eJ1V01aSAwpenr9BurqyQsza1y7LvS
XIJc5oC5fRkqHvIGlkYvr+qLragWjF1G0/8PsdOBaG2w0O6Lv+0fOfhRTL+ST06D
CYn/DBGRGN379yVStMyjZYzmdzg3aocMOHlTx3uP/99eJLoD3dBwbdzDcClzK7lx
v+vyyMMP2w4rUtQZf/iP+ryeVK1kRTs/XkzBq/TgTxLS4XoYVAu0zf9lB4GySo1/
C3D6iMCeirtBbHsEncQcSFO428g3cqAUmOeeNM8UqtnrBg6m7+OJ4+ZTEsvvpX8C
nxcyTdk+6odrPb8gmp414DDu+6I8s15CmuS3awtbT7p9sL6oDIpr6Fm1FTaM9Kld
prbIPEkqannxlZHxq9f1WIIvTVUkr3G2Q2ZgH9BHbySugCsKI3dUy2IPCgGXtHwi
FFZiFwG+8qllRa94l2D9D1hdu4ahGpUriNQiGl0EV+AE+QLD3gQ2O1FwSSa+j5Tq
i70CGAvrr0j0LZrXqCPbC691PuGyGfuaKsJSeCV+WpABnAHoxjWNiAlJPaAi+QAB
5KeFx0VeB1u2I9vH+jg/KVlugRn6c3eLS9ArGo9iJ0P6lWMAA8t9HB9K/Krn9T2X
qjUBdk62xdMi/1rZxBTyk9z22AxHxkD43UizqG1dJrAJONloRzLVgA3nlA3rSKB8
nAqR3BdTe8Kqzd+S3B722t1Zp+w7SzSMaMspMKOw+DPwO4nurlKJP+RCZUFQmocT
C6gkK4gt112GmsI5tG1MzgO8R4uolIg0i+QzYdJX9E3qYty40nUMJl3uePTIVxEi
UpHEkiKwkk85mafc+QlNFAjIrSISWdsjk8qDH/oomh1a/ejWB6rqTNCb4Bs0klwY
hQDyxTu3xgGT0wQme/HwFUP369IQJANFdQP3HqoR8xNhVAoqr1/qyrpelNh8inmD
yEXyPfaLJ23wHD9BvqucQAByT5uvEfbpTK3a2lCNLIeBk2kCad9CkpW1Jzq2XWJ7
Zr34lSIndxVZ/8nnclvsn6Lcwu+ThrNQJDAowvYdEdR7y7g8aAKoP1nRE6qlmc06
8Ql4PwMGkNp0kmkFqym6IGkldajKYtFREVoEjnBp/yahX5GPrNCq5DSX3uiwoWRi
dRCZ+1T1Pr4u8H5YtZ9sE1D62OafaVjqtk3wF1O0iY38DXMh48Rggmzhucdg8tRR
5+Qxsjwfj1romG4mM8bXXhY8w0PNeQjuaIxK4xDk0MKb8No+jOfXt2VHoWC0AbnR
3aIvTnoTYvBMEq91kMQM/CGnGAPCj69aJ5FcWikX+ZpSSsIGAuSmT2P/60BsfWK7
VjGGslitg849L+Xazk+kXJx/+sLrOaPohPwvU68yz/kJeJtFVCVesWIATnmMYPKn
XjQp5fxTMEk7BsLrUtRSo3SzGNGrygzF3t6r++O1v1fnG+qMR4VbrW971aomzdXS
KNBWrND9FJLQ9yRWfhrxuHTAa5CtiQzCpHI2ljXhnv5vq79RvNchWmv8jcXO74o5
csLCYLx2xoJR6xqZtxYZkjOiAaZdGzjwbEF8DduYftpEdlkUOnZZunBI+7AOKIkL
`protect END_PROTECTED

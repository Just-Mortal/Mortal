`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fx2ziSHwVa/w8Jo1zrJGESVvfRNRjTcldIvIF6WTElGHQLaRsW40H0vw/La+aM3S
dbcm4lIjrY2hBqN5ubhDss/A7XROw/k0w4SRSliYhrhVnUMgzQFc8DumHRrxSg8Z
rBAOtARKf5mOA/CxLpw35Rq6MAan3gFX5LNQvsj38tEkWBNhG3v7yyHBqzlaTrGK
CqzQ5JIX0TV+7r7yk9a09NLZqbcfk3pst1tYG732gVAAW5GatCcb+a79GFEudFQA
snDDdTgfeNbb8IplJU0MdFBQsExod/DjuYvXxvZio+ovjwLmiYoCN/vk0BsTt7m9
2Tw/Jc0Jy4wsE9cL3UfMXjW30xZl46sCTwOHB7V5wRcBY6rvjU6QRPddZtpqfRcB
eH6DZiaAc9kZdcb8Id9tiSJUsbKvWGTLsFjaA3KGapWpd+XimagDKsNX5FItUqqV
XPtCIDDlOIe2+xyCzuOgnaHZUWIJ3j/XhdKGtAfgFKPTtGNF0BIty3shRlIuPR1t
jZ6lPODVHNgox76JDUHBjiJDEMApivrCBQs72Mhv45Ty9CJuO2nmhxYqkGfPuwFu
PG7QNtMVD3y1b0QY3u+OcULURFwwMp2GVORMMRgQKWFGxaSix5plC0RbifcgMpql
2LAhXP0jZJxXZCaZhOu9IJGRg8M2gquip7JmYnHB8GJvcDoUNe5J8N30lqE7wtRz
RnN2OtrNxHAwerJSDmejmXyzHzSh/+zlOMVTF28/TRHSNZsFK5pNgnHjkWQSUivU
CoDKYiH1ofITzMCUj18YGG6dzxK/Lr9imBmu1xf8Z/DbR8uCbTBRq7bqTwjaaJm5
Ynt03VwY3xiFnBdYgn5IfRsEdfg4T2g7xgkFuH75zqujnJchp/y+p3JT8AnUx6Cu
YbJj/pN+l8O29vPvGSLvuZd96Pqf8x2UuDtQsX/91I4ElJJ6Tm6crlKmF6mZ5DG9
B/k59LbhiBZGW6f6OdOj7xTjFN6wfV3QUFoiKiKJ61rh/+KGFOAbcWVDRPClZeVw
1OD00k56hAb3vvP6kHhs4uekm0pYlkA0jYRrxUd0QQ1uQCZLU9rsAAAJYKF+sC12
H6a5egumZLiDvkgVjb81tQDEHk6KPlYCZgExEQZTcbv7NX7NoifsOQdJn/Oy1Ymg
Yq23YyULHHJR+oi5S/r1OE0hDys2MHxlTrfYvWWy3+1wL9sVDvuDIoija1XMG/Ws
GCiZIfIsGhblV/7ZOHbjxm4CqixZxmmBndCTOjINVaG5jnv8k/sOjkYm4D8bPCzm
8kPcb3g/MeiH8YB2WubiWk8/AT0o8YniH1Nzs9BpuHTRI6RVguz5DwUbnzQ16PvR
CqaoCccz76+4kJ7Nkxl5Y9bdRK9w9HuQqAS6qebEYYYyjnrmijFtayczfVFoH8nt
AW8ZzpB5r7CXIJRiILpr/g==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXgyTyAqZzulJUQAC9r9aRPvoopa0weMCZCXFRlYQ0AJYQoKd2PtJ6810CTR1Zr0
MJGkW6zJD+N2bpYfKOv9p+rM6yN2jQdhNVP93cjNSdi2T5uYIyrEII/gw9b19rzK
58y4H2o++/FLyfMLCMJS0Qy3G/qxrDziZvXgWFpUUBbpo7h+ehFaDozHBw0FoPie
C/3SwNy5OA6vaM8Pc98A+/pXMnHWv/T1i8G8JRRPUtjwS+/99/bOspJvrJOd5r/x
jvLvH71RFWrsXbo9qLgjfFInyrVj1X8zhWXlEngIcKcQ2JzfAK26whuTV3VZNB1J
+ChSrR5eQDjiWmNm8GQQbxSUM8tbCg64uAWAhv+r8zF/3bmWjhn1ag1q1ZZoM1xa
QA0DnjkIkcm8795KUeSfwLs/Tv6lRjaZ5kyFHUrOzxz2qogzz/Uz0dvg9tHEs5Mn
L6nz5LEygyb1MprBagGSn8m2BRU0y+2C1W+f2R30+9ZdsGhYKWtJU23eq7SVOAwV
Z2VjF/wgbo5uwvCuO9orMVvP2m1CWtbky+9sIVuN9NmxAOgcXu3jgwiAmkOuoBqS
ierf+7HpEvfV0p/1W/1ILkL6Ob3G3rKvyvEqBtc/COK4V4FnNfzhUTxyTHv2S+US
k7Uqrj1eTnk133JSCAI+MOgZLJNxz8ohb6q0Gc4QiJCmmXtaLywTR9S0wd532+ws
51lCSHEDCSz9c5Q9aiGr2GRFbK5VlDClLcvTRx2fS7gOfUmi3x7PJAofWdsfrX7W
lUjkYangErXRa/AyrXoWj72jskWkcT916NWpLavRsFW9pdmZGeAwRvag+LR69hCJ
JTIXClQd01CQPNUYjWRx+HnwKbwKqqDqsq92cjnF0V28pbiOXAHKJnFcA9apM0FS
qEsrtoDEYJADxHxyFLpcSmo6w+jDmoIvmHO6KN1Mii4hNkpwyGNLUaDn+6zbFz5t
Es4P7UtLxhSKzmsUFTRMILpMZlBvE/bTGGAch7k2AyiMk8rpS3BUYcRE24SlybhH
fcL+ay8KOm+9f4njKWp90dvNJ3Z3ThwEpdPIdGmZwcTJn7KAGBLmsqFrWP02m/wE
JjQN5oMjmG0f5rnchjjGqcXXmrjdVJD/R+fWLTB+8uAMk5+YBeYM6OOztP/3dXsO
Ir9py+EPWbkGPztpHk+BW+q1h0/d13t3pwfNrAo7+fddtGX/5s1U59EiOdprsyDc
xsxAiXqAWnKDmmA7RIXf6ZTiLixH6sQ80g9TTD4oA107cGwnyXjwpT0Qn3aWH3mz
zOl0IgVBsQuQfyRrkgTcEBsxxwKq76crKnwJSjQCLxS1NSFgXDu4PENAFSGGV0dk
/H8kgP9Tlp/+L8zeRfDI9ipGQiR+3lAlm3wi9Mw+IacBmTuOr2ajWeFwB9MtX0SK
DT9+rM9JkTO21+UdwSOGAaqua+7nxxHYJV03262koQgz3Vv51PYmjCQZBG58386Z
`protect END_PROTECTED

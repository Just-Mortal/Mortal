`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jbTuB24b+5dDDbmKVlHBhNbySzkbUOetk0rXNRa3Pt+8oFfjINIi7RX9GJD+4uJ1
zhZlxVb09c4/EsbXcBN3bTXcEsp4cvylXEkk5WnlEFYX1dZoOCFdqbunINuKOHrC
z5AiK0K8G9jN9UV19OSXtz0XAoVUbIRD1MMJZCR+Zu4XGUi7miTGtkNXrQ/XC3GZ
sqtiaX9uTInWhOkh4MwGXgQrLhMwgx2Bdwbjv/mw6q5TGiT5rOtefDjL1INBQKCK
xOggqzHZwKCZNr03/6gKjatpl6WfOCWq7SNH/vdNvhWSGNCXFQVsid+PdJVG4LqX
4nv/VzNgNbtdm44hiLdhGs4uzMds0yaN7AfwxkxbmGJKVFKf+E8q0uPpRSuklmhu
bmBQ93wDhUEON1kjW6Lx/aihwhU+hP4SSPr5/Exc+Dy/76BzBjdUnH79g0gMoFvv
QZTmmtlT4Iy6zmfJSqJS682FdhGSrfq3DuSIljATSDOzlJIWmWLQvlrUlDRhQRJO
X/g4yVs5RYl2R1iTUKt/CmDy7Iphqlpm17xN33EmjWnOyMeJ6+/7PLP0HO55BNlM
yo1IzCnePlbS8bKym8St2sZiX9mKIXOS1JDZBU2zYfKOUjUuxb34H7TWEA1poza3
WkBdaoaTvez5LYXw6jnBneSeetMw8gdqIxlS4sfAXCJ+PmOCSwrI47TtZFqJmTen
MKFRIaBtoL/GRanGxjYgKGbmHMJhW7AV3zGr0cge4xL3ujjOUUGe9PkGju96xj7u
fMkw+TyGfbPq9gpYqB6kMtzDlfaCu9JuKqE68jnDLJpLR0hRs53T37uqnGki+isP
AFbg6JzciLQenW59YLJZnQ==
`protect END_PROTECTED

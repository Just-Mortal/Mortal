`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+f2xxOoPCIMRJnkPrPG9xaM2vyfaqOOfpwZdJ9Y3XVwRZQRC73qWhqgG4/rb8aZG
vduRtiemmHYeT+GWRUxit+tKxHu4wH/XNHZ/fnYQ2SdncDwRQYqtQm6jUtX3ishg
KdHuVQgRWbCbEgd59xNYnOsJURNAHZ3xFdFWPkZzHQ/LKCS7xpufTtb2TafRIAM9
MxlCA9etT8b7Jol0y5NoLFR3XdmMD6KUi3DHVlyjsJLhc4Ivlv5s2BaD1jzbm/yv
gIE/vEYuzhVsjnyvv5hiNsKT7v3/5MU7HdQM+MNMIoKNjuWpIemL5U6IaI4gekop
GEcAiEmtJrVHeZ+vP4EcDIEFNYWsttRTjO2dL9xnga3apdC9I0OvcTw+iTaBu3uy
GI7acW4Uw9WATrvaMfYWFSRmDHAqdbVSaoNeJ39oe+uTRhgYhrNO/4PzLI7Na3AK
D43IEGwAQwDXu1WkZXeKEuGpW/kFg1INqWO6xC49cnRAduY3rwHXtHC78ZQptwDF
AGQ9gqrYK/yimq22GwNP9XBBcLsD8CKmraQDsprUeDRjKhB+dz32+5U1Xy3GFq1G
wZ+d8h2V1RgL7nVSl1RIyM4Us/jcLQv9Y9oSD6XTK7q+fTUabAxAcuPab8z/Vc9A
mFrCAYE8dN0S+IcnRbcp40vF79l5/+Jkhm3VpmLcRhil1hWK8sO6O5DRnSeFhzY5
R4hKPdy5n1RbePU3Yh4xQHaXzZwEFGK9I8Lz1fESQgegjIMIDavPqOwfzy/QABDT
wKxLtvDJKZ6ZeLeNUz/DoLmYUQBDu7o6ncHxAag1c4j8yGGW5/FzznS0IbdjRnND
xJ1gu0CmI5huYwSgd3ydbX7Jgd0Zdz54rCUaqmm42JILfWtIKQN+qN93jKjw7WfY
cF86TSRotuEelAb3TTTqNL7+BWVYiWhi7ufzjovbnYlUejhpLETKyyyaXni2LZSV
MFFPzyGfh2omkCD1Uz3wR4yOV5uuxitX6gzvBo42JEqQOI1TpQ74qYsVcDKifYYz
SMK5x2HRsCVfXKy4B4PY2RkhB46M2bzpK9721ROiVl5GHTFQ8VHyZMaY4DlYU1Ju
/J3PeCacF41EHfM5NUn12+LjpXNeZqRe47JkYW17RLfUxl/UCzZpYH5YG+3VnAmC
vs+qhJBodL5o8KT0gQVSeplPtTvaoidAg1DPGZl+7XzpWwCOv3JIXNsQcMgY0fbs
Qa721hrxQMX2nrcZwT2fRmeoExMhUpYXGF6w4KwJhx97RNZKdBEJOeoVylQR4fHr
snxyHnBqXpDWAnZqrn0BSeEBzNIyD7YnqvD5aJ2x8ZD/PZHB7DSLMt/Vo3lw7PET
xanqAJY60NSWXRz4l+JZLfDYLxFpbOtYMg3o8S6sKPbdCgSGNQee1JyRx99fVBQY
SWtZtPyTLPrIoywCpiZ9XE6cpL+xO0nGafnlKB10LFmHLct4tnngsN3ViJE0VPlm
2fzk4YvYCu+aXFnyQzsVFDTK78wvzup02OIQRWou1hx1rqmNNCNsThH65YsrAI9h
tSDNCr8PuORhwTIB8eQB9hLSeuhGRy4K40qcCISG7Ru1ecUUTravwB8WroV/Jb4G
iPI8MLl19fPetf23mmb50qbnvOlYA2KtMgb4ODfqo2iAnqt1hhfFnyXqX96iGRfM
NEiSYuSeicq8jfOmPUprP1FraFjQStu55IIqdIGBWp3OEeuM4KdsPAYvgFahXKoN
EjqpUztxryWRrisgH0tMDfTlErH6HFjoF6wGxofeFQjvXNyEAGuUAGRhjrBVO1ea
DtnSE5+oZsu566+ANm7/xaSIkcvkQK9oTZOA5l0ZjApRpk5+0YMuBH9vm8jqlUW2
b3INsvg5bCpLR9my8ipchjmOujqnfq5uvSjx1pMCv/b8Ph/mUrkN45evQGulFjVu
v6b9xIvJMUzRSBuyAgC2Uw0ybj8T1lPzoSJtjCTEwb4sxCk011otH3JAU2zj8SX4
ivT8KwmdhL3I4rfYCZKizLWTRcKP8uPSUgGRn/z9+bVT7tsamhkykpRI0b2faI6W
YJuXb8yoQZwjYo77GfEujpAPFN0OWtxIRM9jKKYyKg0hfeIDt889qdaAOBGR/n0a
cmz5K/An34ZTsvm/18VPfA9ADm7tcWo6YtKhWOKDstdG47JwAbc/A78pRlNhY6sk
bOVD8xPPJSrrSkfzlXRj/isrIBi8C3GNt5T7MXu1dx1r9risjYQnr7yNRCU5/MaQ
KLAIk/HBFdjvmxPY0Dl4LgRMRQM0rfirFeLHLDNGnCDE1QxAzUUJoUi/MJbHwiLg
o7blL6w46npKTPVXmaHqJWkVaMdZf8dlZddE3egbTzm81iAdZiNZ/rSwjF2haJ+V
uyumwYm1hQlEddOexjov85HZQm+EL5a1iP8VlKb52Uf0aUuxSIsaN2PLmUm+bWXE
9xpz1jXg7VAUv3Ki+cNBGtV250AR8k+ixr9enDLq7RbcEeWpM66pprb2IcsGSU7M
2h+PEpnTcTiZEvMh6Fkk9Z0Cgq3W2boH6wuVgTaqDjHtugojh/cwg2OBdMVNgP3Z
+LKEJGe7lsOo9mmV8TusgcENi8p1odES22xof5x/LdcLqLUeX/UqLuGwE5Hz2b97
Q11girEPwlNA/dN5leEhex3ksVDF0KyoiC1Oah56MvpaC9jY3BcW/WTyKk8D7yoZ
AVpnZjYlvOlgALnlPH6oXlTXJzj8NMLE/myPq3yvMJa5/bzxMNRcZDpsVNU44qa+
CSMYgfUgBVWwyBX/ar9VV4DcWxqpkfqX7VdYdW7rxkngp7lIB0PtVxlGWLZTN2Ld
bDfSOtYTZCTw8moZ349FkdDhkEf6ffVtTFAAP9Cmt+w1xfUXhknK5HwqdbgzdjUJ
iCCBLoAHLZ3rVSyFKzSy270n2y9QVoT6+c2/tM9VQ1BCSnHotk2XR6RJlVUcXk0W
a+h5+n/kbXGw4S8zBNzDUab00TVTq1SRU5rv4I6T0Kc2R7u2WXcJXegWOCoD1N+E
g8+TcAMqithMmRnaFGUKVSAcs5ZaKG44EGpmLkqGIkvFH0BbbHY6CnjPsZokIVx4
PkkJNk5f/cCs42e533vZyw==
`protect END_PROTECTED

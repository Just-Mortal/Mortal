`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mQcGqTr1p3Hde/9vA0O24MCGPnzIgNQ69nlOWkagtwWp95/uo1gK+4z0KchM4q1r
L+OW3ErU+wYgz5SNxw+5WjsG8z6/LGeGXXNAAFruUXNu8QNfxUDHHrgpFFmfMEFQ
6b+cRI4lOKTnl0bYWuUL/QXjf32arIKRmz37hZZcwoR61SxNnYG8O8zyxyfNBt08
IrLAPGV+Eqs/ntF/P3Fy2lUZZCXpaQw9Ao+H+78dtJOO9WKkZFdY19m0M1wV7zsE
hnO9fusVervzV/FEJySS6lRKIW9Fw3M5Tty9jmSua6xezBjpqj1L39VzLI/xDrhR
kFG2y4Z60fkmAtCp9dL3AipH/Xs+oe50zUCR6wA+GmcFk8Gsdob+7ZxA/mbNcCDf
d8/3Uk44L+/I98+MOgkdFSfMRigD4Jxhv6OnsyAuDjboKLd3RJ+4MW5PCcGRbeGK
hln15XrcAjblq+WgM5vNr0QdJ9Nznuuv/n4cMf0KLLiOeWBcH5GUnxoj4+GHdi8c
bRvxN9nHZyHXcseqeHCZcVj+lEBjADrMeTxV7YKzS07E0GvAPSS2Rsv7XRHWMNhI
GvCPYPpCUaTSuRi9JmHEbwC8HyJ4qxVYxjjy0SWK5pz64ai+vjDmcJXGmTT5T9gt
KZmtaS/Eavpf+jxAaU2kksBMCDfG9dMg0JrhssiuYFS/PEHaXulTVlD0JLm61+pO
lBQbSULcToZMVLopKVeC++3AzpykuN7/Lh1JSU1xVVRs2NYaZz8Zv7vSod/8pBXD
K2ljWos2XvB3gWkh3CxTwXTAv+2HtRjfu8TLstFGX+h6MxiC9I0Thot6+WOEsjj2
6OTPx5Sveys86KWk0b99h/D3VMMSJiyTOrm7ZaQUMV+DWtF+JeEcU6XXsGeXt1gY
JGJ8jSDvISjoTRIAwNIxojef31Gt8wy+DR3XVc5BdmOvn70SybG6pfWcvY8NpHaO
jPJ9yP/++KE4bBXVN199RgQNM6itT8tkrxnjFoSO1FxdxlpLexUPhXdfci8ZO/+y
94SIIakWZSkeLK3E2yqdrjIWCcVhnsu3op2QqEMxFmlkl93KGqvVua9KsvY85rg6
3vgZch6KtrmKx3+5ceGIpWSattSu6aXa9xO4fgOwUFvPLRmJ00+/1qihlW3zy1cM
mQr8FDQUzSTHDvH9JlTc1cQwYVlc7IPnpFjSZEz4w66KCkaXopMX0jjD9ucM8wNM
AZVd7FhS24rTASop78vCnjZ0khVOVAQtvYWaK5hiZgZPBPT2Q2WeMGZVeNSyZPXn
GBwtU5YmiHIGO08IcVzmBdVnDtTsUOp7Qe1kEwGXtWc18w4UFXicP7gpTAmpmG50
/4+v9nTuKMAWLnkJ3NZNI5quX74rBUbizF0zMj9YoGT1cqXzwf17q1h7XWGtG9C2
5hyL6qNfgx3iktsrJi1rTQErfeuLV3/XBqe1U+g1zv3wxLoY0AqcLJwhEIfCfTv5
4TQvFYECl98Ij/hRXo1hh3/bpVUnnW4WdYPNGBSIuEyHQYl/JuNqmsUmvAAOT3ca
1oM9hFVXRfNu4RNPbFmdCarX67Dxso8Si1rvHxS0Bc7Yp3vtuqIXy9bwPbxHimTF
OYWW89nTcJ5N696hr0BUfy6JKILZbaEdzr8FyBdD7gLWvAtxcCYhGCAkIadYFYsH
iXUBUMuGIqSn74XOUZcQzjBw3v7NTLRqHvWroRij4fgfmPdR+VlgfGHwiUWpkUi5
BkwEpb4NnkhhblBZb9q7MKTx3/AtAKQMyKDIfbRgAwZoUPv2hL/ZAFfCDTJThy+H
gjYJBiLwYpULdijbF5Uo4b7+ofAxf1sqXW2FAvtoSnjb23t1ZK+k9CmG76lthexy
kxz0muhaag32Y9x/wdOe+iDnkYx8bGPV1VUyXTrXAblualz6U9x1WmTRoBFGiKo4
+Qz4xUevdgiEPrzLqnVx6Bc+mit6eTIHt5yfcd4VGGox1vNJTlso+TrcLbROiQO9
379utxFWY8nRr3Y+++XD06BSIOEXgq70wLNxeUiSqFLna11bt9p2/gJ/hh1Jxvgb
BT6WeNxSSoaEyY6jTV98JaXEmLqtu62EIgt5fSN2CH49HT/gk6UeoNdQH4x5Gyj9
IYbEBJHxlYbkPNnufDltDDTsZzBcOPhP4hrFnZgblVIEvIeiRwRySjki9uHSuUYp
0wmF1kvY2ZvgdOwtwdNejIXQcpn4P8p2VYxL+bQDFc5Ax/GSGiNS218zKF/bmcSo
1qOymOhoKfkwAEAliPkFo5zpT3OkBQ7+2jRiE9VcC7nLSkT+e2B+LBqy5CCh+cyW
qRRQkZ2Hx3sE2G5lG+8cJ+/G+e9dx3iVtlNjogWpMj2FE22sFUt1vO9IbQB36lk+
zdFk7x32RHqciBEJdXC/O45XNYfRmBr496YOfFXiQfvOW0tG4bIBCsf3x59iopib
Bl9rodHBx67eUfcDduaAMJGc/ikpJFP2oaVJTx/AhzkrKoOvFLuwJ/w/DZdVuksX
O8lL/+Fe3csFQz/8Bclj4MfiWgTG067ranOSvmCKVxxqdm8IGjVwcXQA+ojZZrJ2
rXwWTsx8ioDkSPVGJD9X+frKjAqkLW5vEJs1niA5gqn8YfcfVnM7GtifMxoPSImT
9RvBcC4NPre8iyOJSqNwYpVYlmlkqTVSc00rmcNbRmWRYZNAeYuKFjjXxmPfkFpv
y33GSE/9kSFdWVkXK3OMV26FXaaKaI7fO/5sb4pEHHUBPt5AB1DsQY59ph/9Gdgo
CHQ2+v0T3YRvg8LtssJjScRGd51IZBLcgRsMTQcQtVtjWc8IATwY838Rq/ngPUV+
wOqAHPZtwm7EcpRRTe8ETfs33MSeNY0jHfJQN8k/sf6XX8+QfQwQYIPF7K9FWX4F
9679ptXa5nKZOd08j28mUUntGqn9ElepZPHLM5q49yE4rYCygrKTO1yjpC+bbwGv
S58TMyxVvYG0av7GHMLeiniV06vYz0F3AOhDDGcLWe5EZHqYz7vS9CcLxw4mFyeB
ZmiYuLBvhBxRjHM802MoQJWe0O8mg9W6RaPyxerjYeou5haQhHQxLRvRnNxbhkGj
lWBGatNvx6WDM91P2ZtEY2Z4DZwLMJah+Y3zoaONARO9po1viajy8G7EBBR6bKo4
DvCiacZ5HmSBnNpfEvDsyA92p1es1CUIGllS2mJRPBwxHFAembAWX/vcI8aGftTA
zR9ivdgQBxyAoLaf8uuojj6qwK+2H5Qn+GgLkZBVF4e9zdLLCWK206I9m0Ke1KCH
HAzW5+aedvGcSUmMuXeiZOiSNUnlUzTQUJwgkhLq9AmPZ7FQ12ByDhd9aZHXtEUG
XS2gJeW+P8eUfTgPBwhzq3VZkYEgNKZHpSs9PGBA0xzzC6owTIqyoN/mYX48rRIz
V1uXr4I5k+ij1Q6OgHTVcZTHkzpdted/e32cLmXksFLUzeXcYx+nSOoBbukSoRnj
YzsbxdeVKng7eiBK8IGmvxFWZbR3t8hGyqeysVmQ00TFcR8cVU1vVFVrH9XlhQrU
ytR+Sau0pvJVwGLnn5sme+FCNBq81qdfqSIwN/9qAmr72bOdMteRDWGF+uFKYZfQ
+Y6Iqe9bUNKT/56k90uT8nYwP9PVHMai41sETlOIxGFALv4RuR+WD4EQUgdPGHAB
/vRRAu9hCjTXzA0Zd3IOt6f6fx6tkjqVv0zBZMXYanUrBuMEyyNWomawjWP5eKfM
mqaAdz7N90ZJDD1/v1SZe+oYFQDNWfHBfNOK2daOcz3oVjDh0FSGMfcQNLRMk7Qr
VTMY3M9a0PAfbAkXx56eP7eDgUft8JcYhYoOKMj4ohiXGpR+q8mHC3/3P0M3dhyK
NZmr/707DksqaSlYj2fmOJ8F8IEV8t/xGCki6eIBufE+opJ2euklNbVqnjnLjSmz
cVuY9mTxDAko+qB8trNXDii1brTCH2jSclWU2UyiB7Pm0Bg6kjUv/sP+oA0gy/6s
wGeLP01obbaF3e4FSxzGIXGxZtAxM5xuvCbomMjtXw3dnKJLJB6Bu3alcrOwOMhG
K9PRYOXbICB3kReXIzPLsNjyOQhXVxuQEYilXVWP2jjR3wuzEqC+5LjuctEOSqi3
k+j4e3O6vh7YJa8UJbJTdFwnLfr8bAjeTZJlITBHQQjx0aZl5OcXYg6SumitAuiC
mvVsQnI1WBtuJqHB2iZeHX3prPCpbPKJ7e6lnBgj4bzmMDojqHaIJrr9wtk5Pmdk
B+Mqy1BgLRPTRNoFbL+XjRzCMJLIjzQyzFuyIN88ojZht8pMdM7yQVvZGYvjSbsQ
6Ma34j+RHyyUn/wmiJbXxCAKIyyOorkcoMwkHj0wd3WpdQe++o05nmq/7yxnIONx
1TSvF0n1waj7vdlBiEV2v2s3v7L1KGGBCptpZdQY/j1ZDYL7sDwJJFEtmGdEp12o
JqDAngPs6StYEdHf2PSDbW/KlVGVMZNN2D9mgDek1b93pwDpZcaRfxXAjcdfL1PA
/ZTuSuL4HsjmkZkd9Mx9+VlyukulpEqJDg1iJ+EnvBiUA+m7MOZvALOiv5io4CJU
ETORX02uos3cOL53vBaSKg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qBI0QvQPYrj/LNz06nTqOXNkzhdElh6MTvUo8EIJv4OXwFBCtlqULb59IxVibhc0
d730mKjW/fhYlaUwqzlrFEWQFMVNbDjUXehqGtvHaxW2hrL0Gj+mP6cGrQcB7aKg
A9pysf0b54ewjA5vbt/h/iSM9b3qnJxniXltjt8+0QVhIG/5zr3k8qIx4q54/vKu
0dwxkJ9nCzOD7WvFI5rFRvbpMsKjSyBizRLNlaUJUlXaubCfFmuwSsWEziFXoOeY
6SdwOXUxB0H0yrhVb8kwKaOvD5BrdDyF6mDGnLAeUOhBnB5aPQue8CfO4cBoub/5
z0NG4pz/N9vZvuumtgI4yULAiMGybv0P+V7tPAEYoDGt6xnZWSlp+Ch2j7M/7SzA
GQCpHopoe8uPN/GHxsDrF/ofM1/2N2Sy7ew8inUjJ/PLhuDip9BSWFgBbYteYMu0
JlqMSSw242zC5VYhEkkLgSgmoabZIQQN+xfqQZGER1azlIRtdDJpZ2Wy4oxZx8of
GXheW5LGXUGI5qr9araI9/va8MOee/IN6Ba1Gyu0SJUmcmIVG+FdWVbPHWhKanon
5lJnwF71digxWU1Jv2dPNfMW62w39L/N1hDRBKwwselW0UlM69zZ01OBLSA+KAww
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3SlnoNOuB4DuDnpV00ZWCkAIGOA/p5jgeqHwUiaSz1Fq+BGbFbUxfyq16kkaqVK
j9XLEB/lxi1AohBaudwQGVKwFjY0JKFl/Os7bwKprrNVCDcACYokXMYbgRLH6HP/
8JJp5iPbdcN5Lx+puYkfsCpGAmtQW+9pfsFkDdZcgL9kuHHj+84hwsxdDVY5yPCq
L1jowY+F/26kqpfx7QrBH68L5+M6mgBz6ptRlv9bTVZw6T3tnHQ1Wigi2MhaEyq6
vSwWwf8xQfUuwb9/HS/F2k82Cbn6egDwZNmfn/VKWBgry7Icfgb1mWmfFoBTv9tE
ihPai79RCw5QORlWfC5Op46NJf68Ihh8Yw/FrV9an/arkKH8XXT+QwICjMIgPoHi
O4rNiq5yiMyIuiLmbV9io51Z+WRMgNK3x4ktx6CYtOY4jeaHlLPUTjscQ+rKaAhC
Xj/0ySVn7p8MDkfSLmJ44ZuaqU1VCKSXzVbtGHQ+glS58Zxn9RbjZ3hTwfEgtMnC
LBxKTT7wUl8rRwxJ6/7lTqHmKDBdJLVyg9yub4L3HwkYA5ghtQy48N2hCVlM5k2M
2E2gwj3C0nm9wiVByKZHKLPf21vDrmO1niYwDlP93q/gNgNTFmnJjJTPvZsUqdqE
mhERDpJRtQP+NDgO5Gw+9ztU5mekbwF3lTmOk7mULLJuwMlLl2AxqmkmQI3YBGJg
PvqvjXyhTiXqhTIhOKpScksXCE9+gHGqKCzBSKYFV5iTAU1oxLeLQh0h4xstF6fH
RI5oRFkqxCeZ3jm4reRt7991+076FSpXruHRMxvTCdLbMiYHcIUYfeI/QCe8nyw2
eiVJz58SIHnkbt+IU+V+5xcv8K/S/Zk8mn47Y/Gz7ivzAixu+nye6ji7DGU4Mjb4
IeyVoS+x/Y6N0G632kLIjoFawK4esqISOMBBq+Q9khqc9XSk0LjYa9xuIuAADyw2
c3xowo9cI6+yD/i5jnAAbQLQHfuRNPWGf2iC1hohH/3pf3sAMY57IPo6BZ7i8AsH
0ek1fR2mRwVtlQQVX9NKxiqnz6dRHRQeFwu9J92h9TDajuW/6OxiGUFDG3PofTnM
3rdiBHzfFNNHv+4fZFFrfuffJWNRdcwxEBhECcOtjhutwLB8AqXRo+EmvE30aU5C
DAyhjdF8NbuX5LDwjFeeBA==
`protect END_PROTECTED

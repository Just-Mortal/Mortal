`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69oyjNi4RyJ3ZNA3hoPVvR41X3dfwxpPFMk3n2G/sGn/TbJlBf/Vp1EoXgnYQVjP
+qxG0+d/eYcUAy8iti+e52Rs6wnfIIKsL9Ixe4oS9UnojU07e+GxDxE5Szb1Ytqu
IodH8eM4SKU2M7yX8FhQ5h5/YKC0KtwPv1U6BogVuDeEcsOYr8iBqThdx+QPK+PL
yNGpgUwpMb203jXNZVtYvT+d0B+8N/Dkvrs8mLk2ijLfs7L8az8WGDEFE4tYucYq
Arqrxr9gONjWwZz11rg+MzGY3mUcOuSsH/D9h/vZ/ECZ0Lyz8xJM43BeRcGcUnf5
o3efwawqlA6C3L9xcaJ9Ibqa4a+wq2gmBE+r4Byyrv4ECin0fu8fjCzmm3FLQR8/
TRUEEd3djhs/bn+lDBT5rwhb2wDdmlPGbSHo+9UcHCvhBCBhR7oD1yCrMZcButsy
XaZ24EH80EaLZZxbV2rQYY4z01mNsI4kbhO3x8MBGG88C7hE+Nfpumg1XM6to0Rn
30PSaVO7uwEAVnacfeZywtsh0ME/tuY33QRy1Wozovo8n5RrhUxE1rY4DrzydgEx
ZOwQ3JJa/iVcecUnjR8gSyJbmBAvA4KKW3m4vcpt13N2C+UTNHvuJ+3HTi2PkUHq
pDFua6WtCZpYgpcjOEyYS3hLlU1tjr6EVo+9vPgkURJh+wueIe4mFebTfV37fovM
QhTA9WTv6vauyLsx9HVGTB7OZxoeP09H1lv2dFWLEbI4YwxTRpCNS7YcXFGzaZB7
SLDJiXKiGUogqJTDD2nhN4ZLsJKgkR/SnMQKg4D0aytF2Xtu82+z6swp7ze9GW4q
30U2zSj99IOI0So1WJwTMD1b4yHA+qRD7uxprqJnz7If8blXAfuVG6rBHqe+v5Qe
1EsJcEauqw3C2HdJyHxDIDvUb788cWcoabDnDohVOGMRYMlc9EAOm/C//ADSoNYR
uQ8RpOstw7sW5aaCq/sUkBABO0aK+1FnzIPJ2/Mjq50gFGbyUDxEZ45aRJ7Enex5
2W1R72kyAMlC4S8QqLc1gIvso2sLMiK4LuypdDPiGJJVjFXnl1FqUDmzUrJx1WLi
SttQYzJZTFtk3odZoWmTgV2lAgRPQr739duTyq8qB2v9PFo9HO5QcCz3m3OiLB6M
DaX5ot/07e73r3HPizVfL9HZ87/p8ymt9jAjoZ3zVPwHaLz9NGtjwlsompsI8NjA
JKIAjvTUky0mD3nXapmuTmI/JKHvgKM2g53NOy3GtmmAUlbthpQlFPOK70jKuNjf
TSHsXCiI7oCAnfF3WlOcqIYLY8RYKZXt5G/Q71yoFAOdV6nD3HFu+YC1VSR7mfB/
woWbOP/8Y2KdAyFe198s3FjjbkNpOQtV3IX8KPyvNg2n2X1EtaDD9HLthopafuKD
oelhl3P+vWlUk5q6b1731sWAldk4vPhzytVYMVGg83/2YE5KNLWHzOv0rNqhNcCe
gcn7YscKwJsAM988nQ5T83QdW2C2JnNefQIyK8g6NZ2XnKEz1chFt7R3wpo6iDUY
pmM4+Wejt2ffHsfzutBrB/0PBpEAgrY9EskUkU8v8sHA6+RPyQi4q/msOZOy3OwG
IYDEbHXnpuV7PutyPT+6i/KJFgcwLBAmGAHbVwonypX34b27FP50w3JeYT9xuzZQ
wAIzEmMmpLS0AyG5txUicpMTHhyxVdLB9XR8LdgsJk2Ah6v39E3l+5YelFfUt+D/
OCgWnCFl29zQJkiZubaWAsTe8DsopkcMSrlUXodOuQ7HnAOWOnGhWbiTBMYomLre
R0vzAuoVmo9yKMJ51KMvY3+48x2WWZ3rv6ytJ/FDrxbtdi3QRLEfE5ESZ2VGxDvt
22CsW2n/rqtVzY84XB0S3M2tJg+omQOVjcH8p7qOp3DTmYUIlIJS+AHZZOm11WgJ
pjIx8rGw2LdUV+eNyw7RP28701CybomaLF35XK6JLWV2Lg5mXoyGgvV6ytCTkbI8
GFTfAPiqXOrkY/6crYVGpVXMnmPzhpVwVR4cRrCJ0ZXlK6IGzE112GfN3nFrMOeq
NuazUTLNowM9A9DlL84mJX/6uCIukf1Q0y2rO8RF/gMGWW3vtqm3jPCAQ9QbZFxH
Y7eM+Y12vn2qITDxXc4JabMat1HAvkUYB/uQKgCVPMVIwAol20Agv8OlGp7S9pSw
lnCFQ7T9FEPjCyzXTO0OxZ6qkQ5GzLRd3VzBXbBkXNgMs0TPKfBLYod59uwvY6cu
HqgRBT4ynQqVL9Mewtdk1hXN2dzR/GNbcc5yQAFR3iFVWDAlmTIPmi6IsDU++vTH
UlTXr6hL7nfvPpUYHXcXcBKfnz9nW4PXRm5Ao51jeAA73bbXa6PVklPgjNlFsC25
aKs3j11wwneLCFSNVQMEP2VQ/yzr8S5EVlDuV0sOC1q5w6UhbH74iOcxAC1ghozG
6rrEn2nIcTCmZRnl0rDWxT/1Liz3ZJI0bMOEuTBpYPv1CG7YYMSCergz/jc7Zxye
ZnXc4DxxU8MiVmaYWUEzmdn6ZY6E2RCtshbtzkpZb+tRyrTcujrEZoRlW8V9LnsC
cDlngI7WdTunkcN5Bl4P5o95dgLPkzVbK70weM2WbWhqa7wT9cY9P4jZ/fXYd7df
xe+CoCp0BLAyugOfy7CV52a8Lx84O+GJmE1E2sWEk5ICqhJ21WIMI9c17snaNXjk
pmu0MBIeHSvCR9vKXIFx/20NiVNAHYai+HQIs4Hk/AsR24EEksrYWUId0fNbqurU
D52aA6eg67BvyG46PFGbA8GhYvxnNswarwymeG+Hw7uYNW4jrmppBifRvVydj6PR
TqwZ/uw+JEO2gxaif/clO/DJHbDDhlUZeWUa0zx9QxtuMSgdbpQnSQ8GHftAeqR4
KBZkuD6Lngxi1Po+loWiqKEp7ZUum70upDEThAZAqhAiX4RVTl9DowUZuxKlx+vm
d3QLZD+f0mQKvCwScSGOsnekaZ36iZla2bILvwD81LEm55P6qbAK/BTckIvn2IHo
ZOyyJmmOrC/LES0giB/B8kKDfoNE8RfTKF9n8NzjCW8yV3SlHlHJj5D/A2TMg9Ar
y6ERmGGF+c00Q7oZjHVptg==
`protect END_PROTECTED

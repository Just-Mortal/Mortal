`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q++Jbk8i8YBslPakwJB8wSqDOPsnRzRNntSR2+9heglV/05XE4ZXONifUfS08Q13
cbEcZm84HdRIjoECCggQG+x6iPn1SOwnYUspXFZEAIdBy59GTqpgcTxeh/JU0++z
LNocf2KgVLQUS9LSMYTMZTiI1oRqlqQVwdshkv15VN7Fn/EKgy6YAeH66RAkSKiV
XoVR0LFl3F/kScj0C0IcV+uNVnwCiaF6jrNtEOJhhViw+Gfg57Th8u70UZy7dom4
nxFQvXNHi4Srp+CPcpN2ZqN6BkX+VaKSNUEkmsMlk4lvJOe/brT6y0WwCCJlHQ1D
u2S/a9UWn1MuQ1T3PTlo2g==
`protect END_PROTECTED

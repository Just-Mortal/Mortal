`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/XMwcz6p/gwStxkYXOLvxYP0axHCSEqlyZ9hXh9zHoRXv39Es4lzVfrDA4uT/Mix
142XQFrjM5DKyHRYNujvcWSV4bAFBssPcQXheeJcWd9tWwwKjRSk74Vu1zGZVMCM
F9qcFjCtQIaNEFw3gtrs67WzlWsXDZyy3iwLxZghJGoiQCVLJrpjM1wn6LP5krjI
6p+wPr/2HrMsY7G8uEHTSGUD9s7SAIzBja3xv/msM/4S4OeiRVwq55M3ZAiYkimS
WvSRuaxOBG4hkeg4sq8+sngf619wVLvlFLMnbTzU5V/4y1bbHbZ5g3c7NFcmy6Mz
82A5nP458mI4XbI0LpnfoK3MrzG/tJEpGxWPGqy58r2x1OoZ6XL+atsLiigR2E3s
Mpfi77+8hlioAoBgL5wUDkBbAOJgzNy2zuJITSypU0fzGg7yMv5gOVuaaGZWjTDG
7faEQ9ZGGaUh1XuJPYRDq/JbffzcHrNfucdw+C2LYXy/cXGk32hySQoYytOSpdXQ
qAas63BBCj95vTPlKAq1u6ecOzl3iy5hsihFwfhbksQcgp91KdRmuIqkXJEjcJsB
qtEoCbdiE2C+EGypdf/QDeLY1oGsQkZw1VxBG5dHcTCFhkCBOvuF1LCMseKWOGYt
6S+A7PKnztPbAamAX2q9ELIArlfu3/187Hye5GtxFjQAkFvVDe6L/bAbxWgrDqKl
vCzZrEGUveyB3n/2D/LwNejVtvjpjPiHN6mOqlY26xu8biqZn4NN0Ok5gIA4VPkx
kAz8/Q8HOT9gOFWouAHsU7SQ1c+TEae1/MsLLRFePRDiuv/J7mW4+zmQmkt1nSb0
Mpqdrk/yaHDu1DdBWDIToNNKZCHldyoFc0oLwweHKDJe+ueH32Cgo7l1FcVN89kj
Lccc/AROEdIU9Q8fybhL29Vt+vqIAkMGAVIE9BB3ueV0ANs+9Rw5BJhmqK+U7J4j
1wJ7EfEEAtTAqbPPZ5CE73gwAS2SBBOY1+2iGGyGgzJ77dRB2jxgMtifOcL3yIPg
NhiyLVV9CbOUX/vdTZPL8Em1qd7REtLipfq9Z3SBHGaTaD3OCtui4qml8j06Hsbv
HIDK+0Z5z/AVKiwwLz+fg5fA6arSQW23vMNY3XMkU80N8RLEbqN0+EPSbm6ueCWc
zKpHjAPj722MBlmxcqbnY2gBuiF0v9b/6QgY3QB0OiB6907PmK4TTebzs5Y56SI0
aR3csLDFVhWUAPhMR0TLNQ+IPkhX59OZyCckxCesgpwBskqwqtnG7RPT3bG9dhoV
oZxSfXDsZb6OHpq8grpOcePeaGvNZ3WV7SPP2SehI+E/fR5XUShWC1jMuukUiwGP
5j1S3dRZRsLMCnvsXwSldMr0aYF7YpsjkFMKJ0ahOsN7ZBDpP9gudRP+2z7E8PNL
GmspiMzf/cgX6nuTBpDhG02VkZWiyXY3KmcneMLVnqlIjb4kGaO+URgsUZOtYKC7
DRr3Iqc5UgK1FRv/eO3hJq6IGvnxBL1INzx9+jZQ4zxN6gLRy9kbOBjWV0wkxAm+
d4M0BPZwuU2RN519ibMWH/4hoB5fS6VqH6E10HSMfCbrYgXHnsbXG0cEXLDqf16R
nldsnZsMwzzef90tZsOqDmwbargDx4HrPQ1lX6TUJ0FVVby2LAY18hBp1JK90ZVZ
gkiV9hjnjcPSp8RM49HNGrp2vsMFMQEnfErirByCvJ5N1jw1Avd4HQ3QaGhAjbZI
n/rmG0JTy9JcAhQ3zTDdSBwVXG7Nr/jnoytgGwMH2yvX3pKhC+ryFk5zb6QvAKlB
XGeCskau8YLs9xk1S0+QwGOB+UGSvFRB4DsAi8f+XExYCV8U7zFMWvBaST8gJIAX
kt5ZvOb2+COvAWSA9lyNRBk2MNNXrbrV7Wc/5QWgapQYWIHLGVyyW/zZlhogwGFZ
m4kSQtGkC3MQAlSwhcX+n3HnNbScW5xlzLpd3q1q6fRsaADXySMo4He8oCPLerH+
n2trnz+S9QOJC0wXaPURnz9MhvWslGVh/8pROn49BcuhUHOd0YyA2Nx7PgteD1Tw
qoqihzGILNHU+BaaGWqaIAA3w53wSQjTNBheR20WZ50XJZAGizZKToCPHhNHERsU
XW2jjalDR1Pg5kECbqT7y4yjSN7peymDQpW7fcuon33N+aFx6JsRvZ6/bnZzqmYl
v4To7lIth/wOYxA+jlaU5sqUL1tdM/8QlOJ6u2VSQdItsjJYKv3JYhhcVdTuWxZm
FpPEV1b1Dtib/hkciYJG/ry1nffX2t92ydhwEzOrRhOhfywoovMSLUz5nV6XRtA6
ZhFooAvjvnj9gviIUvV0nrBiM+di8rs9pZmyY4jjSc30kVuCA8kp9tcePVADH/si
+8E60PdCPoX3GpBHqrhJP6iNYH/5fuuqCQBm1YBDqgGcB79JF9D8tDyPk7FiIMwz
Jl8NbwDHjxGaQuI1mUkGWkqsmfPxczMD4HWuhVSWXd5cs8UoE4TUzpdz/5g+voYU
wN6dY+aCIIrVUAoGKM7VBLmM5kiIH19ZzQYBSwcsVSYh12OK7xhWuK1RCtgAwdDT
K6UG/LKg77758YyG4thiE/pBjFyvx6QXWdj4qR1tLzzb3fcXEb7Rjshy502W3oXv
rpB8VhKJREBsnMScDFleiMVmaqLb1cTN2P4bdIy159eE1UlqTJIfdlhlQffuDdG9
v+NysJdTSuEaKMpn8moWvpXBCPv9WOi/bYHcxykglZHVF1hyK9dEzWAhWv4HkDQk
2dpnkJZmSSZR/Su9/MF0wONb8igAnv34RJkJgT2uI2g/h4BviSEjrYYMTOjvJ2iH
3P7/Uz/OtDFG2rO08IsRvsV0OKJdRK5JmNw7rqj9xdUTUf1qL8uS3WBVj1Z/5ydN
dxqxOQP3NVy1a2c3iYLbP2oaWn/2bxqcK8LJSdTkAgkbtA8KcXQbYiOWkKbr/SZG
mA39sQ1dy6Lg8hXW7Uce4OnOq9BOAkhdRmq+OH5bcEn/EZqGF5RW4natwQ4sdjNJ
bSDN9RIXhFc81lr1xQyYklv56WosKN6K8PUVJ1P/fiLh4piaXLCxB6xjoDwwUCob
r2rBS3qykJYEHp0MJsDy1BsnePLhc07j1xGpWAVp1Vr2/oM7NonbUuDWQN2NiREj
2j/c6EjGy4XR8W8PTAYg8KSixpM0MWYxYxIMOWHvvUffeF5wMom2Ltni/EEPrNTt
f7t6ZOAei67FQrGNIHWNcN+c6JbE7LT+qzHbY3pxZWXsO0FegvODr4ICb+T1aWth
hcSPy/BChy2/JKWHvbzKzFHtgDiq0I4o7YGyL/F3r3+oxGm2DWmbp5Ou2K1SMu2R
RVEFWiqIOMb8aBsI4j6D+4j1ZKn5ArVc7g0m2HAKrRGx/jl16rk9XAMTwXWtWKaD
cMPkdgPcsTbthkrfOeAfh0Kb2hN+NPEy4AeWAyIv9mGrZxkwwYdNIb7Skk5gn7yK
WT59lN81y0zRWwSFlzWvGFsB/XMAFDpFbCR1RTxQiw7xQNjXRz/uvGv4dyC7e3rh
IsZ7fZ2cpmxisoasXVSSrW9JGVkCRvTekdXmGhKqFu9GMhkxxvgGQ2M9traAWOpB
qrRPUVYgdQCD92zRyeLblArTl/lwIPmMCuAcldIC63cr3BcQi5SA9vRDUCP2vKwx
yBcfepkzX+tCADFRe5UmsMjFL15qGMRDvnQhejAGrarYWfXovzXT+euN3FDrGBsk
X8CZmqed4xtEOtOkc1/oRTJEPG04y0csYo7JUS6PNIHrmpZvxPite2yv5Z8nPn6B
/2ip7S/d6vXCCsnJ0qxN1HwSGYmTSNDt4sB3QvagnhvRf4u4eUlV7Kjc6mHSRr4x
3/NKHTfjFDoA1HeuEyEfh1Yu1P0g+XxgomfPlmD+p58QtZEv6q61Ee5fz0bgJXNI
rpTtHq6KVyOE1mLDn2eVAPOWPHYFhv157Mgxjw9pZbBoOSXFoztEspT4vBmX2UAn
My2cmRbPdc7FlrBKgj6u2SpCLMN8iCdPgp3YtBcXLI1p+4PwXABKuS8u1jcm2mfh
JPYASPmo/xXpPAL2gbGdKZO3hY1j+Emae6rbbht3fYyS0pHG8VrH9SC2K1Nlt8ow
pgXvqFvdxkh/MkxFxF1CZIHzdT1szvbbFRCOnMLPhmyu1mC6UbyCqp64XPBWq6lf
bluP6w7F3TTqppNKmvTSckQ1nZMuxjJzmHjeix4Yitjm8I7nv94LFiCwYkMbvoUL
wEqPpIvFlFBid49WZcNlmA==
`protect END_PROTECTED

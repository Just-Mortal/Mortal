`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asQ+2CC6xnKLCT/UNtgvodo/MQ/DKPBjFOY4W2Brb95RECtsKAjSMK2hyReqy6gY
074fgpgKSip2LAel73tkDIwyRHm2Sw0ZsksdW3yQBwzQZcQGyJC/6nwjk2MxqmkK
M2f++0X8UMHPZltNEw5aArHMnUSwWkxlPNxtUs0zP00znrbyVcALZPXt8cFaKed+
LebRJPbLpsyMEFfklg9xKpxuY6vH9I5ArvydC9y9EPL7fuTsh55rNjwmUNdybdXa
FK5lVT97BAtCOrQ3n7yBv6lEMXhH1Dzvjozb2nXzQvNjF23rT/uZ70CusA2nfrJN
4SAozMAADnKQWS8C6TH7TPYfgV2xOzNsTJ+Jy9UH275g1Qp9CoxY0L8ih/qsG2tb
SiRoNaiP1/tPyopU7uQVxlwBJo1Y/dISnH7u1IdbFzowr7vlu+P00HRcimT8AXQ1
4eq9YdKkpTZANdAPkAlDr+OvW4Hed50KIiUse8n7mCN4moZAooP1cFPI/5TKRc09
bPWf8XvBWjrPrDW7zMf0ddE7xQQ/RMnppmm8GIvUYsbFqhCxoO1l0LZTaDn9Fbge
wvZ4jYniN3Vdyhc47+iGUlBJi9stgom6r+cfFR3SnxL5v4LnwGWeAb6jb8jxzX48
gY4HkowHlmj4tduD+AhXxxjFBqC6yNvopX3RJZgXZ/Ce6CfKuya3Usp/rx9S7LWx
ZUsxamNUK7gEsKXSIHEkBAuqOsaU0saGPYBxRk4q8peSa9ocWYdAqPZQijP1/9yz
pVBNl1u4FjdjneQ4dSwzffD4f52eswjQsvgsYQdMciUHQR4fysSr4wJAdR8J/pwO
1rMD+kSidCkCGzXSIrmmYi+uKF0F5d4Df5ltaFD7AQ5ojYQZ449KdwvfhoSRLr4D
/z24QB6MU62n9Fifbe54c/iSa4OlBoGej9GEZiqe6iGOXAzVlSGREp0AkXlHBGcW
jz2hPrnoRVVQ83yHTknLY/+ZNJNeYrjc3/IfC1pBbtmAH+j+bhe3JKI7ARNb4YxN
OMiYwEGuJoHz61FajdfyXQt3Qdmow02V4QJkG8wrr5nGBrn8OG10KtD1hFHDI5Ec
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TCgP4X0feFBZs9u+QYOqRBJdAXCegebx2Mmq4bSAkljnLxpVfmGh2j/lYAskZJTg
qk4DGEOZet/1ZvONrusWEHaQqIfKCOhc3+ly+T40OGlJTeInyCYzl9PAuVSN2Y9e
aTNS+bCaKemit3n5fSjuKXsQaFN2PwZiOF3PDjZpfC3wiMvyOgySSPMldG3GmK7P
BswxvL58dEMKmsq4pbBYS66431ebmhXh70tWxrm1RydwX9ThVlGvpT+cx/4rijfq
cj6KrC4UdOfAhLNvbhnkpG3/er7skQXpTldm/oH2V3SDBbMpnt6jb4cqtHj9GRLF
PbGK7j2TGzIMN3DuBDTGX8fTxTo78H/ChFvOPBcUcZjUGFCLOhqsHzH54dxt/70k
khKZamd1Ir7lu4bsm93ZT8mk82D9QGW7sXhs2uyI1IWZnZgBRMcvqWA+nNOwf/X+
pTZ4Ym+mLOxGD7NkB8au5DwEf+HwXdSClx1w0vBFsI617CPU8+PcG1DBIz8HREE5
HaT/tK2dPrHpqO0EWBVd9HANB6gUV6MbPIqfuAN/aRWNr10ZLQ6omL+5BCmKenxN
OmRiJJtVAEtwxXdcMRoJ98rCybERKnPFiw6N3F49WWkiVj96DMuGK2nS3mkAhqxT
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OizUz2OzdXFg62BcfQ30QgGBaXkxaDRktAfuc323mpJDWk0n0f2pGnKZx/lva9Lr
pyRgYZpug8QME8lPKntyh0y4TnfZIZeiataMb44UDAPrpqI8EEvWojvloi1Dwax7
f7uz1XNOJgfiw59+S6Ai5Qo5wUwbnpi0cp1y9VxgN6YxgeQIW+3qLqYYlmda5tfC
szGOIVrPQSlJm6bOdvVFTA1xeOhAezf0pJGpEea7s2XWH8XoZGf+/KoXzL4LfcYh
RM7+kx2sqb3Z31QkTC3R1Y6bYdlLy6x9qRY8sFpCHlNRSJrJaveRG0J6WwNaD93g
YydupH/MAEnEuAvNA1ldTk3lSe1GgTKKFvS/yHThoTnDFMHk+q5PKJa3uSgiiH93
d/GZ380PIlFG9IFka4EiLBpEXR3mKL7wA9y1HDesCpTHTTwCdabvHmOKsSFGHv5Y
miotPfF459oglh8fv9Hd1tOwlnWP8EcRQj1miQYNFuY7n7lO8qBI63KFDdKyw9u/
wkQfVo/dnIUj27VYSg42EcJmWisvcwmyNf8L/7pko3F6BT0jgxYiKLsQGQxuGnCp
xSohi5ash8cjcdQobYuMHJTLmX70dp5w5jzBw1wWw+RZRe9XhcZq4FxxUPxoXxoY
NJjd5jgJ/6EuacauSy8Bkwc6YIJf4kXyN5l0B4f+PKn7H55tEalC1kmthZRB+zbj
9mIMRiVPRQ9uz31AZiClUDuiQYwuRbgSb/5XPC0zl9OE5+W2JPp5riaylEr9eghQ
FGMTrsOaaKxktxH/Q1bbg5HTfNjTTQO+3LQ4+CpEcXbFJvnXMB/7Ps2fLWl+zWUg
A4Mctph/InDECt7ejGjT8hPVNJY/4xZTIIW5FgwTlIqio0rWpp8xYACpoQ5/vSvU
MrMfNMbGSMESndtTY409Mzacur7r5BW55piTi/7vuwXiQvQUcE+bvHhCJgi/uYpf
U2+WZ+U4Ks2Mq55jEhAbNPPk/f0bT9pkOMO0QLSArLa67azoFO2nWe1FnRLF1qD6
enu0rSoAjLBlPnbDaeva24pxXjgTfMkULc29v0NKr+l0KFq4lCDThBOP7TpmilcH
R3SzwEWi5vQchbt6my+7PaQ7hw1sx9rrkCn4ksHIb5ZrNKRo5ZkqhhjCwVT9bJzw
rxF9MQpX6Dl+3HPIPTScoUTWdFkRvXByL+w2eIUQCwnQiAT2VscVKBRs4crqT7Vg
/79eWkozzIprppFYeLfAkeokK+dxOnG6VJ99UTdOSXKhaojfn6P2OzXsDXwS6hEj
jTxCPLk6HaGomekYsPOfmbd5snEKzof06pSNy49txf0VSaBiJMpB+0Oeo1OPg3Wr
AHeA0wPFkAegccvPJg+DFy0jnYKd6iecoJTpt0M6DAJ/73WHU9RWy6j7Q4+rLGSD
RKqa5VctSdH5lP8ANpgl6pih6HxRVcYqLoRPa8R2/UBYI1qMJHElrwpTiuleLvPs
4bdRcqnQoBlZ1v2h41rGkcMm8r/xiRfGX0KsDpkIflbzOsXhqsLY6HTPUP9aFmbv
KD9qZ5aIDDtKULaDMZBOQ9lc6zz5NSbP/9F/rzZRovza1PWzKBjVSwOgFmRPizYd
mLNEHWQWYCDNwSAQtbW0j3aiaBLj26KueZE+lGSASPkKDKclhC98ylp0zLFgx90O
4Hleg46AzhwJP6tv7gtm+WCHwqXwUYZN15ZlLYQWJ3/l6qB2dIrMBYMhy5kLmMSU
eRNQCCGUDY3oqjQiPXBWJRA8xov65yF6oIAagokJbD3fy3xDNN8ezoFmOYofxd9u
ihwGisAd39frLlKr4seqA3ZhEA2tGqKan6raRiLe7CCz0CCWKZa3Ft8DEil7D7XN
UXg16ExCgM133lezQe4tM4cvWIii4TfYeDFN4BVDnTyyLTY2NOialIk4OgnlKJuR
iAiwLpPhNGiMHdYJzLAOEkGESU20JHV47Hew1UiOElOp3Y8tdNMBzPHJ1ma7djdL
FYYdqW9hbz9Lc3deyKqF/R7J9JHR/EqA7P12+0b+iJUGZZUfgFpo5PCwPf7LjoRL
s4jbNpHWmQFtGR/6+MHHRdU3PRML7ZrxdDhJdWFrDdmGTAhDyt6fjzUg0inzvAv/
c1nzYxubSgP77lJUK/PAHPaaMAaf38aep3PcxOwS/GnoxD4cDzxCZ2dze5m39jjC
BUjv2cY1Ttws40ZB+qvV/XN2uddAJcgCrin9PiUYeA7KRYo5qsJV1MVvlfdO+nUv
+lvfQBWWyuqHL6S5L0Br7RE4Rbn0J0PBctve5iUiW2RFFeRFkhHlJnGQEEoDI8Lg
H4qEceW8rm9gSXwjtZlNQT32Cr5qm4VIRewVsY9S5yq5hfMJ+OxQOQ+E3RoscqNT
OkvMU+MBFEFyUlQZOcQO0BdDRo+QME/L015bqwmRjOB+cJEgpFdMY3ycLmaJJlhp
6dKSEUDnyv7IhUCO0JBgADrhfKBdhKMQGUCx1mEUsfzRjKcEY/I4hjqQrDmP6spX
ZikQ3gZjNCEvn6dvT9whYFMC0JbRET/0PSsjEUGv9Z4k/AMhTzNmu54NypnHh1Wq
PztBhHJ+KC6T09OIUEAXNTRySRDM89U/Eda8YzSVibDEQGqivP9npa4dIoNXcrCz
hTg7HrmNU3q3ByyeFR81g6NA37t2Y/AsVhKJfdlScWSM/wbhmbNt3z92HYEvBknC
/kUrygmoJCxUafsnCzUE3Xo3C2LglidhE/mN5YSIDxZB/PYJkRhZSdu8M1gWBjWA
UDkoXcj/wiVx83AcAl1RTW91vvSOAdyqbqCZNpgBMEFnMwjWlOee5m6D5CQcaD8I
3d0cgoispdwveguWBtkLiNMwqbbzSxDjIYo+IqM8EpAACED25ndTGLmN4aFRyaU8
E+OTgXkyrDD2XUdnIHvoNTXBnxdJ5sPvxmGUlR9pD+7EJbbNEAWxIJkXv1VCe8Bb
ZN9y7yf77XSks2ouDiP/9kQPrLe/qgm4rXZ2Dx2IL068mugXqSy6SmLNM7LnaucX
4l9tSxyjeKzW/2I4957EG52W5tZzw7DPS5XMsrGIw1hmny+jD37aaI4e8U+9Bx5T
yw1/StEZypaKDdeOaVtX9DZHw+PNYySwwe3mp9zMDjIxtEsMIW2bGgVmeaTnmeiN
oVzegQCHFm+WdUHK8Sx6Zgck8Mzi+TDaDPDIKdY/BqA2V6U113Qzyo6O2ExEElFY
ssIxG8VFrwVe7UbqUnsTOwGs/5jbFygyHE64YGMe4PNWxYTP+4tSwSKn4Rnb21Xc
HUwNGw2f+BGlukK6fGS7ftxWpZC1lhVhnIHDolN/wzjAYXc1jRkuo+x1iurju9LO
7MzfWZQtn36S/sxvzUV0P7iVm9IgfAluxmRLnts1ze5K3k+pzqIQqOiDpVB43HqU
uftrg3lEWUajtqjiirXn5NL1GcvmuKQ5DXka0KKuGYM6gfvdgXnYOzFw1jfqdY/d
iryB0tGVcSfcvyDGvjgtrnaHLQPjCxh1sYNxnpTdrK6PmbpoP7fzbt+TItCzUehn
Kn3+G5KL/ep/dpkjCHl9ugYRvVSau47PLjRedfVLkn7Mwzh6lSrkgubTIzGZUsVr
7DYiw3PhTD0+L5Yny9h3qRiCfaKmuOVUhsp2eVVwEz2raOysCacxtxjIo64GVan8
xUQV2JY/thVdDQql+ryQClIEmU3EJMqDnOkcMyF5YKX6ohsM7mxMvxrW/YE7Bt0c
fWzAWZ3un9XrbTsybbB8KLVfolw7csRCZM0x3edOeQSP7US9o0Nx4698JGjoy7RT
VuJeb7p/7fIe33CNQ0xV4p+O/gNFW9Y2Mp4ATCXGnJKtbR/kh7AwkLjSNSNpfqPn
Np9bX11pYG19RA3WRRTWUKOKdXMJr9Jq6fpIRlQRL3VJQzxcWsstLoGda994L4n7
/M1mr7NCFJ62tRY1mDauMU2baGR0V3gPs8OmsYlNP9pqp7FJYdp9LvKxLHlglwVt
2dsUnlC2nzAiZoOBWvqJy0t838kGrPo+YrAHlKB/v8E/kcUsnGYcl/2hqpl4cAgQ
nc+o9PyF/FG07gr2qtFuLTfQ5iALODbxYYrln32Vk0kVybyZsusypQmZfFrGP7aI
4pa/BhX58DAKck9fo/FytZgIWGwZ/gkVDsyhNeGWGCP5ycLqMzWlT83Pe8ECHhq0
AI6tu85+iopZaHyYA/Oz0wdPVP2MqGfKoAlPVKLtpSGl2X1efj5KW4pHkqOXnuXk
Q+XusYwZg/wiYmrx1KDMZmY/36c85aWgPLbZE1iRlfCPAQe1fxPW8jXJJ7Yj/P+y
LRxNmpUJMpPkRy2gC77eJIYe5FxzU3gyYz73kghmGfSfmg5+qPxxba8UtVELN/u9
/tju5xx3pRpeQjeAYjPvevbzsb/YxrV2Eeyrtpbq1RgkChEunVZKYIZ5kMYdouJD
6VJJUydGlaMErUIp2MqoV2idqRSKlqYJIr8oGI2QqTcxoDtThWypFZpG9183vNbw
kQ1Un3CtgXtSgYWO8ZHkOzg4VTwB8g1CwSUreFvidUVwZY9LZKfP8fizORVXEYjX
g5fuMH1yKdhdLrKY6i7HIn51KPmXUdPGg+3W99fAoh4JFliTpwDPAoCwdHp41Csj
a2MM9DenBrMsWGvu4w8ObU8F7ePgd+1BUTVsx0kX6fFDhr+q3GoeGZNsq20aFZA9
x3e2Si6MdnzpSlaI0XATbn1nc+CY0qL2JgPiuAD2wHdLC3erUjut2iRVfX5brNaH
HL8Ye+KJdaPiK9daeasSAcCgwuAlcAbKOrGM+eYmz3FGUYBHETFAphhL6a2dISAn
Jlvb6ePyYGGmBxteHR7HYWiShUjL2Hk4xBRcLi02UQ1REiTcVjmkEVGpxF2Ga2UU
tF65XC3yTNaBNsWuUdvdIg+Uctg65DaWN6fQ7Ju/zeNEvN2EHA5E77kepw0lzHRK
fVorNM/aUxecohY6h+WVXCczgEYczgC5LBUk7vUpcR+MQBaoCeqisoAjvUVMPQcd
LVALgWSRpnsbnrbBkfgwLqKBiot9446Yrqo+EbGLlz8MXPWLixVL977mOI65048/
EIJN2XmpHX+kblTRwdo19jobgH/KzOLtqMmZ1Xv0q2vUu0RcPN5k9g9JCaCrE9H5
CltSGPJr3GH2RVSHFJ6qTiQvLdVCxPmOVmVwiNOMepCxtJvyCzo2HR+cT0ZWBgXa
XTfxNgUUtAaq7MPN5MMNaXhg1/yPhvLyC5NsxnyNp3xeGxSfvYfgwvtZkKcmUBYx
igMUK3I4T3saE/A8xP+3HE6JlSdTdOohJMM5TVo7z3uQMB6hvS7vk4e0jUrCI/3E
3eqdPgGelTQr4kiCHNfM6OBH3DlU+U3CslkCHbFSShfeGEv6uNgE8nifmihYYuYF
VhCmm2KG5+zDTJC3427BFQSI75T/tEwKtAJGKZiFeCWyhuToJCbb9TkijFEP67Wu
Ye1AzT17SC/lZ2ARNINejYf4uxs6guSXvhkpDoUqnn49qYAuFxGV7Cg5cI6I6mfN
Lv8gsJPewws40Cqnvqj+frpJ74TXZ91dBewPOBBuQJNKEMOM+zriIQDKfjYnKgH/
REmC1lXZ8/KejLHCS6T6wWxgnuHZ5ZbQFxcAoAkGyvFDD3W/drw9UKFx+8rFMZ8R
WHlEN4TuURVz6MSfdgd2LzcRKcn5xe+AgJbFcySsioNbB7r2zzKb8vF9EpI+HFCm
3N1ifTlLNbbUuKbb/N/CUg80ASBoilF0qacS57Drd8Xzg42KrC1R01B4Unj6wOUJ
wgM0PPGIfaux4HrgzCLOD1U00TSkpsUxQoaB9dhZJmkYBc3g/KJzA8dsXDNSrxRz
vMshFE58nnPaqCu2D49+wHCkK73JSxgaZjLEUI1w8eqAqVek2pcOt3LkqOFfiwYf
9A59/++FsUobRv+us1MPI9QoS0z1k4HdFoz1pA6bd1MmZwyLYtlASyShWXdcfDRj
vICaFk64ChC6+SQWlSgcsk5i5c7aMlMcWn40LqWtN0X5yoD1hCS+twxCS3ojLcuY
jBL6rCJtCIzym5R1ptn3Dlhm6rRfHP+0jMyNGV7EfahNwprlGbnxFrz+Q8TDfIZq
+4q6E5jWwXhvRa99pQeSBGeILTDKQCn28rn57j9TnZR/b1hionRdmlQQ2Sl6f83h
4HdNXxJqJmpKA17SxQ9gZ3WLzxIIlhbIWguVzoLf8Gq7l+c9CE6Jq7hXiaiFEWyk
+QL6UrsYdXgZXcMjFlbHwTe1wGt2LmGZwvmmSkYsmy1M/3D0v6R8xGkcPLIAmhZU
lsMWo2feADETNcM0uWihoA0e8aDDs/AuriXxXL8hTWi4Jk8zuO/aMZ7aCj+uI/my
Wsmvk8+i9NYzD9L9387KQxkzz4D7+ajHheclMeYQaWXbXYt3GX8fReRknr7O63HO
JG97DIZJpJ3RKWpB+dMhpm2N7q61kmrN+z/oAETTKlWrGyDfrYe6XHbAnReyByVi
Fu1Sg0WXXtclB5jaXC6vlml2laNCOG75Np86knvii6Xpcw6fRSScHdx50jCZSPeb
c5aM3ylhwm1tvR8a4x0mblOV7fNGIirKi2i4Np+olrPA5D14W31iF0r3SQvnGNyP
lCb5FBwbL+Tzj4C9MUetm2bUAaZVYwCl7oGJ0z8SctTOuhu8lmK5vqKP1NRdbNNv
6V4x5UBxyHwwUuPOafwjahrTC4Q2SROZAVzGf1rM9x/yTr1K7w+KHim990EwC7/9
H2sVI4+iOdIspOpNL8ENpBk3xs/eAJ0gE2XnXGjXpZ0lC00zpiuJpHH3Trxor2CY
qJCIRKCx5dAe3tt4gwlQb7wGviNI8uTQ5XR4gSPDqk6QFsc3+zV+fAAQnQgXLe7A
2Lr99TYzcYXNgGh5Ob24mUdnuUWFr+qr0Wvv9R1U1kc+LneTQGhElBfis1DYSmsk
y30GReMAqK1C8mCfzxS8jZyXis8C52n76ywO/ZhLxc7SS8Zv0WhTyhgbF8AnxOV5
jws2lbNVKz91F5qPDjMFQx6Vg1hF20MKVhWJ0zdfEwymm5SRGbyZK2sO7I21Jqb9
IJZFmBsZ8BmZtXliw8YlotcMo5H4pevqu7SrFAqrs7eDEC3nLvDXFqldbUXQUWII
NaBlcASg0hPcx+QP1fCqJGpxk5G+mdKO5kFzHXtsOQLLwZTg8mjcLiRPqMBTKp9y
zK8NYCVtRWmQclePF2IU0NW5bRMosqI67GKJCCpGyWA0gz0ltM68/F4ikEdDemU4
HpOg++4mnQoZYLmdmdJcb6Hmu8sS3f1rGjKUYbLnMc7aj1EVAb+ZuMHE46lTegCs
rix/2k+cDqAkGl4FCLF9UVu4UBiwujnZgNqMGfhTMELoZyW33OReLfuePoALvpPa
qfHEV3Kcr2wQ0ipQvHwjEQdbn7sy1dsK91GVzrpbm4K2zRt9Su53k+axwVsActHx
5KZIRYlnSREm3v6YxtaBlNulPNm4i50Lgyn+T/Y5cFvy8WeiRadh86RVDY0LjOLD
GJZblmFIoJ1dXHHrjxDXH3Bmn++YVULepguchi2pq/2GZPjM45vOJLwm6earpoMl
uq8LxLrHNsLKdhnva+qIZCuDGIBEkm72rWu6oS26PAA0kje+veOIgyOy5JH0MFi0
emVOPwGqu6Y8zoRpUiDxnDJ4KwpB4haIXQ4AtrMzXwhm4AiSzpJXGr12eCOGnIah
VyLDH/LehDqv/VPyYr6bM4Au/8y0bnzQGLL0Crf2V7Cgt9ZPzBjkOnfftycaWfWk
RKfubDxFXYzZTGpNjpmr5v0fkFNF0TgGQaSBez3Nfdx88wuLNzJgnNds4yetu7Rx
m8P9zRRpzbEaT8qS0j2jc1hZOcDaoUUXqPCxTx+g3Mv1MfIjgcQ4zadO8IHGpig4
k0AlyfKLSMS7aPEfue2vcxiu7BwtMenOOCyU5YXUzjqWOxoESgM8yYAU88oq+Rb3
qemdNpGvs9UsF4mbPiMJfp6KayCKmUWIKCekqGYBn/rVJb5niXBj7ZD3fsBz6dMK
BRlP5tg2RbwoQqcuNTLqQk3K44xAr11bYQHN5+rQ06/Apb93gvM7B1W3j5BgnGOa
/CoDQXECxlEnHH2PgiLuXU7T1o69w6FjekL8F40wjBwP+VxZ2dS1kshkr+/Ved1J
DVSAUlu2gtOFgMXUUaYa42dg7cp4qYfBA+9CL4vFHD2g6AcHYuTNwpPiKOmQNAzN
6HdAWKqJsQwZ5st4iPfX7Nx67v9jaVYjo1RT/w884EYsPnekw2X5VteM0joU4AYu
lx92wpJTkN3DPWi9dE8SrDP5rf5Xy3KLn2ozETkrRsWbqppHt+Q8vE5Qe0cByMNQ
T3W1LK9X1N9UxtJ0Ob4tqu66+EsutHRUjj6l1q0/P+/k6Abe7FfScM/u+XRZ1QwO
wSdSPJ8TvE6a2VB5doEM2xPuHIsdHWG3Br58HwqpvracEWm9Io/P8dNtv1x5gLUJ
l64NGBZpDsIgWiKQoK4Lz+CyqQ+BRfmMouxnfzRDtfsKji+8f9EtVa9URa2CmWv0
BHgjkt3Gq78J0GNW6HKMdSUEQe6hASWGRJdioO0v2aiqM4orzydb6bjfJAQi+cPN
u1ONS4adBGoCGxANqglqFVZyEci4zmh/ie3eP0TKzLFFhIbz1A0Z0fsPZz3L9Io4
dKGd4T67L1H3GMWILieifz7WnwWExGCeVbdDwRjwVuCOtSC0DXumBx0GvcfRZQ/+
mfrGImxqYAsFbOWiH9d9eE0BnH7S0d708800F0cirIJvBDg5H7IQFuxK4/+nP3SA
KAmZMyH56ZM0MvAcpxhQ0em562crVdIk0YvSgpsU1EcrCAw1eIFrQG6CNMedObEI
3l4owSZ8zL3Ehe2pNjcAKSULCPVIZ+gNjOVhBnXX3wBQsjPORMu/c8vNSWC0G5wV
4r3QeNiSNL6yehG7t7FFnw/h2nNQMboCfDq1q5zd1qlsNVTS3Q24bUx1iSVBtMc8
BCQLz5jtQaSvVPf4jbh4QJo9Tr/X2+hQ+sTVu1B9PdMPhyG2IcnAdFX0T5K5E9Vc
++jsoMcpvu83QDnuh539KgSBelDSyssQJhD1Lky5iu9/2abhPmZ1ZwAcGSCFH+vR
3OFzAeosZ008FJHkA9zB3PBzfX1nmWAaCvZR6z6iOfWmG7ANuu3AljM2tahvVQiK
Z0s5N9ZZoDJrp0FBIavSIhuSDhdib7rbz1eTrrnn4XNyI1FJEwJ+eZxAD0yU6TBu
2D82z5g0Z+Q2CZUlNfOKA1dTF7oht+i/JuSZQIXC5dNKrPCuhfg9eHeJ9F3lEhH+
BAY3Ym583Ve2hbXIl4lU71pe9asPvOlUur7fBimyJCfiym2MsGSXCCI1pV4w15+E
LYaFWEnp5AYHF9I29Bc455XXA1x68SrLizEacokOlNacUyGWGumlPhh0LrFU+RR8
NxuH+RrZbCKnFEwzIAYC0tOl72gwgimmuozDg6r4gdl+8H33TWauNcvlL+IEU+Gy
NxG3W69kMWE3Oq0rfFWxD2EyF7EX42D9yFlrHFWJossTaq9EpXlwkiT7cYixVXJB
j+5fp0nlXljsmiUKOWjh5dN6xrUqg1I6KaWAryvklWeFbJL2PUr9gX2Nn4mkXtgB
xX8lSjvYVwwjzCRxR0B2k2+P0UBNe1WWu9UPVbOO1F0Nd/vKqkUD0WLqjjGTYl19
/EAST77RuaXAUT20JYyLe37kQMivQ/sl7pG12knnliHyjBu5y8DF8nlsEcG5SEYU
XNMgdPn0MnSaCTNSRyzaIuz/bmG3mpCCCQss1Bo98mZnMCUp0yFe8u3tnt1VAgLK
PomttL5OCc7UKD/JpQ5JAsa4t8JfgygyikcOTUYKaZaM/kAUnKMZz9qbfvPSzT5P
bfJ+aG6WKOMNUDjMO39uXRmX4QVMQ9WMP8b5yrEv5Q9QAi7vS+NJO0hESHgmbbKE
MUVpycRQGFupZWVtSCOyULcfeXZYNc+zWrUUK8WyhpFOaMKqwSg2Di8d8pcczZuq
jekEx5VILqzYJgjNgjtseN8G+2j1vIj4E6NAshKupvrnz6sfmbv+5pi/hCIe4Pjv
Pg2B5/AJl/L79y6ToQLkTZs+3aOofFj8/kGUrGdq7GVvvWvbTZOijJbpfrMUa9WP
hPfdNondT7cAcGMFSX/OAs4V0Lm2ibNpilSvHsDQKAQdYHSB9OwYYQLcxof0gHrO
6/y6uvFkUQVUHAMiswteJ39x2JMcX7Fm2LNXMzI6ZyfEZqczdfKD1Oy4HFGvmLRk
eLsQLrejw18gnhn1EEajPxa6Z5eWcFk5fM4B5HA0QyYE0KFLfnrsDB+fNfWN19zb
gDkCO3wWR+2nw/QjdyOQsC5DWlZZhJUFj3RQ8Iy/10a9nTcSqSGCtpY8vsBBJHD0
OeY4vmex3hghR45p2CNs/TCoyox4/P/4jvOFVbp66KnWUDaqubX+1siSPimLosFy
Iv40IJ5oGYl/Jq5+6tOCaCRXftEq0s5kwoTh3hGuTa/fE/85QMSplFQBxS7TiKdT
uYocBBCqYOaHANcYqGcN/UeLvJXtmpzPnmk+ew3JJEivnWhj1g/PvXSlguDvB+gx
gYUmhTy+itQvshS2CIcigaSNhgZCOEUX1S2DWgaZ0PdUIhhtHEUqPyy78q5eSwrp
pS7kVYtSGg10Bc8wc+JuJye3zWrkaKn1NSx4bOyAiL6qzxLDggwfZatJ0AYMLDLv
Ars2URBZdwDPvIiHwwLpMalA8Z8vjDwRKUHEG2WA2PGgEV+D1C2C0EHriMiMWRJW
YM2qzlJCD3O2mGDxt5v0FTVUY7yjLhk3X8n+mRaS/ojAX7JNrbTk+EHxq6TBey4T
lUjJTEDCtZk8e9/URj2ewmJ1WZ5EfVjeo0FhOHMLFzZcY0Dk3YNFGIinHUzUik0q
9Ns8cKzsojQqnjA/XX3zKz+6+FuOOc9A/2iDPFE729BaixNsnBsRA2sKQZBV4hij
iJRSdXAFMi3mZXWf+pnIkKbooxLj+36GjMcYEoE9m1TWsCdkO7s62/6a6LtqubT5
c5vGTGGAwjihhgiLVE8EHAAfzYgD+OQdqykCatko2vjTL9qpKyxvoDIiDdbLjJi5
rhut/+Srs1iBOyMkNtjJlQS5lH5CkDTZBdm/xyYjK6SnJLaxfcSzG++cUsQjDcB5
D7MtHmInZz50lQeWBIRALzlSrF/lipvINNerlpidcPPxVXAJV9eJYyV6xiqQ4KZZ
voMes6TiSI5dRPrkfK6NzUa5uF6k8cPoUerzAS7OE8lki1JMSBYHA5zMFC0XLZIX
SmnnMJxeLs2s3oWLTL/53ZAupVfHZJjEtwyZXGlWWoceWy1zeHVX2PjR7Xf1tjFM
g7gSANE4QSYyCcv2fg87s/LhKLX/hKPy+by+AD+HoDmPrf1Toahvs7aNkZku1uAq
H2qlwv4WdJzXVZauDk8qJ4JefSCa6o/VIp1EoVWwzsSCYlaJvhFVtjM2lSF4DlcY
x5P17vB5pD20xgpyx8i5OofAoSsvt41Y5J0gK6Jp4W5mPKiDpTt3A2743PiukpZo
KWMbZbIGHDvoJy/I7ct2vkXEAxwrDbjYJEaLuRfK3qfFW4mMRaEGA5nAA7wouvY0
DI2HMoYISnquRDuKN8G/XcA1Cd0ViCXbR2++opMFm2yBpKkp2P6k8rAR8p5O9N/n
p1scIy8YMpJhnLs07+9nvo/oEHildehDD713mlNtHqDharRb0UNi59Ij+ZDLaicT
cDV03Jp/gz/rxl/KQhxuQYOp2R51/0q/40sX9EHk0eSwxmMKxkgAL+6sdBm87jhZ
6fb+PdPh8yK2PMwn63dCMhAnWttbApj4RvemLinBK7Q4Fag5qGiFsUv1CtebUKL+
dR8YjXv9O21Ho3lPqj+ppuGJMC2Y4rsNn8eDwyc9/KyFdbgrr2KOMTbiKiPLEUG6
jDlCyxrgwbDmnswslRFgTpE/u1QhRCn14lGHJf7KQ3Nib1j41X3x7djKwjc9QX/Y
qEEROQacMA0xowiEl0a/Zv74ErW6E+2qlNDMptq+MUCi5Pt85ID9JEUepI2RKRCy
GE3wPGoLHXsntDW+qawD9NYLTkAcXnA1pKqqMs4uQ50ex1Ot1zdGphkp0g0wYs/V
7Qd4BIX79vdPWtr3N8oN+cq/sfNhPsQctC70y8/EU9RBnKHKOCsqYHj8QDx+xwUT
ZZtufkAaO1NSCXyDGrS+V4RYiAI40jeqhFAAu8upN8LBwC/BVPFUtXSONoHloy91
aaqWxn6sJtJTUSIbWuF9q/XBJPfb+vXrrlyU3NTHRZc+lCx6ghYTf0orLr4GzUp8
xA0R0DvO/m8tVXpWoR+C82QeUusKmjjmVcd4m98Xck/MYHXYyDpBc29bJkJ1Cx8H
eIUmy+6FHiIGJhTuG0JnLGhMlLuvt+O+jL3Ur7R1ZT0gE7JYSq9BWd6te6gE052n
rpPphYmEAF9s024xyZzFg+aBHzb0/fjFHFsErgPy5iEsNzE1cMszPeLHYP2SjYuB
X0FOUgPaWsZkdHo7/1ALo0nnDjrNS5d+65zEsHFJLlO1c7eLW0Ga/1DbxxjraQ7B
mlva4BMk+ppYWBQ0poLL5DTxULhvGl+GWjRNe3tQwXpVOl6ex2Sr0WRjoLKcwV7B
UC66uXYIHTwpHmRrD0MWjqEM03vZHctrvk4pquTaPMXzaz3tpilOnXO/Uu3FBH4N
xBehGJoK2PTvIG/J+v/S3DTMEhkJXE5xMjCAZbp0aEloTpab6kb9yDjAIsQjFO8R
kPYITAIiuvTFWB9Q9uScJBBCPjyp/ArbC58h9HGq3xf6Uc9GQs47DE5XmT0O9DOn
75zNHtmUQud54T209iY30ywLPPl0CJJ+AJ+i8UMPMyRD+Zt267uVBOQtZAXzd2lB
rJsB2Wuj1HR1xtmzlMDlK2Vb2+7wTlSwQ+COEP6ei71mq0J8Dw9eeda1h8TrVssl
g/kmYT0E2V7cMsJc7XU+c3jFDQQT2QVhZSmvD7TGvoxH6WWF8iVy+jh0WhWLnHHK
DbtufltjfS3am9W0/b62JFjYoldkTw/kiBebBHwMGUUuF5zfoNnEmrHyot5+zXoc
eoy3p9vSPyqWhmnldvDlh6adqMRfBpbydouki+LP41emcDGMmZ8j0eK42AqzE1Uv
wfl09Cv3adoV8trXqq39xArFkzC9MOYc9dXt1kwFtX2vCiqe+rFHcoaAEv0wJSzN
JtMAd0XO/uOtd+RP7fnuQNPzQ0tzjPAmMfF48Odm+m6J+Pu5qK8PtthvYnF1RUAg
cWw9yClEc0XUE7K5qktOTsg3FPQNCrYllC3Ga7XIqEFRudQGr8T9vko27AmfGlAV
zxtYfU+T2a4RKrCHXPHD7N3CIljt1FcDLYMuTEsq+0tFYKN9wj9ZaQoE5ogSwyKT
N2Z912NgBQW4qg2tknfuFSY0uRkJ+mXb6F41qXvsQF53xyRYzN31gmuYm7wZD6eQ
juFZSnkABzAyrvzLLmQV9IClBJ6r5HMwl5i0i04AZwGo4ksAPnlebEn3q7mEvb2S
8tGZHiorofi8BQn6LlyQhzmRaosutJs6CDCVZJ2LYwrLx6jILkEJlMAMSIZ6x8xW
9JnigJTozQ07xIM3hZQoFS1rbc6V9sKduUVh49IJ2VSCFd6WL/rmZv9UaS3Qi8A4
70TVHhTWuct0prumY7kt/CZ4FgLM5YrLFLH8bWtQAN+shSDfIxH/tYDCFIxLWLSv
AjCwATZMRNXwpNj/DINI9G8IRR+/srBo1UTSgib54KnamUhe1eNZWNHHG3uWYXXT
QSWnv4FXBzGe0vmJrH4bDAC/VgMRTsV7kfGVd/xjkMt7D4lIG4KjIQjxHctUGcFP
SSTHQRlfw+moDponY9mlwjKmebK6jhulJaOMDSRwRth5MopIZMpYI2jXi6X3vyUg
9aXmqdgwf6aZv4YLwCCeMZ9TITcyK7RaVo0h5Y+e1FleAGA9Yblo++0KfyULtqx6
sREoX5G31t/xqJWRKpJoSmbbQV7JRKT33/DcRnjzb29YUIMd3kaVpIP4/6kzgjeg
ZWmA95aF0c6sbx0fFmeRSTmqIu/ek38xATNXNInzMdVe3YuHG6xlA4Im40UsfGIv
ZY2+gBaZAVKi/bitkKnTFx4a1FosAUuXtWri5HPbQ+RGJdwCvE1CEoZY1+Max22i
H7dqDsEUV43LLmfsyfYqynVUeeJGRkTpwRCgU1G6hkXbl66+Huy0eLe92iQDzkxc
zIYfXrCG3w+blAKczqYzQ8XuNhjkNzQ4Oc38R5mcSh3pwLg1OOwMcfU/f9QowAr/
ri8ikHbsYf14XA1bY4BZ0ii4Y9uqH0UEQpZb7ijsMc4GsKQF9Rhw+LKrwnHea9QR
Ggzf9oTSZgxr1d0v+xMLqqcqtv5l+w7aqBLCsBHudBTv0uB8DGuWQTKVZqCu4BWv
uclwQfu/jxsXDmxKSEAT9p/OA7j+3BtfqC0YWK3x4OUBPHfy9PXqw5JYH2/EoY9z
fji+8hbjnVyZt/iMzPShRPo7H/xnRvShLmoXTsuygQ2pEeEzOXqICvq4qcOOYKf6
nE0N20yboosz+m10PCclAg4X+Um/z9HjPUmOE1cvW1niP4Lnn0EsSlkmMTRbb91h
UCcxuF2BWb4iNmGqpfro2DO5OcyYY5L+YBLsYl+1iObxsUFZ9ScXuQMTVeUkAECS
BbGsJYHKHBdVHQzbDUrZWVkrAxShaMiIyEGQb536xQX6EpTKLo89VAqXNxZhmyQN
HhKX9WNWvqDuZaKQI63CrdJRyS2nTqeJLtN4KHFdesRL5zJtakEPNYzz4/RouqJt
ZKHhDma8TStGmcenlrHz+QPo2YrsAvML/gNT94i4ghSSSdJ9vdCilL/eAaib80hn
NwY52fOf9HoppG4YT23Th+1cAzS/32FVsM/eOa8k8VI1G3rVof1Fc3JWIp5ED9RA
vRSy1rrlGZGs2nCieBTlQ9J/fgSK23o3QBDIX5OaMg+IDPzqEH5tI4+CySjVlMs3
9dGFtD4H22gMq8FU/HvtXvP9oenfRzoj0/ZcrRihppCPqm7nkGgdQuKjnxVPUMzV
RE6NK3GwTK9W8JSvPgUiJWg/Dk3t6BfMCy5QiXdCRKMtQkM6Z9UFbwNKph0xh7Ip
yUThVNeGG10jcx0dz+H9MfpGDM2pmMXJw35dfymDFEIZDtCHxlGxiZ+JqYZ8Tt9g
Vf32FPSJg0rGNJmwUMzEv0043IIkDYsDB4+XsX8sdB3uLrnq5YRKg+nklqH47nFx
ookWVLgw11+eJ4OXHTmUinwgsWMf1RbgTHmrMss1O6yfro9SCpeXBWkIJ11bghSg
NkONMK77PZ0a1VGag8XrVZRmxiz22bYEIQ2EDLT2Nkijm++NUfUv/9nHtv1++o3x
YLA+p4rxH15iO0C5s5qugkpJQ5FG+ycbHKiAIovap0g5zqIOFT6QdJOXJs52EHzc
w2EFPDPRVGaei8x5Qo/qn4NAEsZFKrT+pWn2hfqghX6t+7vWagNhAYuZ6SeTZEcn
Gb4SCxZUivvkIiVhS9NhE/wSeaol++oARUXuC2GNFUZovo8Mv1C/YpSsbiP/kH+u
RieeERDbXB53y/6nKnzvvCXS4yO2MM45vzZYiF9AtLlBtean2VTULTjsV4zntzPf
KM9jVPS0IcWMIrM3RKMkRmB90ou1ATKYMuNO7GKfzJ42cFYiX8kOKGbQphogesC+
nZP7KWh4e5zUbj8sVdIaTlvQc6lUVh58pGBrbPeDeTZxffvb5yTXYqIeucErEcO/
JZsWJXbzD8Ei7bHg7wGP9lIPqg7BF3JklFh9PTz5eBgnsHMIpJpEnkwS5XJ3EgAU
cRQXG/sh2bPdqzeCrTJ5wpMqX9We1IkJUEJ0TkQROoUDKQl8wKmF3QHKb9Uk7gdI
zqiNFDZ/uvvdJJG860OTvyk2Wp9L7Cmgms8s1uhuUiFaW0DnLhNS/VpgQb+RwZ+M
92JswNPefE6nG0d2/qslO/E01J7LM3lBy8Fr+miTNL4WZp6YqiSnLRMwrlLXGeUv
9nmaCDSwQuY+n7KzjAQq5e+rIyfmKXy4pQc+ir9r0pRw9CG/1yNOdi6afWxiEAKk
i+4wWiyLXba8UicuIigOkoUQvaHmEFOnXtA8+bX2HmlhsJWTKCh5Cc8aOTs7g94J
w+YNOqamIjZb/Hy8498P4wtCNDjo93XsH4yCJYtf0Ppdl1rTwz7Egthz6uNENJUc
NffNYHzZuciJJsOU6rbn3kutgxcybI/mHIwqijcSKq0rP9Vda+XAQKy3xHbqtFO5
tE8UQt2xzQkGWmjuvBkiwlvUa2t3y7xflMmIXC8pslCw27zq1QBaAm/JW4vyd0Rd
pwLmzam5AFx7Kz9VV1rHvJrb4sd2a6sXJUF75oXHkEPI6e41wO4zS1NZcTaTAYIn
NC2mpXBHtx2KDh7LvzkWkam7b4lLpaANv7mQS5duRT4oi8o6aP+suHH0njvPdTu7
tZOEC8c4d9OaEfjwof1ebHFuWKsMQBclX/40zQU5t3rEFeNDN7Jax7nQX/mipky/
J/ta7x29ebqyz6MtD5m7USoQZfIfOJQwDmDJHcl5bG9kMMUl7OMt/RuTr218Q4M4
plw8C4g51bSZOX4AoBCW8UaQd/soX1/g7svjKJ/MhQVJpAXSSIOeYavqz9UK3y7/
kuw02mA2qyN89Ub+YNqIYVr61hYmjoE9NvSDvIrMjkd48AqAJk4gOf3cUqbPrBNE
k/F2ACA/kOwuiBMDIm9IepF4M0nDIknMGqFGW6fHRSvmYEfuGaMJ0YZ2A4TAr7m7
E6rcbuZozIoPzxRIDgOOuQr9QmC4PN6Zbm+HiaZWRKAVNaZUv40yuur05Y116myO
Q+ir8K4Asc6VkZK3Kd7wAdQ7ujNbLbYd5iBIWdcL8UbCu9EA+OzzALVXbrsrDlVj
f7t7InftM0+QScLyQVfwgyxUrQIZzCJ4Ft26e4jivK9LMnKPrZvoeV49EABMTxVl
Wladtp5gUHVAydG2Bqscfhg8iN84IBepBVRA8SGhvuvckzeSojq1k6Ey8VTeeVcW
/irUBUcw7ej6Qo6eyCwPA7qiKRH/5FRgCWi8cSvKObTLaFOPnyAMl4uVaEiAnBPV
OzNGAupS8TMs8Cl+czYllivS82w3GzJwHNKa5hwWgAzBu58S4/HzkH4m5HgkvOiK
qYoNRBkiO/dTtFu0lTvCeCoH/v08ZbT4oqsMX//B+2g2dNSBQJwkCpWxJP3Kp9QQ
wjr2ttS2pJoPKuBVNUgQTuTetL2cSdeQYUj53R6m8nHa8PojatUb3MMHBCjMho5U
E2vk83QhAxnv7n4nV99sNkDt3jNy+PBxv0sGFBdeUCh/cwTktFLditSlVlErkGjJ
a7+FB4FydN/f9g34TJ8tF8jHBtbSdTrS9XCh2QTbl6kfCKiNQbQIA4dt1IAjBoHe
RwSaus4748VSNL7CvD4fLdSwT1NZN7KZAnlNNywk4u19JV1P+Jn4kMaIK5/0VzBW
cNY6Hhp29JLftYvvUu1yivbvTfSm8v0me01eJv+K6CqSQlM/7jX3lyK5go7aPdpV
9MFHFyxmGF1mZOoe6a8StkCObphQ/kt4/51In8P6qrfHYfpM0qx6BJGsv1Xk9Zvl
V1jSkdES+2pKZ37pVDTNUcWkbgo+OnL3v5QuFW80tc25ywJvqZegD6plu38gBbs2
lG+7arxYSRm8iAze2PizzwSOqCNDWaJbDrSXyBlonA9KYYW8AGupg990s9b1evU3
wXQt9nWMPSWnnk0QhbT5zpXVTWcuPSqo4eMOgacKi9RNnDgAihQyFNvBOcbUufW4
oBLZ+302vdF3ZrFYdwH13ZV4OLkqbj8tYm/65WjeUaXMul0mvxsdlV1CiU8AcYpa
HBLWvVtZvaJdutUERnKYxAydaFf7UGYoGTEZQvBIyyvj4MHxVTK9X7LN1HXXiQ/Q
Q+F8IzAgPiAZE/4BES7j7bdXh5ELWKzXjqrLYzHwZty53iBO66f6uiwTECtC+tva
+wk/m3X62joC/zrWs41qC3CDWxj+x9rw7gJWEwVUX+MThZbZ2BQI3UFelkN6z3EN
cyO0b9Grpn77FZe86Ps8BRSQfU3lt8Oh6R6b2q8UQHfqaQLw1IV6PHnOODv+Nw7h
9+v2IuAPsr9pjKnGvXCFPy+e6+VvJ5fJq/j9zxrH/3nj2gz+f6oQUXlbh9/DtWox
7ppcxueTjbgGa5gGFEKarVLVu1RFnVNPKYST0sMjm4dLuG76j1WinXqdcO9mTC/y
ZkdmiQt3bOHljkP9BhmuOXY/kfRTg9U1TpgZY/em6Nzvsj3kQnPeqvZu1B8FJ9Rs
166zHsfXjnv/sFS8yJJsKuLEFWjFkvlE9+3yf5FMuqCVYsaoyKzU0hGBNUPPHZbH
U9Y3DQV2Fe4yNHCOrp7mi1N2OIAc7SZe1WeggiwUIt5qY2utRp/sDjGIEuW4Id22
y+R6Vola6HfnG2bq7+/wKN/rLSrLSVqR+eYTI1X1vGfekBJAcBWxY5KWyqmt3kOC
dIXETH3zJ0k5+0qMoWmKGYYQsI7ao0fxHJFiRqtWHjqWnYoHjqh16h0X4v5iLK+4
EghyXLWtdgmtYaqxG2YIr7PNeIV7QgVuP2QMnIbVsiuqDZ5XSA0t5rNvWyuwYBnj
oFvQN3qgWmA848zedCPwcN4sBbzJxmHVQ7Rg/OmYJqW2Exh8coF5F13FWt5Osopc
4VVIvQonWxJdfizH6LFPQAwdF5IOwBD1oLj8EIjWW2HubdVvAmPcBZH7OJc98cuu
4IxD3unaZ15glx4ar3565dqXwBqj9TRqB0qNTdN87cXN69nXIjn/JilfMnjJJFj6
+I6sCGU6B2GcelkaySu2rAFusSh+S2bdugjKFHZ/e4G9gzptUSkQ4CqJ8A+5vhn4
CWn+B1RSoA8c/6ReAkWIR9qnVwvH6ogGuzzDaNMq8XK0U/pDV0r4kqDyOel3bmZy
SKoULlNTUbHjiAjxEhjRDLyF4plQn3WwGtWk8KlKjUe2u3skK5mK8Ia+YlXbqR3X
GM7QmtwRjMrQqceEpTFdTiM/Xx5o7ACa76id1td2IrIFA7QBhvIF6h1phPe8lDJd
9JNNQi98XGEZJsf0xtRn2riP8xNZhUNKMUO/gzqZAEV05B7Kt9kubwzikXGo93jU
KVeXBE5/xPgF0x7li9EwlP0jDiA9EFUiEiQ+KHKViXOMwyPC6j3rH7vzealihJkd
8mIS/XAEdP9mOwKJQsWBH9eC1BZlIMHINPg6073Y4CpPS/nHmNpw29vul5reR4P6
Ve7qQINUYNhB3N0ddQWObrTB94ioiUpZTIWPWleGnjBMalyI9Ldawmr4GiT44KNl
SzAQjrvLw/qXOElxET3UX7dYdd2YAcBrhsl1n3L4rr+se8JPYP9Gi5WcCeN3ZNWs
wC864ZgAaJbcFW8h7m5UiEPxLZPFBig1GY08vADpSSCBpyL560ffrPETMj0ocdF2
+LFIJegTkppQqPywIiLHLZ7K16WUbo9lwkpeT/rKtSrLf5D874zFaYc24r2mmwMN
EJl2ps836aOobNRqazqnnQqBYZNmYJ2wRi3QaoIdMlb1Acd5YfAd6od54tQlenJH
yM6ijTjumV4PZEpPo1X7MCuAIOCrR0nzNJ/dshu7VMsetRe14R+T8lJWH4ShEtkg
Zb00rHPku0gPQnPaFBowS/tgUMn4rHwFSx+EnhQCGt7TeAYKIFqwE3liYKKnzEZ6
at+yneGgjjPO1vJAIWtwHYWQ2XH13qGrwFPUo++O7PEjfCxZvltREUhr3JxXZ4tP
GeeVhQBdjN/R2HT9ZLUxX258QaISoM7JkkL0agFq+QsloreEbUHKI4/2x4+pzDzi
VTz08Qed98MNbZpRkvmBJw4PmY1r4aP1LGdd+MaoGB3NnnRYFNqwF2MuqvlfO9Pg
hC+93rIkOu3FEkDvwverFoRbhMdbSB9FgNsy0M4n43Qhihmlq7BQfl67+fnz6/kR
BE/mvM0H4lSUWD264uAXiXmuMV9/yxMAEyLZlFdrMI6Hra8jfZ3DprucbRhinjjj
vb+APBI0IxL6t/nCr4UekUlos/mMvbWv4fBZ882Gys7QQnu4dpewGszaJ1iylSFH
ejdIz3Wb1dkZnEQA9Nb/MivGTgCktlH4Bnt0D1Cl1m7VPDpI9Bluzh5xWnMBjb/A
6lF7OpJGJtVtwzpiMKIuAd8kagj2A9CcuDzOGNbRsYxL60L09rSnNzC27AjLvITP
1gkhKcC3axTFN3oeB0NQ6VXa0SoKk18LgQ0vhCw5PPidT6853660e5wB4qECQmRI
TR+X/CH7YIIxiGJgI93TZoT2QkpUjBdpWcPJpfG3WhMsQZcpQKe+mhqd3Q3o5NM0
/MfSQWveLDPB7OgVd9YOb4wIMAc+5bbop6lI9iQ250OiTLziq8KI2iGIFWRQovSu
pe1evn0IpO28WEFTF7Me/L16PqoCFcnh6yFSFRp/6RPKupUV8MsNEJ1dK0q4/DXx
q6BkvmbWn7eCrNPEZocm2BMZ2MnZ/48VMy1Fzb16rdACbilM4FqThDC3KAS1MYhR
ym3xWhm4+fibjSdzzknzQpxorvjEr4Cqhrco3gu8FWJRTPymFIY9G6Jt1dmHR5Ln
0JdIdIE69f4mqTVSswUnSej8vonWrFoCXuDc9nm0F0zST5VGo0svo/nh8bRXAD4L
I4tKTiabh667YIyCVL/JNWFIc1+MZxggN8h94Vg7ZFYtXXecsfG34BwIb8SAPb2R
yLxyL5JIcie3DcMxHewMLFyCIJbehqGc8f4l6335JK9PnFn6mTYqhoxbBPLHTt6T
8ckzi2VQcqWrbnUEolPd8jK3kKFe0c5JudWdLBOsrIUWpn/7eqZ57+WX6bUH5kaE
nxRNtGtKMdtKcqrOEBH/ikbHZ3Zs/P17eJL3zaLfKVg/lb39vED6z4jFLRuyqGl8
bDf4ITaNUw3ZjTHpTh76j8sfyuRCm2vCwqGIPZU265uA6mrRQe9weXzHo4IXz8cG
qEyK98cKe2PJgjhYpERd5KwDIezZnNsBOZF0Sm4C0kWyjs/5RjrYE5/hG0rajWKe
103pJBC+W8ywzMlrh017/FOj837nrzvLWYYlpUZyPBIo1JkxqE/bdPm4I3A0rmEv
AsaymPkmT80JtA1fP7IQ/AwIIsz3lBzqJAaEacfNr08EAbyX7h4bwiQ90DuthhW6
rtgDoQoItjimThxVDB2d9EncEQqHPLCqGbiQc3djd4v574cUb+dyHq2ixPRtY8wF
88Pt4ibRxRZftzGOaJ+amiED74S/yHe9ehpMfdd81+dK7rFWlw01V1xeELm0JSYi
tE4ev+N5LGuhIxh2fnQjiWZTOg8knF6k1BM4ixhlG7uRacwjTeFByDg4msql3gqP
/KAg37xDhZISNtoBGtDoqxehueUm9VPpVrNKIy8LqGuCqikPxc1F8n0JmzlT2MTO
ebEad1zoz42e0ozFgZpNrHj25oESz0LgJXczGOsy7szVkLuyAImW3eDGao8OQeAw
qKiFxXlfnHjeHuP9wOpOdybcsncQRtr0N3F2L+Ftg2BFz85GPDMFBQUYKSetRGTR
TWkOhUFsEBl9nRo0XjiZbBi2G/oFxv8waAjbYqShMFNGnlaJwdFiRpDRXQihlpwA
uP9WfGRza0d56ADqPWYjt3ag2UtcLsAQK/m5XZosTIiIIlhDr1ccZSmEdcMNA4y1
3TBihaTPS9uq1Icl5ReH6oyG3GPEmqQpnDOavfzjZiDAVG49z7B4HVgz53OlZJWP
fV/knQXaraCB78YHCm875PPNz/yMcoBL8Ae9QQ4+19buhGOGs7sbjJu1M96ddNHE
ZrN09gimwSjPW1omu6U6A9p0RDDSbXhorkruBIOaKpnGFAV4UVej48Tj8b6qOlEf
SpJU51VsuO4aR/AYanU5NUFSSxoX5oIWYoorRTYj5Dleh8Kudsy80Rig0VOj0TDX
pm3b/WiHApCYoU5z/BqEZVY6ZqNaDJGCV10vQ+PhJR4vA0E/wRcaYuJiqxBXd5S7
K0iLDK2Nb5WsaC4Ox99xhTSmuTScmtsQhxUll+IdsbxqLSA7cr7m6Dl3sZBYU0sJ
knH/YvLAOWmXr/M5WMRn8ey1qVNnW9zkeawnzY+9vayyBBRPx29YaTiqYmWYip+4
BIL0n1/wRxARw20sUruu0wQbDZKPvbvZuycbCkWpd0zEvubHt+xs3i7PblMppMoG
uAoJxtxKvvjGVNLSGqhAuoe720ELYyg2txA224Dyx26Wph0153cf9pQu3EW+0tLZ
FQh3krRw1TnQjn3QbcOmtp2+eH8doQ3Lz/Tg7i4KmrVm5EFBERX0jjQ/EYnmNS95
AeOaOAULlBH5VGh5uvNxmjK/zzp7EQdgSDsnWE9+mIJC2IfPpdd5cEBBCJqb6WhG
EzCwa+c3w2c2Hzcvfgj0w7HaBFScShLNjBL+MxSz4AxHx5urMPSWrrxV7guMspq3
gVh9Qd8Ul796qN7pRvvp1vmpbWJ5C+h270n7g61uVXgxDcUorkvaRDd2uIgtPsyZ
LU/TvyA6+Qz/8P2KkTA0uVcZkQTTUbYNkRc6rkiXXrYQ4aahYFFfoNWPJuQ3jj3X
OhwgsY5g09mac8qpx59Q5R84PjC0W5j16FWq6s0O3G3hui2BwjDFBOA4RHGDaJqn
RHIOivDPR/gG+l2cCDfZwUqUFxip5/Ym3rPV1rS4nkDoBCBqwRm4E0MBxEsNrmZw
RlUw/9lu/vkKpBDT6VQ78s+brXzU3AcrONBu+ClqbDokTNlDWm8AOkNaG0lnjnvA
8RV2WJltnZTcqFnWQC0H+0KAf3A77vhHZCOp6KfQHy+qKCAO3lpP3lWHPwrXvNkE
qAg+WuddRLcZEN7aAbF855Y0nB/MzqEJCwS+V2n3NpsxKaqj3JZDICmZgRKOJsIr
HOQ9J2pRnvc6kgAkVg/Sk+sFJIKuJ8AWQ1KGQg+EDHRx3HtV4ayX31Cwzo/CwvLH
hZ3/2r0PZiBcgGpE2sewIuz1B3gI/quMdKkmYGfs2VgAmwZI9Qr74Z47Ikda3VND
tmSe5LWC+5C37IZhd3/AAH9MYPjSOBUCgYFZOaF2uLu8Cvhff6ZcytLImid1KD25
7Ylx5QDxEIv1G8JudSdOEfIS/s8AF6rPReApqFFEPTrahk6PZm/JzBIGztqHwixB
5I+FwFlgU9f58jqw2eeW6iyUH02OK/8+n/0b5TCenJ+YErYelS98UA/mlKU5Gnsr
l6gvXzI7oVbW0oKLWVctGX+k4m39WbFuIL9alSEd5sGwtrcIZ6EHCkxkiuwhIPmz
10PKNlYfdVsKBoceobrXEVli+SdSRLFKqXtau6LKKoSrHBuAslK4VZ5nvXf1yYGk
G5lWZ9Bfntq28XNS33LtmIadzGo+upJ6HYAjwqJ3aK/9ksigzjN2tBiEokuiQy+l
6FzLLKBI2q3ftPuwN6U3W6NcJpusoXtXgALUi1A49HJWBgs+Ea4njI3Qq8+NBewM
Zbhu1jo3nX7nKAT6W/fBjn7y+nZVMurzNdYPyI3TdziDecYMzFOtmgB0q1HdR9wR
7Ee3Pi2/o2Z9PAExoozee2UUjfOOdMn7pM/uxBriGdsxPLWtjGg5Q+BKvvSkco3b
nnoD/a+BlTReZIdjgiGRbh6KJiPkvaygMEidH30Ef5gVspNj5nOVta9DJk5xXC5M
7BWwnXhJcK3Out6+xbtCU1tWSkJ7CuJwjOdu6CAecoLHk5E1Y+rLWQBFSVWXcnKF
pl7ilJPYfo3GQEu6fhf54zaqghn2DjU9+qYgGsv6uWjzzwl6ftzxYyEyE0O+rsYe
+NG9Wj6p84wmxM1tTlhtP//Dm5gVMQlTnNKo+eV01L/DwAeQXQfrMZmpfQqDoZI5
LHAkbbawGMp1ibsCHI/9N/3pfO1yuqxk4hbCENJ6ugFpCQUWavmdjCD57xUOcdSM
vQs3FbrjbfuI0dUhisgQwzuys4HAY1twLBs447k2HPilgS6lb0Fh5/liZdtnwK40
X23wBUG8koeZkDwrNg3XSDWOjyKpd71IFKoTQfXMZrOm/Cl4Ak/TpX8xV6cgq4ot
55+Mqq6gGH9vIHAcqaz9O8nUAGvcif+H3ZMMeFBy5DTQvUrlSH7FQViI0kGoU7Jm
FY36zoxwIzVO2rDp5Ajw1BeKLNw2BNEQMkBfrt9upyJh8tROUUhwlIxd5FaGiO5M
3aVIk5M6vi/XACTMJhu0M7pYks0327i22IaUCUD29GO+VEfXGSXZde/GCwBPg163
V2v27MlW+WpPStmPtpdOMWl7pNtYppJ2OGDAcNEIKDERhvcRrCdPpxOghvUnME8a
iLHCIm0wBEeT80MeMKFOatXZQBV6/Nhvuf0YhAtBgXq+RkdyvPaAEi6lv6bhNmk+
8Zp11pysS7E5HKY3MjXGq1IIatmNAVH6pRVQzwDPs1eYhfHz51GxWFVRx7DnuqoQ
o8WGoW4cCIatEhV0vQRVOrqLY+ax3q8tEtGT599Whtwtroubi2J2v3KpL8LIxsoP
AZ6D4hc4KOOmoIxOAGh32VK2cDErQSWKXqEHLxazEqYvtkR5jT1X8PfzIr0uyCsB
IQsXtjjGzNIjkgWNRcpFb+V4XI+peuK2oiqyfS67lcES4sUJptLlOPguRLPVCWef
ilg4DsITCGvoaqiBYAaIxdqP9oLszzQg+SF7+5KJaxoiRmvEKmgKSR2nR14CqCBK
KqjfnpeBnzbFVzGQ67Umv4qXHW+fuqhtpvYTsgI7yCTe+GcKRK/GZAn79cY4OT19
ATy8p0nHUkeeHXRm6buvye13NFdIXTcVWgRNMdhw04+cHXu3vdPTLi1K7hLWUuOT
yemDFNVAl6ljEuQVEsWJIOiHH+TUW87W1snmQB48Hmxa6UyYB/w8T2h2dx0AfOHD
3+4eLokM+eV3z8L4zmtzSYS7EXJ25WmpSHG9d+E/uDUunn0Qgev89DDJc5VDvbJN
bmnhMoR9b6l7PYJUHQD+SJ6asZ8lnNiz/nfH5llRz/6FezW5XNxb5LCg69UUH082
nNpXDkPT1pOVnUr15y23q0EonXxp13vkcO4IaulskzPlJKJ34mUcodzc+HrIcJW2
Y+FYyWTC5+iEdVXo/nx2yA7e0/3PRBUE2bRVCXJbhSteRRXT8BOB4gGKhI7ky1e0
bfvWmb/jaC44nDQTfRGRRNFybuKshGgRYBsIkoVaUgEGvd+T6WMfG9cr5R7S7H1T
H6N2UeQ1VgXbJxS+O2xAqMKm5zQlbGYXWbCY5Ofc4EaJDwAwnkslCmoG3qfalh+9
rV0vKdLUmBG5hh2TWPtiS6tTi0Tqlwu3CCLZeFLv31gQBr1FFt50D9ZxorflzMbk
cXOBiGKes1z23aaYqDq9JURLYqjqV7RucyFzHd/iretM7ihnrMhZK0mIpekGjL+E
do/APOwlZD5O8QDerjJ2YDRc5DuuKIqtzZrywVJs+NmGgC4JUY6K+nSlY3u3HcAD
pq01jT3nObxPeggWI4LtgTr0ALRfE9pbSqN9bBO8pHFjEebnm92J2eggfRPahAjG
b0vu7k4znkD0w5KEV3+Y7eIxYRatTHmmsdIwPU4/j3g1SPagm+FZb4FoaM2wkTS6
rZA4l6q1Krusl7ji6qYVXMrKcVVn6MNRwYDOasznLlpjREoKil94Wo6VIdTtXQ4G
YedWmGHPU/ihGlhiLpdqNm1Rx584qnNFCrfdXEbSrM6kE0zJiXmDW4++leUMx0m3
YIKFZsObe1DN91Aph4DcplTUXQz5RIMrlM2u2I5NeCi/psSYvPfv3kWrW5nqXQKj
LjgseKh+7IngcDUhvybLZ3lEm5caJSsnkiqpCJGEFbTJd9QhrSPhLoDHWgqwtYjT
aQrAACKCsp0t4uWDE5m+qJMuPKOcEXCKKKpaJN7qeqX8ktKeWEc1aYqz9xxgf1xF
bIBT2+NAE7/a2GGShxFDhwzRcX3B6IJ2OcPxyzMxrasjnOvH4m9lIZKUZuZBGN+7
2o8E3UsdvUPP6fNlQ51uy8cddEaf1dfVVvO5NwzZQsdp807rvItHP3Y8EpJttQnD
SokA54lZLrzvFpa8kiQfa7zKTje0G0mwCmsrosStD5ei37IVCUAwK9XT2XUkCpun
JDubhR9ntsm1LCvrGbC8RdhCJCbGw8yXLBziZS1+0aCpEuW02gVJnFs6ltWq4dNy
7tcTBag/muVunSm0o6r36eCdITn4MOVBBNUF5pCqTaJlpSXfPrNgo539Np+D5hmg
i39VZ8aCJUx0VDyR+PEAg5gon+UBPQY/F/Bdx4AglTHg9VKsvB606u97iXNiFOPO
x98CPxpT9wzk2sRx0Bt8pPD4kSaNQ5T29mbnBVqxXU3GaCSw47LQk0+mQ8HtmKfm
GksNFIAwJnAHHCRxD+1+xHMfPWNo5nqpReNwfF6RUMd/OMJ7syqP4AAPoGoQGglN
E2vp495+93OG9rKO5Yz+mKuq9jNS+19YaFXuSIhbwB+WoF1/QO03oixiHcd9tp9x
qwyYBIKDb0DbNa/LsS2EGc2k4xizhGg5EcGJ5mK0geLrrB6L/laGfbr8XcRvkDhx
cdtmJFSYBCRcsEIn6lppboAe+Ll8Z/BFMxblzpGFkWYPzZfWoyiF0LBNO9UeDAm2
1xBnSpjfNSTreB6hj4lomNDiUu/THvDa6Xa7WnP5CRmBvYbrhpg+mQvQlQuNnxJq
qpm9Na7JrGRlTf9zrsT5/wlz/Hn13OXor+h6LjkallvK+oq7ZrSMCSZjvI8YXSC6
8Wqv8tEouVFgsD+8GuxhWwUkiVfwU71cqnlwKQwySnYxwtH8nHWjzxo/diikgPz0
7GpmM8ZnefP+SyFUav9u/mAd8yOW1kD1GlCCMpw5VTuCyV6qYzQEHzKreYVbLp//
GDJNUyTCjgMirC7Wa81udxXSChy9AcugVnvHIKWd4RKbQNCWkB17z6nArnIx8jsn
nZhbKapTtu2C1EV2hub+2SU+5dEsKQQYuyno4GRh2YLpRRxtbYGUh22aGHgEKa37
ZQpEzNhH2WUu+Czl3SwNuUyemFq4RySYz5J35FNTTnSafYf/PhUL6F3GlsNDuYHw
HcYBEuw2MWP9fp69ZPide3YamX7co2Wie1CVW8y5t3u0Y+SM/Thav9+onUYZuezS
FoDvNFGQbJ2ionlS2UdQKS7nPIajDc1JuvCpliKgKIXqv7gZpGU+Iro1v9kkk1VW
klclTbACaGIH+6ODOcwbuDfpRsN6DW8Ajn+ftz53C7KCz5jnP7EegFqCtA8uLz+g
0nPqcU0/I2upbjpREjV7wwAHgizXXQOwWMh0/2OA/oYq1ZFz8z+/RehxhN/tjmxS
mp2FNPs/XhIn2+sIW2nbbZM4Gq10RyUGSpQu4rQ4+zAz0YHrilmW3NmuIAt/4ewM
x75iMgP9HKSSSPjsm8YdIp4HlzXsUq6DP9sMgzr7Or0otS7Smwl9WHSZVingeOe2
g+iG73ya4I72Oxeks4Jf39iuselbrwC5xoea0N1PZl2M1gdLk+Lb+Kfn9NXZ2+eO
rG6Q3Mkh3i2HiXS/g7sELcGwdIRWGHp2yTB6D3rf6cR5v+2jzN6qiykwlGwu1Xxd
5dyP1XpbdbugG3OUjsjldQXgWLBdhsO+m9osgp91ePmHwuNVZVenpBTMvA9/TJm5
FFqIDmI/oBuP9Dz108ZpCwTRZt54M7RqUmepWSxYXE06oQqc72FuKx1AfdfFyBKz
AnPHY8a82tqV92KjHmE6rNiXyvqRycsahjiN9Y1aBmwPSa5341yp8dezjiDTj9vG
jYC7YIlGvHCBNUA9W0e1w5nC9gTTk5FoZYITLWwhoh0CmaLFrudayBYxtV5tHF98
mEHmMdkmfNJaXnN0mUzIFxZ17hDw/hkI1lH9u82vFF7ZsBapb3RWH9R9ddmwPeNt
ABW4IYwcehRNT3TjGKPbT+dYu2NFdBQ7Z8+Ck/xM2/P44Bp2q1QG0rY/ISAUPMX8
ikdDu6NeiIRpA0wY8jQS+sbgm1X0jTtASA8wGEq65qLFWTdaaPgIvw/Td61tLkMX
CuBByTGl+GRvM3Doe0176hwqk9+fPhxV1HFHFevI5ox283s3Ecdpx4H5p3eRywF3
qZLWZitfU2u88svM2g5S0xAGGguJ6d0BTuOeb6U4JBg/1xkiLi0fVbAGU7h8kQX1
svJuS1O57pc3HYbTjOCI22OHCKFqMH39ikENXfeNhQX3f9MOryc7RZmTTSqoKsxM
HmazDOGe9CnHB3TWIJogWxDpWMZ1wwOFaB1qfaylNid2m5lqIVK8bMN5qtzPuaQh
tVbuKjqOMzZYxfkYvPTuJ5DywwASCqDXxeMkBZ4W0czH/kzgpMhrtuhgIQE/UbqY
hXyuoHjdzHOHZaVDV0IZmwIc1UaX/t0g7DbWeNWVYZRfNInpqZY5gjEDEkh9oWmq
gYv/1KzydHEad3VWR1OaaUb3ObH8QfKaiFTgPbjdCEe/7V2wPyLe/0hp2G2R4M87
jCMHirkb+1maIaciueiW5Wpjn1IGl+cfMYhwfzOGpDRPu8kHhsId0LJLy6xHx9N5
4ZRWNsuVq+gi3/9XBCowU3LVZ10ETiQ8G9uDakjhxyOMYCKw2xmjf6enDH3pWLX4
jR3oUhYy0JKPywhad9iZx+5fk8ehZd6ltw4vUOXDsJSnICu4nDCsTcWy5fr3HKDK
/r7XPHdqhVKqigyX28DrpmtVEuyRjvIqtO/PYtkFoO9agZQgggRcVCUZxzvxvnN5
vhu8LarHbd/IoiV98/a8mmdxFGVS9+68RQSx9J2dLy32mRH3+VShEOs+4n7EikFh
4XKQ40WlPqPiPveimrkoQ24aY6IVZrrfyt6VptIds6cENx4QQPN9/oHanHx43e0n
Z4MVUv7Qp2NMWz45oUCAn8tCYfM/Y5e2lrt5YuQ//hx1qUc5WqK706fCEhr3j3Hn
deUezEutvYjNxq+3bv5DRp3O4Rb3ssKrC6q09IiAzuR1hWdSlkDnaMOjfO46WtqF
CT7dcUunbPcUPkzOiIZcRd2IAK9ER+drsiYs95S0GSDiWGp148dRrXSe0pcfMCSy
xRjWbIOm//dBNgHUTuTLvVHKWUTFuJS8GftduXbck/352A0gj4L4LAEBNExrxUI2
Y8qd9mjvHvBdvLFyPOFigruExiKT46THEIHeaSk7uHcFuCAWZ7QBJn+E265VPdxn
nbwiJW0mV/K5zvqW8yDwBLwHJR+2cr/l+iICUxx4WfGIoUDnHbtZruDcVRx16aWY
bBQ0hW9wwPXv4vjSGEd1HwK5Wyg7RSu0Mqgf4TxzUtdxuMNV0WH5sVcPCyhEjSVT
QdHk2ugWtWJm51wyVJ2j4NQUMBNIBhfo/eH8mTu8l1C9zmsKiRWJA6Iyp5hdVseU
jQVWjBXYdUtJdfYpvFBLN6bfOJ8yXjC0xWBu7WxJ++o/6QGPmPudw42T4dcjNkrA
R5chA+Uipaf7GjnNbBOw+sqdiK86Vzks4l/fw49hWszR4giYZb4KO1t3Fnroy5cO
8zLuEWWGeGgX0CBt0AJgScS67aakdqfSlxU8ea+EBoIT4GtgzM3JTevOS6oGox/v
CEg76k+nLZ48Ju2w80oUVsSp5XAeOXsKamQmmRdwZKyjQwgiyKNF2RAf7Q+DYei+
sM9yBV60Il5RgdXWrtwLqkp6wAnCaROhMHTNymYm5feDa1RMQJgz0qN4AeuK2Zld
IpTdCMgdtUge5JKgVAh8xXlo2LHvc2HnZwCvIcbrnyupKBMSeVo64HTkDEtzzjtR
o1UUGsbjCFngO+OdLUslMIPBDONLVUzWTyTCf7QHGS3xcLvLfob8NHOi5StySnhL
ho5z4YIjapUbqPCcR58J9rpD18Plb6Uf2i1qSak4+L2g0MTmV4GcZkjsD1l6gMP9
Mhz2p4Hkbb+NNd/4svWoROjKgc8lUgrEuAneyF/XvbYasQ+cdgGpaUx7bfIfRW0e
qOsOami0xg0H/8VtHH60PdRzbcsHCPdjW1xKeauFqg4wc9k8C228BOag7MQKggPh
0EM3N+yxo9PEBcZkVgenbY3vUC5+Fu7nRV3c9dRGW5jCqeIrDuQ4tI2T0y44F78d
l4twXqgIc9CMY2wTM98c1wz1mAGNNg5Zjuy4hDmIIJvLspwL7PpH/gfBDRWHn7xP
S+9ypeXlko5R4pjKJNHjXyQc/MztX0A/LQefo68muwIVK0P2AStBa7x8mPLRjGF7
g9ZwdzBTCxWpWXloUHLKIP7o3eSnZF0oXu9dJPj5X2k5cAkDv4CTAbkPTd8TswcJ
hSRp4+TnPWiJ09WIbMoIli8C0BQIgxWvt1K1I83BR4hQExz0baTkjUS5snjJkLEh
ogDOcReuQYH7gPUEXk/x200tSnoRAN0oaxdxW2MQYnh2403LTEPfQ6K3ArvnaGhq
g4MWc0/3lWcb+8/w0utcKIAutoao13mvBhMdcMO0Y+XbmG13RWSvY51HCg+S9nD2
oJanNPq3gJAoHkRV9q4sczyH/AQQ07FEvh1esbnNg5A9Z6gxQQfPlJd4jU04Zdnv
DPgEvnq9wpDDyhr7erdRIaX83pkEt8/zYLYeiT9AOmJP2aKI9zbKnrjHF/YLZ0nu
rf8ynPtwXNwwpWaOp7LnRAaUJ1EPUC2cEik0LnumxwC65Og6XM3pzdNeXH83uGUF
1YdINpm3xNc5DNzswrPONSa/hnGW79YLNRsKGk92qV0W7+f2dBLZpRkCIoCW+rzD
5paczfExOMYDI9ni3RXh0x44cyxdsj9H2L/C0hW2UVP8BFK2V7rHiPIJMc8gJUlR
WUHGFd+gWbey/U1mmfNPX3l1OU5FT5wryM5tGwwcVpeJw+hAWMzmkOVVVz2LDAyj
TUUt//QhYK10WWOi3UjiaKikmRvJIWNme+yW3zWr8uQYKiRiWaGhUewwFzQU5bpz
VEWfzFNJQy3+CnkFpVKQNz8xv214caOG98E6GxtByEGVelvcowK1kcq47Emp1/Wo
DBSgYDZ1Tx399oJwHoNdHWF4fZNTn6UZxcA5udl2ijJzwaKgriDznmi/CjTInrpj
Z2br6clGdvSx6NPKTzvPD3SvsnlHKhTgVuR2AjMq72Dd0XJo2e3BTFbW6NCoL9kE
Ucetqh8bYBwbasAgGvgBt2MEEJtOodtLLRUiDfUPhc4938pTVSbWA7HiuH9HySpm
qbPboOCoAmOHffuNEk1jp42UOYlNiOrYAIRT2GDP6JJrSt+nXM1OjUhhzyK6Mot/
JPBEZw86zY+DzNG9DKNHedErZtgGq6UDoHSevS8bkWpSd+GdaBQ2KwZfdAx7/i/Y
DQIyQRcwGWouhlwvmoyQwlpS16LnZJM99o6QGlnN3r6n79obDKbCLY9JUgcD0awj
ZkOxJtBkTM7zjxYBkMlRtGQpyGVQIqsgZIsG0XLmjLLDCXLnfR2D+YL9YfyWn4wR
023d2Me2VKBtAKMnVy6LRWtnyyQqnx2VwyFqr7jVWvK5Fn23uv64uV1LKH5hERTA
RUbEY4mc42zgZTY/VtkSYdVAgO4w2/FIr8W7dAlmQ2X6jzhSlyjMxq+mlOCkaMLe
l51hd7smjNt8AGmhH7G0I557jYcj3er4KhoU2Pnp9+bb4f6fgZnv6domtWMdARcy
p69jHoaFW6fBKrB8JWN8t4iEJ7ogjcipcg2BHSssA15mMC8XDQkT81omkkG7u63a
U7+RXgQkNmQjRggIuZB2nWk4S86d7Xq7jJr2QXJmnq9DXwPu/mgV+Dd6ajzZ39sf
t5Rig5FmAVOwXpg4dYG1DzQX5eKY3gtQ04OAXYXaKR6mA4zDuIikZr19QjVMp0+b
0N7QIVI5eXO+PQf96pT83X/sR588r8t8hMrUxuCcxB4gx+/mXGsKNiTGxHj+zCCf
f92IQQV4F4RvUxkPf8mYJmKzVbRwyJiduxug5WDhW3K0YEWlAm2KbTm/bavwOtSp
JLN1apxSt+rJCPYVGYqHgrcKN71QlNW4LPecIZudUlW58XKin+59rLwPycP2PCNk
bUTNxug8PtT3PmdI6YjQIIwuOz2QNCPFZ4HIDnWVlE2V4I43zigirNII4qXXrbr/
enG6Xmj7y04qvHoK4US5g3w1yvklUA8nGwxJ+IcARPzSpQA6Cc3Le7KC8KEUsyfF
gaMqCU7c3RE8hofBmSjgcvGY0TuE1Mr2Ks5I1TmxvWcfUzAbUeS0gwvlWum5X2OU
axJyUNzTvoxdpNI0tmv7h7P5ccg69zH+U1SsvjukgGu6BAIqpc4OUqzmgKtjOHFk
dNrudlWggjC2vS7//eEieTeyGdJNee29YM+x2+vxjI4iviYf/khkxF2pKJ8DPbLR
vttndAbMClKyLpFRn1On4IKg7sgSH3DhSirCz5B2qBrtwuWwlSgaoXgYNBJLm6Zr
apWREGdH+9C/1dwLCJy2H1jSVhLrE/+Gw4BXDvlLnBNZV9LluGSHO9nmCagSGV93
4sUfZ47ApigeQ1C2dhhrGiCNBCpxIeGmNASh7rrULTChbIohquKx87gWcVfU42lT
X91NK9utvHDTImC0ldZQv7/KPbwkwCkfR/n8Gtpz4JSjc+bPjFQ+8ib57ZEiaEFu
vRrqt+UZIjn411YixS/3vr3G2wsfWTktKZdEc6AoRyVGtzL5w8K2w+5I8dUPjnAO
CCO/am8tI7zyc4BoAyP0roGB6nHzpKjFt1su0UsMZWCplmnmmak6AU1NDtmuhjLv
/UP2NfeN2kXHK/8PBftsx5plQ6oWeN/iXHwxUTbMXEKohoqAPsIIvWtgnsW1Ip0f
h4MmkG7hCnykc+WpK031EOF4i+loFNCB99G28WmJgY/F5O2YDhPRRf0sEQKS5k0g
E5XtGDjEeVzp5eqREr4dXOXFSL+X3W/77pxpGXFZb5rMzziBphWnVHPbgfTNVswT
FuCWyg3ArbxflkV78oftxcq5BimhoKi0iBW32u+pgFbZvn0zLLQZyNAkVFk2cyZJ
MEb7F78FQ5CwivrSy96aEkTd857TE/hwt1wlry4dBm2avGdan9dSGGmgSwHI+XjF
FYO09cNJAo7cLd933GUygIExGUTZxwtny5L/qYm+2fd/lIrib1uidGOqBr18E+Gq
t/x96sZeUzZ+VC5HFmd12ruQTekMSMVHuGXbg8k4tRSoLNoNVXufo1lkYF4tdQuZ
Bf5V/bqE37vNhE1Jg9xMAispYefYCzkmJFpVkLmcauccZCUqKLTRi4XnGVev90NW
NMYJwKYaLuEt/H+qj1VXaHxiE6WHnGj2xjoSBmywLfemwKDi5uJ3WdYgdyWUhzbF
XhuDwNBvesRQV4jdljhyn5wMvcVKRtwPXQRSDKeCsrIZ5ovO81kR6hhQAULIvQWL
yXIEzx7c01MZCnLiZQXA2VOM+R2UqCOoeV4rnQDudtL+RJAqDxldNKIu4PwfS61h
K3eKOcGwR9xtEqSWHBFdKOR0GpXd5KD6XoOcYig5J+xfiBa4ZwlrscljHG/9jNZZ
zSkLtgchbMwf88CmNUVGi2Tb4CzA/RAH7lXmpbpkSEndrCPQ90BQDoYIsjFq/bXl
tRexqL6fgYze+7bV1m60vferFx64d3yHgD8R/Rayiu6o3uB6LwvJBmvpkPaACWye
qK4uLVLZJOryNyfsBOuVsaOOXy2AUBdS2sDlCBWmQ04bM04flqbX1HIOdKpVdj0B
qrw/Q5mtppydZ7zqYualacHdMWOt0D3jjPIKXhSC52RDSRNQ/xqKPd/0NxtmOuIE
eqVwZVFDszfAT6pNCm/S4GhRoVPTzQGsXycoATUUPSCzjHd+z46LRn9ZggSrvWZm
g+xPc6iKY1pjq0HKp8//ZDQYXWSYBZcPnWZwaNkengvBBc8/g8LgOf1RYPwQDaYY
xPV7l2G0NSyEHVf8oXZCY9w8LxZSnd+s9v2hstoUU4PTkN1EdR6LsjD1wQBjrvvZ
fhBMt78ajuem520iKrsbtOFxiKT+8NysnA+7SYEpFVVvQMTtSGZ8HOfO0Kq/gyvh
kpanQBW/qcs6nzQ3J81veavUIn2GCHeA0zz7Xe4ecaVWllI2Dx262R2EbG7eBUmU
Dsq5CTCVkxo+bzeE1lDFTC5NRHJwdclOZG+CKhdi2OVTMQqSdtfQSgb/7yzHtJwd
WskJlVVsMPn4MHl6+N/ePxDljGkqpZHx9MOJkX6yBLkHKOQMN9RAnURx3P3OMP8d
APV9JPcxtn48xtdGlQg8ZqXuGwCv3EDV8iurm1iOhAW9wNGEnWjvGvlwm2rrppIn
N/nYkMAZRWz9UH8hWJHAwHELDciO4IGmpYl28sDDXPUl9gCps2bXMT5MqAhm5n7l
8FNr65baF4kbG6XTrV3mzAQX3DDAQGkSpcoG/bIRRCdgwX325kRCaOReEguUpKxS
Gj/M8reUKBuOE3jTdSpTns/ntab2b1gzp04BERmj0rr6YBKPjJsKVNSejCZhYkYK
jT2pYNcdvFfg104RF6xvjOO3/AOtjJaJTuz2+lUTuDaVVfBFH8sLgxs/0i7keigL
hmd8Q8m7q6KmqqaYv6ERhMKAuFWTgkDdQOYZN/e3cy7/U7nFKvakm3ETnoltojob
xk9P4UL5UMYSGeE3UjA+jFfrQ1h6UWxDP9FjiVwTqOZYVnq1ocr+b9G4fTJIuLTy
vVIFfZMF9CtdDs/CQopKHvTyspbTf+ois8gi10PkY/1bZ3ztdGMBskPoPQyyA2oJ
OjSvVGMHvTS/fTmcmgCiySBLP+qOPOBxv3v0CK3tZpVtMP7D/YKnaD2ic/UsXb9U
jvHYEWyY3sKi9yjdj9ONXCo0CuyrdL0fRgWOUlRZBKaV0P+/G476Hoz8eRGTp4Jl
dc8H0rwr7uDbpwOPJVmW9ytOFgYFazK4QFstBa3DWGH08uLF0E7PHrIoZYKg2xMF
LFTbid+ZH7Ik6LGO+nRhwPMUGrVMcy6L7W/niwjgRgs9GyguEUgbQRGalDHPNlga
ZlcMJMlfBQKywy3d+tBbiafvf849QX9QkVe9yA6jgUPUZlIK4bBOYUfNum3RNlP/
hX6E5jIse80gCcHe/H89wJ5AKEwUK8GIQiPn/g9i57yPoRHCxcSVK7AxafRT83Rb
Hx6cNEbxN/ADe0zhuv1+3fPATOzsa4GY4gvmTlw1suV8rIYQrRg6vU0UT4a9jUOx
pI1Yqzq/QchmL3iT3Ko6M2k6TE4bNHJCCQl3Ng3iS3RdGIEO8DVc8P1cd24qqZee
fLnMxRhYkc7vDHAMxoNKyfHY1HDNNo5TAIvTxsA7Ty/Kpk2SxZoyaW2dzvwEZltH
Ur+ip2kFgMANvf9FCWeeSBXqG2DZxGN9jqJB9lahc6TgMkJukpTBz0FMvUk7fWXM
SpECve08pOhcss0MKjD0yysZB7Ga8b0apgfi4OrDOspeNmpu8J2yUw1uVZvgYKKR
+6u7n9gafRN4RH3dNqwlI+2GTn2eEVLuMC4WoChdZF3/wTRe5elEKPbHH/Uees+1
EEkLoAxIg6Ov/yvwjALt2UZtAMvUJ0Iy1xNL/VEU+OpN0giv44vf0gnE31GCYTpa
M5G6wwe8St143OoDCQW873VYqqlNgsIaDkhTG1Rsjhk3m2yUZST6y9wStMopylFf
dZJqcNUPbbQYYsmlhL6VG59WhXjG/fWOorae28ImACiT8k+ZoknKir5Ce8CPuqwQ
e0Eo3p9iVSUkeKjH+bE+3jhP0pjCaSihwo29DLlWAvDhnZA70Uq2BbERnDm+3g9y
Q4+vINybaQvIob2iYRT1Z+DRJ92nMMKyv71Mm3QamNISVc3wlQTalEeEK+m2s58g
oPaEIWzDV22hzPH4r4eDvTv2ifbMl9x5k0pLVWIZvottRJXsXLol351UfsQQIjnq
VtTS4MYEsKfxp09PCJiciOdAusQYDxKfwagy4d5cYNXAWh2jX7yJ+Vvpi0gpMAKQ
LnVPmqnTFJ9IH/c7nLI8A+gaL832kvhh1v+CSZcu+/9aOiCJx8txxQLiNy/9Wbxd
n4VvGA6JOuGNn1mANuUSYJGIHijBrqtJcjiz5tv7CydQ6KAkXXaN3csmjGmPc1U8
lxnQXPecrSsTGprVNPWHppNnAbEGdsl3gqO1KuFOJAtSVIwvrlyID8XmX6z6Y6bf
kx2Rr4CE3aUKUVum3oMRQI6eehGkXGMN9uCSRRnksi4cDR+v8kFfKbVhV8D9Szz5
fv66j3redvJaBjBuIfl1AqwrKMExJ5JiNar6WO8L6adDi0FR2Zl5jBje8QuRZKvR
5THnNnm7GP9Yorao0qwz6SvogeNnBDTewsKpLDibtlMNgIc3zvmYKME/HYRuguVU
27+pV5Po5KPMl7G5US1CnWkgzhDR7AIWPYR5+tjjwCU+r/eK5Rzffrm7zvf1NHRN
htsTu3jjc7eDFE2zh1tTko+264JNBjwgmvYCKY20KK8APO939sALSd2lTlAu8MvR
7qXSq1tBEXbXhVDc+wIfbkLH874Vbh2ZILfms7q5QEYWpFloOoaDplzcVL7W3RaW
i7VmoJGUqqhQX2K/q6qdOgdllX0wrJsFrB6V23e0ZzF6HPhIKR/sJxLtC7HSF8Oe
sfqmmudiGEuzIHN1EF97wvNB8/iG2gO+Fu/KKW8HDwX0PtZD5+KOlfhfVfEP5b+X
2a9E7zMt1VSpiM+JfkYVIG97KP5/TO+dUs8aOIbU+ydo+QwFdbJDiOmFZOrLrQV5
eShlnXO1maclylJLnCz+dyD/48now3gh/3Khshn55L0AVWexs6idaWuMJGdfDkNW
N4W1HPTyMIBIMnhoJ2IoUB1uJgylraSI+D+ZkQQlGWR7h2KZU3QjO/ujyFTYinq9
MP2NP8Jc5KCDlDYzH7qWKY0R44QgoivYhFGTb8SUFff8SuoON/42LYxNsm5iDX+i
72+lUx/lq9PDFC7alb4e4aLrna/ONbUuemOFR4ukAoqlkQRQ0dLVgMhgG0Fkdrlw
lkGrCUupnuk86MxVyfdNkSVVJjdkFau5nN+Qsf7kdLsxwLQojBnnquYFKEoUr3l3
747AeRtp/PkaXXBNDN2VpIg7zO6/Ww8SZlfdDunbpJJwDPgbcnqEwhq8Jj98eonv
cD6vjJLq5Nj7y+aKaOrAWbVQGzl9GDSmKXX1e0e9liAD2EdfQlRWpc4gbuGh7Ult
kD9IQg0cwaMzxzK9vdaDm/MZb8QceXHwhg+KAPXMEB99aIt7tQ8hBPQhCI7PNztL
RzokXGgX/Ss+Jsr8Z7Ii4mCsJ/bxRSI67SFHPRaFptzXANw247Hm1xAq76PPV8Y4
JqFoUE9nEed68zUUvnSTYWQe9DcuchTjfQDmyHPBmiP2bQgVLzH1rvnCy3F0VBWV
EqjR0eilW7nYTorXqzd+3GV8380guPX4kKBRIvEffvEUphX5435wgB+1AQ4Nc+Z6
oRwWPx6InsnSGSD24lDMdw3XbwYEM8oO0nlJkf/qj4E26iuTYxckG0QXCZw0knni
o35dJC3cftVQrHcGOYT8Kqm4xAE+7e2Iz3MTjohSicaOofvCWsibCE2lzGYNIO0e
E6G0XctUZo/oFcHj/5114RH5tlGiC5aoShuE8IYOzsLP0NofY55GOmtaSdfsl7bc
t3/dUYSmiEYsjEjI2LC1j1jCY3QsGuUOYanrNLn/XsfXhQ6ftXw5eqC2xxworGed
Nb60SpNmiG/yqOu8OAxSjKzP5Lm8Us6+8/KfBOrGEeagmzRwWlPdEI3elCqVw9qM
JovJvWUeO5rS+GL2+AN+K3CmOK1VRnL30/XNW54Wa6oKKvx4vnxOqvjsMdVbOAyk
RIcazpMLOGYC/7sLn8ukTvhdZBjOSSDHTM5s2SOjJIw2E006F+5KmXQ+JuJlzW8+
jLcgdXWDHdmyg1d2C+VXyjyTwPdXjDLj/+k+F5SK6P4008zJWsvaPQSSJDS4z8JR
Lz0cIstQW5L+y5BKMaIuLg8svXDgNXb1TQnG+j0ydGYZ2dYTW4sHQXm4fYh2nsIv
UtrNyfSpohMkHXJm0vakQX2Tdoe2SWUyb94XOtdhAXIgsf14LpQ1+CJP3WDg6dvb
+f3weXRma0nbYC9VMKOLFqAjLx/UO9zk+vLyX2TLrAE3OKSyWTnEycvwbLrqZcp5
aCQpxe0lKZzBoFNdYpn6yWSiruxxADbM/Wzxh1cu7xZk7c0wbvJCBUSsh5EMbdf6
on5w31c0/JGx3mOkgURSwNo00tQ7aHlf2sesIPXFVLzx4ekKZqzMTTJICbWTNysF
oQ9yvMUUQT0kNyRPfI1+8+HnbJQiOt6BwmHEROF71WKrZN/l5Nu1AFddZxkQZLke
L6c208fGeeqOWSfL/lSGVGwoikc8/MHRJKL4JLli5onFtVQl8gqpkdyiRlzLOaav
XGqIBbRVeBkBpasaDVe9qnk8zHAmDCg6bcQxtaNB2z6TAPGh4A6SxjFlsFSh5OLU
9pQzsvRCmkmTTmbugX8UgSdnaxctI7ulYNJnrhGIgvJnTs8/Rdysnpd5xrCiNu/m
YBn+OPCIZN5q22rytoZVGT2wV7UGGal/vS/iAaFeAa0KkaVl82uE+LwkjN1Ltvwt
Bb/FFCorPghdBLYkUSTskH9QX7/X+fUdsw8Fc7Ut7aRaZQKNd7wyzKu2vmHg2Q+h
XiY3fRCPUr0XApB/lMVGGfP3drhxj7ayJIK3WjNscpictnxxvtwyHlg+KbYDBS6K
GoMTkmfQ8xGh/cMm09XX1MtTm0GNZFGskAHksZJHBwZRovrTYA0OrUm/MRzkTcPU
tGWvoe80ekab9RkSfRNwBA3V11UXHgeOuA3fYz4GF4cGR7uFHOJzm9Mo8NR6jZKQ
bzx1zbV8X9CgJUHLlY+8sgi7FOdN4vauskolYkP5OCVUSnJypLPugC5j20nvv8UB
VH4xV+YCJtkymOtuMUYApFjt/btFQer6FxhpxB1IF3IS4NhQ1rMD61BQ3v1/AfMA
aqfyGvPtHCP8zRJvqpe45oLeGcFUBq+5rrkbZhGzS4GYg2nfsQfeLmc7faaTZnc/
YhyBql+wxvldTxrA3vomw1lsyUnU/pNKl7cppWG8suMwWPiozZHQBv/9aevk61M9
tWM2FPDLEs+fop8ZPBGufc5bh2EsLtHgK99BvZSjWrErenYz8ZfqCESpCLY8Eoel
vOcDG0ral5Q7BtZVKbnpNWMiZVhB7tNK8WwTuEyAXDNv3nbalplPJ672O4JdqMaJ
dUPVE//0IJBGoxEQqXjFlx01XhF8Zwzt8loivS1N1YtPv1p3lr5uuz4NFcE83CdZ
5iiYJ//ZEBCvfXjVkKiUtNm7BnjC2maMMvBxSicpJ7MkrvvZ65pmcAIIhwB+2yu0
nZMYYAS3HKB8pnLxxctCqEdulvhsZQssupoMZ19fYEUZbBFp5pPoGf03wBD/YNcM
EzwH1Pe2LA3cvErW0idBjy8nRBMEpMhn6lmvzJen8FDnk5+lj0QWEUBRayrYNTIL
4GSOAbZIiwSak5fALV7uJPZ2k6xP2FwpmHal0vnFdC7jFiSIaXn6sVg0j014aVz8
yakJiqgqEpgIEWvK7C3d6TDhbmXbX7QJU3NOfTNj6Job47K+2wsgI7vrokZzeaNU
rMhAY9pvaNcZvrJ3wdouerN6mHQlKJlpb41DUxAC9KkuIIclNUF6IqAnf4U2h1z8
rs0GXwy3YxRoOrjJoc5BMckmyGC2agJayBkV3+5EBYavhx2phdKhx2zT6ChbHKU3
N5oCC4+D1O8enFYWZIPD7b/1B7CQrrJJFWo6VeUGH5gW66lwgDXKnHYkHbgEIsUO
mRascHwm7XROZM9BaqenAS8ailo7LCrTqQiV9lliqSelYTjpqqUnDMHRycTMXS+8
TAmGVB+EPmTP/q/LiK+DRpEW+K3Q2d1XjzBvuwJPNWBotyqpFIC6roXs8APxdNwo
haBIvR2vmeuqSUSMayToBK8ZzlAqdP8EkLbqf9TsN7qRIH1RofqysEyTbRDMt0/4
hq88MyrBZO4N0jTD2nx0uou4fNNKTFoh34cIzqK5sVMaMJgaPnpxXp8jSDTgFbcM
1RAEHzJ8sFKopRLj6+l6739SJyOsGpzH9t317kkdmDXpfZukEyTp4d06YSKxWEcb
DwF7Ulp8W0WhhBWuOO3ZS/8dvFr4CeVdV7l42AcuYSut3Lx2YiO+2tt+c/FOfH0d
Sh7WjKnSiS+SBGvELgHhj0yOgcUY9WrrD7y0PfmiohJiTbT/lV+zW3B6tYCljP2V
HPvbfk3Lptn8uhjAM+pG8UfwB+NSZw3AvoRwQ/zVjt7YOPVOVi1QIhRMykEJWYzf
4uRA1Z79idtM/GWg1x99RQVSfWkaF5ih5mLjBp1fuUFCyv5mQeIcMEheqR/JccRq
K1sGJBBoUOv64kNlx9CIXG88ck4EHYQOhpIPdSHyA68gUaApJQSF+pO5VXRpLs3e
XvuoLuH0SLVKQB3lEYDv0fANfh3UpohbRdfAlEY+YASH6oJveCkkUPxFjiAxQ3pq
vMgjYVpjwiFOkTn+X1Y0XirME/ZP7mGycEpFTjuwgOhyVK63lnEojHB8I55jb677
LuEy+lWu5XzvYf6tEvBcjv4wWFQvEE/N6b9/MKRz6iMfS2qLjvMcWhUgqHa32M4D
qIA2cLsJmWmdfi7w211SDP+wExOO6I8+6Bsjv1RuzUJQ/5j5fw+4XXK1xjVeG3eq
/JmlhjM+4XMDH4KSF00CWPNZnroAOl/zIyLnhG2AVTbvlejvQe4foVEwxUqCwdH8
UXYmi61XY86AfznbqfyYJ4KOOzOHVN60if+RgE3XoPLRr+ollXNUh0WgnOlmwFAE
PPQsDbmhDCAfjdBHqxHYPOJdXyNnDzdPGPtoIr4Zbp0BVw3cTgU8nbubXZiUus3/
6BUL1e1ykOCqBtCP/uSFI5tHhAuBFk2W8GTXNQezlFsgteag7nRRdzhf1sfcq8dF
qF035GmasXrSpxPbh3NxBkmxPPRHEp8iVouPxPivBKsSSBMXaCNNFf6u9lgiMSQY
WBbx1cb6+9UBzrBbUWWJ+2JeqeaLxo07YUCAGEiA+j8YyYYcBz8Ri64HnBf+FSMm
Yt94YA6rvneV/f/9Kb0/SRk2olE9glAA5Fjj2PVazY11cuK7Gt8yMPT9MrPMgKpT
4GVHyDfWnFgrmdxUrF+3kPfkhq6zopZsDyah/YlbPLa9ci77A57wqmoU6YPO7mTw
omGhQrt8Xnt5AFZzYGujI2QHRuLf4/YERomz3G3OslhTWie77+mZqC1qHlBTKBiq
GkAvo8VPUnyeDtjHBURp+Ba03ntDXTHEzX8ie4X+UNpo2m/PZGKYhpFYx3BLlwl+
paK9qEnsazTajZAIOAAFnncmVLXt4y7/pImEvk2T4lClyX8678RTrGQ63h+KiTtQ
8Vw9RE0sHrQliD/LUEXWkAvEYt0TAfwTBHB+CpTYxA8/OEo9F3rs2cQqfWp4Nlb8
mzMunB/ZZuhkWGbBThnZFg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U79cKD2AdTBp9u6T8MCSC51794EOwHrFUaoLyyhywsfro9USVSKgDXPDzZOA48B4
pGsFvA0Cix8UY0nv0vgMNBmjvd/F2lGzzRWUeS3ee9cYEdSsUtTcBr365bLQV8By
XJtdbODV9OLa9OisrZUZ4Lk87CWslhVE6AAvB2eM9pOoSfUgZqvQw2K6acL1Nc1Z
SZv+kj8KZtu6E3tLFZ8aDnIMqgSaHwJtsahy+7+ru2CzsVZCptRlldd0/6KwFgJZ
RldvJhqkIYXcmEF/j671U2MSZYNM6icYhDBZiL692lQCez+r7IxZKwljwa65gMK1
X4cQ88clYW63mL1YAcNckva8w3VaGYNzjY6uwN3zLLsRgPt/cVZsskrqebbMBTZQ
vfOiAkdopiSdkBiDL5YpOJsWGhDDShr+7jgCvBhlvOIgbexoHsZZeZolNn34YjZN
Pwn3OCX/fIgEl1Ahtvv64A==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r6wYfXGe77xzxs5iI/EWukwlogfjo5/lQSJhW8EfVDeQ8eb9XZRFwKxm9aNB7nyM
OFh4NC1p8yOqNslFXDyRGUyPvrvck1exzZKDVhcdaIa67wZ6oJOE1erMmG5mVjdA
OssRLaleOPHgxuz2rdEs7zGM6lYqxnpb4at3Mzwxj0rU5Kd82/Z+wf7NCxaRkJBB
QWTIrtGoo5aPRO66Ksz1GMZh3l2Vit59eHOExfHbDaqU0mxe8SIsiON+CIaVCha4
Yw2UqtrXyKjgvLU8AONPb74DGUFz6pu0MegISj7u8Grzs/ckJNflXVB3LKw34YpT
YvCGA+W6ey0xrt7tDs04QGSUDOpL6KlWk38EL4hF7cFEY215v3PxNBi/0ripWVC+
8nDNflQCZq9u7xKHtLYro9yBXSUO9MuSz4I/ri2jRr1/lW3Z+IAoh5Dil6uHhgE/
a9cmPuP6NBX82hMOdiV2+oXSi/p6y0wZtdvkudZAhH0Xg5EJU2GCG3PeB7mvMG4O
4v+Il4eHu1CnflNJmdQrrY2EwuXdC3EbdLdaa5TaaNIUUHuAgFnnT4PN6hUGFtNu
jXvF84K+R3KCZ3ez8GY2yEoisJj0OY0LOuACEhtcHXylhtUSKc6fd1G6sB5acLKh
j5S4BZgjzK/I9ECyJRTRE1MmKlcQ4PL7166mPGioLO9+IRUq7VtPzyb1dfjKBIwq
sdDMftihqHvobNyhpnff9b+MN5CoabmKa4+SAveo8VFwm+o9TjXE9y9/JUuY02l8
qZYxI4OSgvW8s3YK/e5+W6ds6B3YiA9cD+kzRIT16x0IX3i70rie8kGvmpYidNL7
GLGKXMYBtQuK/vm2nMUeyzp8b3j92paF04aGSrlEJl1fFAtoTH/RwXu2ajc1gfY9
T6RUTd/Hte4sGXNeyvAryFjj4mIzNpfTDimnOdTMNjh7Owril6z65EI7r7MHdNPu
lFbitroCf6H+5ghBi7/f14NpbzZcI71AdsTv+/qEOyT7lJtW3lvLZ2XBvSh9ATMi
/TjX7SMC6uF/+ct0LueDlEiA52ppk44Ot222uuhkDb0tb0qh6IKgaJkj5AR4QMHP
0IzULvBBb/BFOMseDiFablxN0PQ2ugjE/Xew3/IotegGpdfZPGPYnyCunsbS0eV9
0F6OMWgM6KC2iS8aa7OpvwzQGdqmUEjRnqwULqAxrmzJWpBJwUJotEY+aJFtnsjY
nLYi4J72Os0If4gA0wp2+ESxJd5s1fjbZXj2Hzw2py1ehxfto5rFuq//wYawt65H
ocUY5r5KKmiuY3+XbPHXVeyVXX5olthD+K67cov97zqvGsuUPEgYpR7HU/lfstxy
B7yQO2aVA7ysVhK23KHXxF3zlc6XxBd519sIb5gzkOy01KBit2+CkFivM5JVB8+g
lAzJOsZOd+baGOG3mTACDez/gBx2qL27JiH9Tn45ms6GJyWKpzQBvp4Uooxuoygt
dtIcQf9z7TDlQog6i54ewM8Qw3WNQTc098LdFz02fydxwpodirt9krmvL32WOi3g
LnC7H/CEpKxCMvTatKmN7mXrj8c5E4hzBLzJZEXwe8NnK9N84mS2haQRF4oybPNm
asw9WmqMf7aAe6u2EHQ/xwNKy6ip3DfVbeqYcse40F1a1xnHvdCb5iLudvBlaDmW
5XifTPsNR2aoJtRCNTP2+eE5ruu+Ap5IlLq8LPLnKBovE+lSgU+MNGgAe2yshOuA
5uyaOFgetvYw+Mbetqo3v8GCQuHZ8sY4CtB/yytsd7C29AYq8fzWYzCDI18I0AvI
aHXn67NBFS1kwwLj8Bsix0YjkELpyekrN1GILE4BQtlVYEc8hdGjZx2LQRHcSmJN
YJcyNs+VSn+ZArwbmMg6wB/wi800PAnhMow9/PpOJ6qP/MQDn6BnQ5GMQawB/1NV
nZstH2jh4fZGf2weJB81Lw==
`protect END_PROTECTED

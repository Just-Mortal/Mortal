`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQviGnAq2UKsWXSHuR86BjXyKuQa87j2FFWQwZkBXEZwhJ+wZvaLMOl4xvPWboD7
8Tn/pgRyZ+2NIfTnEUgMybGuzLKgeQuQ6lsEL2yMYMrBQGL7UIVMA6cabQzhQtTh
fmRszyuUJo5oAiTOy79TldE3+LZkLzmyo+h4cAs0tB3lGQZ70Eq7ruMIrCj8jq0U
BxQY7OjxRMAIOXZRXUWAmrf0frX8d5dyX1emBzy+s3eHvF6SCx3jmSr8xV11n33V
S+RMfe2/d70+kG/xNmQwoDpeoTAfTtwy5k9asERDyzXjiZdbA7yY8wEZEUa6z4hi
F0fSV/V278lZxjxuwVpb0P8iAMswKwTREtVFDSZzMTbFi+mfF+FTwyL6rJKKanQv
41oXibwC04b4eqAZ4KqfYKyG2eAqha1xZTZjPY3pnXwk3CTXk6JFdfmKOnMM8tm6
SkEliQlyfleESxkjFZuSAoLv89BRk4IWxlKVrLCIxr0vR/7JTo7RwVpHMkAupztQ
SrKCeLsx3C9Tti1KrS96MQwubWneoqNVYbJ0Bzwi9eKPrIya/zkGGtZr88kvBOGp
P9fst664gd8f2iDSWEbSn/5l+gh0DA5wQe9AibE9Oh5L/LClNNFcy3mnfmUFAm9r
rq4bpvsvOpApfMZpD+v1oSoM0RB2MNRXZW12vk2ObOMH92c/t1DubU2XfYpe8Aqg
4v0XYCbbA6p/zqRB0QPvg8cWPw0LK3eNrbT/lBoxYGytILF9xDI1j4xU2Q66UDcb
0BNFEQsB3SUkRquW6s3irKXazsSg6TPyg23OOceDZczKshYNKsIF7MWssWQbEFoG
lpXSkYpJVR/nD7OTJOkDdMgSadv+fdbT8Ig04e8+lBcGfrs3C6tZkVA8uJHAwcmX
v0MGcBbqRLFfwkjCLhLbi6oNWovI4TzIpHc3eoSoTqlQ8AdmDjT+/x97xooYLEHK
0I+iy0VS1tGmH6lGOn3roM3OQljWQs5pL3AX2J9+/6g4FKUgBsG5+xNYOX1BZS1P
1V0cg7ViO3DBJ6dFGzNXn0jr1MZGeu61nXtc3HhctGq7iLWJZd1JWo0yLKp2hb9K
j0LtLD0Suc1ayle8A/hUrnTqWsJwjvNGNx0frt/myXO5an6VPUQ0EnaOJpkos04Q
XR3ic/7TRY5VP/aK3aziUXL5WR6UzTC+Xed6aUqKL5XFQlSr037ljb/NHNjey9nL
d/8LGfKeAobNP2PSraa6nH5Q8LuMzlUZ6QVM+9+D32wYKxYYPTEOoQpxUmFwMGrV
zOrbpE4YAmhhUrwNSkWNQIQwGSpYdK3P6bZNhr+t18CUhyEDCThFgUgiqwMYoFCX
Ro38G5BBautshbrfZQBp50IIHDxKSpBOWC6a/MgLrkrh5ss6E7s2BX7CMrl9w7PG
xPBJHdEFDlejNjf+/5uD8/JMONlpbOivEg/uS27ssGHq8I1mCxVTEuJQak4MThUF
eyu8AwJ5rX77wkXUhlreThgDIaaKPytFdGOmGxEPiVJixQy/Vsy11nHirKZkGwCB
MOF/ivuaYAcTosuMv+JYwKUv5j1hq2hOVv3ljJLD49tSF+kru9wbvzL5FqPMNUY2
o1RYtjjjiSB2eL6Ha/XaGzhQOcRAUbyZFOfcqck70N3y4RL6ISNJ33VpW8gRr+8q
O3uZuq0wT6mvPmanBFwFgyB+ux3rKhm6dGq++U9CNoK/Pg/Yk07ZlGBpPvrCTCek
yC3myT8hWC5fOY0OqBf+atWPrPvZFfGqv4Rb0O2UM99y8546wlOFppO88iUF4/ct
qDeXPLGa6ny5wRIfOHdOC/RaBNm2slMRgzu/lpa6CLSylz0/pdY35uJuvLg6QXDj
oagpdwz7e6Jp4mMWSnzhtcpx7IqZ6tkyClZIztQkbHVd7cxtDdqePRuOk5JqRTfj
XEERrjVJ8IxGinJA32G51AETdYVF0laHwCh6wE/ty5lmwXr3SWO/pcoUt/8V9YlC
mhCglFLnjLlwEqfs/rU41Um4nwNhky+rC8qTaVsHfKqNQtkcTLLuNsD/6z0bHBIU
uUkIYAwwrfMjAWC/AlHKVh/6Xyzpulapmq51YTlkc1goSq1PHlsTVl+fnh3bIGvP
CsEPTXj5nsgLJQp8J1ed6nVRiyrjziWmE08GP6uaEdZ8t2N99Qgu0UPhdQzbjjQM
WWSg/OPPdZCX2ip8zrdrKB2AJvO73LYHmNMPF4hUKb99hvxGPg0VGIKn/KXIP7Uy
6hfXqozhM4o5RkA4krHShfQt+ym6dwMgbTsfY17VUnhv1dPjwacG3NuL75MUzeAr
2fTTfPLNPIfaBKvaHZZ6n72K9n8CqpTiF+nkWWOSwa0MBn4l8H/YBmK0sbQQDbTJ
8UonBUH9QiuVGykp4lPemH49yGdpUa/gTVBcabWqGYceoDkF3bBYJqZ1IANBfoac
JmaSqBSahJ+XBvvhgiqGEdskxF/wBT5aBRVKB8O1SAzuvi+IrkaJrElVxTaEfDwS
pIHO1Bz+qkQLqgtbz8pRb41wUakYlpbEotcUaGvPu6xmddCJbD7UsfU7RYsMfb9u
vHN4E38Y63O9RqsltzBCRvX4ijx4kEWVG7/aVotTx72gmUwXxo3Ufu69waATI3sV
rZ2aoTKh0L/I5b9XtvLnFA0rQVNAgw93EdiBeyuWUm2Z0or92AL2/x+SGLIsKgFI
PU/BrLxdqMjLrZS7+KLQizlwHKdjojrsZOEBvm8QJ4hvB/wwYFVVsOk0uZ+/gbKe
oGdCdBEQHb7j/f94sVNvnBXU5ARU3IiRCxIAQp+EX3UHT8IYD1R7luIOkhwTkeBw
1f2+xGemggqhUgOs57pKRnige4LQb8B56jwRq6Ju1DsqxuZp1PqLMsmxqCaEdVdQ
YZTvourMJSv5uO1DK3PRfMax6c9JJZvLUHk7bbhOpmopolHaYhj7GSBLD5igTEP2
4J8Arq3X7Ultrl86MPqKxRGAKiW4o0kiJv5MJTnx26T0AAr1esI+1baa3YR4C/rM
IHtVUpthRJLmir7j/Tdyf6s9LAAN4RQj2kSG1JaaAdUwMJ49X97Muzzf2CRVZS6T
+7WIs528AMcThTJrR+/8t8NH/ztoJDD8HsxHHWRHAqUy1qBCwwjIClXhLeS4xTXl
OI3wBJbVEhXyJtF6K+wgKvQHL4PKmGMcryrFEbGx7xEE9Av1d9i3gCSFHDL07yno
KLClldWdMmgfVMitxSfrvUlaa8JW3mkHfg2FDVjuY/tDHr4p/uOJpBwXHU5mRfkU
vALxJ/XcTrZlfGgyElhsVycA5Xu15WPvd75zVU7oqlEFYNSOQMq5C/X4VGd6zzrj
N0wXNGJH+Sqm6nkXF99D0PWZffIFnc7pzHwUS1uOfdVmw0RAsspKglxRt1k+0eR8
Q8nvSVVzWbnr366GbNKT3jlfhTMpEnPqUcM3N3aX07YDmcS/3ekoRtaUFJVtbT5q
/xBePRhMgY2DOtNlN9S12kedAZPKNWURRjggOUgqI1awtGoPrNfbEyiuu6c+Y4is
CmAKEyqokszgUvD6W9IGOYsXt1AnA+f8bGL1kNkJI+AJ3w0V+OZGdpeI9JnSjLRQ
iFDFtoTRkk/RfQPvSTqtvSMZMAvxTJr8BidAm70hJMZAVpIyurHBOgC8j1bQyyMF
zsnE7yEQFHHHDPmllpH3MHT9U7gsNQACq5vNbA31LsRCLY9Up0FG2Vx+zwhmLauM
t21OQfS3kOpUOREIekd8JeemI1xnSdPkLXYDc4D+QZKiuDQzvKtiWRX9AZpWMAgi
nZswPJP+/L8jxDBz872roekUQLgqF6onl1c7CuIDWSbeah7w+zFIGVcxF5lA+2FL
CX1tkuhWGGEZpPpBZ5JIvU4gCHluKmBl4QyqVWYaMcY9gN1krtODl/zbifzr3bBc
3AL/42KQEb8jtajHkJUCs5l+t3bIOetkyMIMI/GvlrztW1Kml53ReGRlDQGYQGNY
Hir6vxfwIbYSbsjtjZ8USDgIWiZMXZQ0eOlVgTtvBWxoIMnDAcaPqPvhdVjMZE+a
sOqY2dmls4F1k8934El0k1rof+fKMW51j4vcHd/nSsEH/meHWzk1cRmd5b6lIoSO
6Ci4x5Z71aoJ3KL2+n9PrhosgtImbCOp7sWf8y33h4fBjngsfTSjt6fTxL3ZTVMr
HIQYtzgz8Tp3y+16K4wa59CsCd7H7+0GeRPNeEycgGPLaZFh8AP1IlBovla/MAvT
Pl4gMge9PCJNXr79zyAOwCQEPydXa8qvvHPMOcHBd1WjW/bFW+RRjgJEdvXwD0RA
MB3KEBJGdsGx+1zmhoFi3sknmcVau+PLLVpJ+kP05oN6gNFq0oqz2jaTWuNwd6EJ
IbmMQ2E9/pvwF4nM8lOCy16Y8b7xCmlG8I15N7h9MV1XQBPPUgBqDmx9RWarILAz
pJYu2Us3F0XeUoaB8eC1GKp1T8kAlX12cKZiywZX0jmHEkUy8g3TaC008LaEDzxo
x6BU3S4+rvwxq/DNNcv0ZkDkR0HUGhYlgy/S7y583Lq/uO6hJCY8yHwZhcKkubaf
GaHoc8fUNTOhOb3b3mLH0B9424e9urmomddddF/W0jObAzLtga1YPF56EwplbDPY
gjvc2a3xAJQQJBd7yzh3uvxKOoYIgN2SDygZWsJFmBaPdZSKZr5miSDF4doUZJNh
QpeUC4CGw9KfE06XT2UZH0bEZ6yW/R5lJaUUfsW4ITFofkQyu7gy6uqUazlUJrcP
5MKyl9UeOUwqYG9ng2UWyVBeDdhFD3faQ4bSak25vZ6VlDhAx0DIAKahg1eyAU6e
6gxdaE1Jt6eQgAtVQmewaHqwJPkNq6OvuPbYtnCXSctDJqElcfrnOWCM5VRf58in
WwGx3lyq69fyZd4Yq2xdFLqSzoo7yRV4np4X6t1rFRbpoTu191CD7siLfXX2zGUc
+hYoJkx7jMybFOp7HPryTgkv5j4JVT9q4WarUQf5PA/mtthuPK7gPDme8jFEJvFA
ZkEYbA6kksHlGC0yjE4iVjGxScsIYUiU6QTvrte8qtALcZB1W8v7s9OI9it7GNgQ
O48ItJG/NvhGx18sgWV4UNrC/lKJReOE9LuH9EC1cUTWF6NaLqLmi9YaEmfrI196
GhX7smLZv/tM7BkS5XFWWq1cm9MsPvI6ebbD93Vi1gJgk3dKOdeMSjkCv9yU8WyD
I4f7eixTn4CFZISLx3IQ29RnHuCdjk6rhLJ0v1KClE2ie7V3y0hbLajVaW9Pk0kw
VEjFAJ0GPWXGhoaDjcql1ZMQW5Za8syXPDTPyIBgSKGGwSfz29lqwte67sOWYswa
TTLQ/9F1TolI64eyO/BUdrqH/v5zOqKd05YPZELVTNpgDZzgyWJBodIWWsvshLUn
W/9NmF7U+5DcvK0PnwGPm2f0c6CPk1DXC0teBNDv4LfT0xu9w68GCAV6ZR60Ga/B
v+Sk8e8T8mbVFCfo8nPzDpRBPFZLyQjJDzeHFMRSGGddlnmHgZ5vL/3GCvx1KAp/
amcPNHpoCUi0zXf/TEJ6Bn2qn/8NMDFIt9s2QdOLYSv6tj3LVVOmsCCoZULsDvTL
6CeIF2ujLoCUVI9aCA8AWznO3mS2ku53eD5gd4w8oBgHkCGGFSLrNyVr28cqUieK
+Wu94tWSxJUqOXGzR44/NlNmsEBrcBqgxHAxAvl07EXjo70JhPl4uvqJXdTnr6kf
hH/MRMukHOWVFOIEpiZGDTvXCHlYED3/p9i5li3loqXqX01TQb2Th+f0NS1UIuDr
Sb9/Vy7iR/b4oRpUz+NlFLieodZ8B2jlFRvnSCEqbVCU5oxJOL2nHR5IUbU6Wmg0
Iu/gw2RYFUdJfOeZXzpd7bsKJXK82UJgrZXGjAhMlwoSEQS2BN8zuaX6Rch/IcS7
7KJGk2n6bEksanx253dH/7cUASTGAYH+G8EqP4TtujcZZytD47JsTKSUX1EocAbH
MwzIEB7ascpto92JbFuqqpWh1VPqzPzIsS44oxp2rUe5IWTnHcaWjZ/VX84iomDI
IIuuk52ZSzRtnoP/oFz2U3e33u2IvfSHUtf54rtmL9C+N5zOzMHSSg3PSobN8++a
tO7V9bguqr65yeGAGizLAqE8yslZt/QzqkG+5CLMxXxWIorVvMtGKyzkRQwGqBgd
jfVrp0sdvga06fijqpDaCLNcXme9KTu4UHSpuMxwwZAVW+AVUAqRyw4Jc26Hzgrq
ZD0l0rV47MvcM1PRdKhZ6XASPzkrSYWukehmCdEUeZ8mH3CdCT68SRTydnJWpmCD
XudS4VuLwKZ4YtlyMsn7yh/BJFIxljwsdW0UFpZ614pGBXdfjIizbDdv76TkLE54
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uq5pt5qMQjK0MHB58jXl5fEkqgU+el0lVvfJv+0BPCZyP1UYGb07oGLZF1K6OW3N
gYfEvkwZ9djqqt5JXa8eUPC4HSwgRmErfKkVgXS0IpjN5tQlfShdhwkd3W6Q6UCk
l3MoDrTO3GxcXjY5KW70y7E31qs+YIs/YYfzyCkwseVXC82+vgl+WdMSWLgWkYKU
n2WPleWsBzWoLkeUyzFnj7S/0ijz3toRNaVnHk2gl6jmCYez3J8Z2FFa6jzS096T
U71xcmrQ32ZKVJwpsBUHmBO/pFTTP6etbxkfG/xpA3QlsQ46Q/Q5Itdx4Yxx8vSc
jXXcwuHFuFXAG/O2O4fxecRAoHQpF520+yL3ZQc0UKnmYrCscOzCyoqNR1qV6RaU
IvcDvaGOOxmElXbP+hXz74EjKIn3mWLozUSKo0ekJvVRBjeqRElz0D4aIAkF70MO
Qv2U45BRSikOtgEilBGMtPHjB4pNoi0U7QjLpNlha0neJFdI8NnubDyv5jyl/rSm
OslNvH71YRRMJh3W/RZ2DPtUttCSzobj2ZaJPVhbIWxpu9ODk2NLC/gjPRma6XCO
MM0zPlqGLA5ipIo1HwS1NSLPWLOvBfqcIhuoeI04NG4J4XJGly68BxLvlmYLj5tz
9lFJg09rqJk5htAk5t+DLpCSRC1cXoMa4wHw/p22ls/sU1zBYHApnUkircKdiPrO
r+Rz74ZzBap1wvNXopMIOgMCMxJJ2zE2d0afX+fYe6xKcsQHBBQuuM71hFUZ+Ep1
a1/2+u20ijJd1cyvRWkxA4r4p0fD2AZkuLCEWr+0VrcbZl67hR+Pv0I6zyOy3+9F
eBF7DkFV+/isJglUfaRVZw==
`protect END_PROTECTED

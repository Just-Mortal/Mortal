`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7llKvEdkswEZmmupuKWjrYeP04DTxE2qysZdWNxugsaobnBo9VONzHO0xupO+vH+
Xn1pzQAZcJqYAldGVPzfkOmF5ekAjMwrY3s6Hv9NcADBtvxy6QV6HZoshMmjq9ab
Qgw8P/QfYECbjzgp1vgg62hngu59o45b5Eg3Yd0OOWQ2hfUZEViPBy0ACBUuH08q
UDblvYB87Z46GsUC4Rf++sZK7Q0zEuGV0PLNbaYeSSFElfBHZdaT7dv2/fPhZVym
7WnS3ooC9YTejiuqbp+3P8aWLVSI5h0AXi18QfTxEpXA+zO1hCQEyc+DZV+LmuWV
+E248vQ9cMYkabdlRiLYRuRZ7++Jc1rIo+Q2jSromU8CaP7L6uN8R6INchmIz2RQ
G+p0BHtdJ0ZP1p9dIqvm6oPW6bTv2l0Rbz7AtOxp42WvbebRemFO5FS7rEYG1Ple
QyB4rHSujn06YnNZxhHZt/xGe5pvKTWT1hfnU/uRcElXKeHRRXqIIxzTJXKRga89
352bioBm8Zyej1V7yeN6cX73EN49sRJmx64XvJUdcMdtSwzbYu0ne/Et49AabfDR
1FDEqz9EhnKAlfL2/TalYT/XSsOS+wQo528MLqugUlWxeQf/rLWib7oU4I63fQqE
Ad+LPBJYwzQjYY/nZ5JCGhdVKRyrBq+GLBprLxkUobO3J9KgchDfzfJjg9UkJ1Qm
fS4KP+eYLptPWdZFMYxCnfrqTxZ2YAZ6KpCDsMZdWGncyyex9hbItmnttAQIbM6C
+wx7rAyHX4lQtsbx7Fu8DyucvQ8NMedsDiR+zPTPj2Y7DWrxNEOSxeC2TDVyVMRb
cWH2y5h/o6HpYh/EaEqdwYRO2Ly6vrkBJ+XxWjp+te2ywVWuaJaEUIV+XO8c8cM+
dc7v+2L5Pkkzn59FvjB9ZQWsTVTzgaw1J33zNSdQOoOq8Y6T7MMFBC7RiI3siuVR
TLzksd5XVm45un8a/7xkD0NI67JeFtqBT42gbuse2Xa/586OCzJbpF4y9e2zOyC8
wRkh2DImsuqmGodxp+kdklEnPzknDhzqFWK8dIOVf2Er5YjqdsClZt5mur4R1iR5
V/xoDZWWPXXL4WPJFt0ew000LSFZS7gIniVOlk0k02j4iyOEYHGH8Yd5raLp+c95
wZoSgePe3mRw4EMAX7cmFshqAiwnLqiwJFqrifxOcXURH18ilIDiBEJ8kD76R4/4
wQyNmHbLU9Tyx7GlwB2Jks5aUL0Y6wzFwNHGVbMnWbFAFTHu+68bhUENT+7hpbPS
H2oxuKTFMGpEMSF/0YGhd5tPXuprJP/NDlh7gp4TweA0nGx//krYQjhSHJwt13dV
dIR4bz5Ej61DwYDQPy2GyInswfbW1BFycuI7iiFXXMHZTCaCu0cTbJoD/cYrpTAj
qnO7cupnQecMqWMW9rUKrZxNbp+GvCRYA2XDcDkpHm/FgdKnj4MPCN+v/d8OeuJi
V33nH7hPv656yH2FNvxbJ4E/NVCN3tscn0pkVfR1X0gaJRApobz2l7TAjgCDzyCs
R/zXiQ5tW+aKjlwx+3i+AJYWdiObZ6mvPd3BSYCUbBwO1HQIbLULMtNTXMlIU6oT
XYdqxXyZ+tABANBaB1iRlaIViHGWt2cbN24npe66Qn0k/0bvPdXehaOZdK2zrAtg
AkzB3TZTt9AMLzBqgyNvNtRyCN+eAaLqoBN32BscVTiDLCJdcUGTuYbKIfeD+3/W
zL1PfBcojBulA0JWer0zseRjxhfJTYi4eV91DjQnP7HbOKok6lzgJ7Caz9VAODOt
6ONXWR/fNxy1WFQWlmraDv3Mnz+qCLhM1bury8y9AU+RnDoJ6vScOJPrJk0ulkQf
VL2WDh+Q5vYO1vNnWgzGQTvXQtCyto6DQeR5Sfxvmz5kAZ9DltQvCbnq2D7CVaRt
6dmm6E9NPF6IuD4yOlRuKSqhf0LIdLROE+6xgc2uvTWo72RV38AYzuQ113QclOWF
h7kmBcdV7Tjnz9k1+rIXDne4rFn7X6GldRvLjmRO5NuG3RyJbN3GSwCefU7yF/kC
YLfqdWRGZBR+Q7bmHQGtfY6Barno1StyIoH7QxQxpBdKdlerWfqAMVoWKp2cacY6
7k/Sehwcav6s3pxJSuOEvoWXy5PlwUQwSc6FyyAUZtZhpCTNqSgE+AMk9QdRbGN4
hpBzrFcYmCj+K/dDHiW2Df+ULyj9JfIAPm3W5VYzSEk/Zuy+d88psWOqRwp5sdFg
QVCngwwjIIW0UAMFL3Y8tJpREd8ddr+lFnQ8vDzl4hI7AJ3ckIR/eJyDa3dXb7Gv
lZgNESfCsoWmJ9wKrAH7+Gqlkrd7j+vQDZZSsxXAuyfplPZhd48ZQW1LT/z7X3bf
+QRt2vkQOorBpNDXdK566IuZ3DD/oje8rVSPnBnPVGlI5hpW3JVyAj1Ayz0/FhLf
kb11nQcv++FvFU2hMy3GoqjehdQWdUBVFKX7toQwVi8sjZXEK7BEb5jXH0Ivsmik
wmfBnB0vWCgqN8RXpxOWbaC+fIu/kx+d+ZnHR2sckQ+Acb7C5Ebl4KcQzWXvYCBj
FLhHTELDls8sI7ulCDjtziR+sWoO7XoD/JpBZlLBtansXnBiUR0zHtUPUiftqWJZ
6QpsNuJRqwtWCXPWvZaqu2quEiJ3T1fRE7dOQcFdXgZrUwGa3k0RnVsh8kNfweAa
LLphE6Xaf3e0g5kF0v1hj4VKi+6ZmNDLAKdvpN6JehUTPPXM0Elb2G7FeGxxhi/2
ryQfu3sZ02RmjiQ+7weezemjQQpF3fnEqqocMhahRp3e1emfJ8BjX2jKMULe/h0u
ey7AZGpiXi+svH3+KtdWwBJBNhOlYMVWcVIjKX5RrqRBN+6/joY1nB/DfAyc7heP
1muD45zA10oF9SIlJbcjTvbxd20uMkvSc6c8EfxgtPfvqjTPZT/EtYuyJXZlEu9A
B/fEnOi28F4wN/Xa4Bu2kCKUTygQZXJu+SLyymN0AIR3ImuxxFOfjGZ0sHrTFjPh
NMDjhjOYCkZLYi1BEZHQkOqYg3NqADylXotImLaTWQD831SL6zhn991pu6CePGWb
RpxhAMM7mhWHEK2SyC+pgaualv0UshzOWKyjIK0OTcyvlW3JM7aM4klTAiAVxh4a
Dh7oHw44WRNg1+9J3PM4N0i0aneKrdA94DpKz7fKokiIzBib3kK8tJocaTNKJqGh
kpgkaRpec9vbcDDBjeu/HUXZ3LBkwoLJbkXAJdvLOMchnQmL4ulY86QPZ9ecQqlO
2lxPOFQ3tnCG3kGeoXrc5hoaRDHA+h6gKXLhJbqg9hb2vcx+4W6QZMV8X7t4/YpB
u0UqdLKKzwIWpihs1poUkPEbNonoK2p+K39Rmuuj008bKU92gUA0trEvDzLFVNCs
GDHY4qKNAiYpXX4dd4iaAffEdlUxZ/r/kxjxvJnZ4UU/a21CQtlVbsv9do2h6h3g
jE5vVO9awndrWDbh3SP/iw4RF/QeIp3PXyjbjoS7nLgq64xCA/JtKSAKMsT89KGZ
+pG5VisE/6pVTzP/TBDDZCxVfJbjRlszPOadac5gd6uVaRb9sWUndZ4+tFm8g343
npL3HhXSyHInpeZNNMX5+BTsXwpgEbTK17Q9cH9kQ42Jr1fVL3/MlfFxNQzrHjjI
72sFLQxoCaUjIqr2SOeFNT9ojSlF9hy1WMF/FhynfferxBLFQxIYrH/d45oV7eG8
vpFnjXVdOt4fFD5fSuCzDTNqmj+wI5HPeNvgCwUNTg4nau1oKESqzZwOKV0wmewE
GCAgQ7cJ7/rJwxOWof5dQRYKst2Migy9sS+facWDJJ5j9SPhXJLE68a9cmT39THK
RIWeaaNNTNSBNd6CXGK47g2nXpdAFF76zJXWOa6HlhBTMUZOY/N1OuUEYysVafLE
q+E4XOiZxC++Oy8Cq7y9lF7LTI5nKhhtX2W+1RiYHelylkImCnEIGcEBsTcmfJHs
a9QUU5gMVhEvfPtsKDifCWa+oIzFUG4N29ItnAiSVW2bZfUi83EtEWPnI1tEJnT2
v/1RQVGiJ4YJ9TM4iROqoujkhCEasd8PAIF10hrJlJKfF2zpXWD6hTSOgaza3yXH
KKrKCu5cRNVJRWMx8NtgNIdtwzpPinBqoO29cDR+k7fOB+bjwn30Fu9+Hme+EKZF
QCH0mMaFgFIIr7LH3ObF+nT2leTsr7vNkcRBfhg2/elyKYfVIYBoHYaqUUbZAGn8
vIRP2MY1BdeHEG0g3/tepm1cW7FG275a3zF+8cg68z9yWABBhHBGt800jzJqUURV
dGd9BOn/A0vFibDr2+zX3VvXYe9SskxeTmbEgxoOaabUmixGd72TEk+HhxYDQdWQ
32XKwPqrcqrpNy7LNrPySNdYXGsLmD+1OWLN68J5hgWTqWSLB7dLmSisuRgjgsAb
ewZzfv8PBOTp1DoVc0wkfTeYEYMOugfKoR6Ulen7z7Ra1yrJyiNG0dS+93pzil7q
eNK6WYwZ7nXKFqXbQR3L95xEQA/X0xKHVcdQIMfdEFMqrH020bNMrzPd6Lrzo79F
lZ/69RjeiOl1PLCGKNwN7vIk5arwirLWj1YOUBZ+lArQVGzqbwNFVqbH4H0+fS9q
aofB8KG7hbmakOt6e32qaag5RA6nV4rw371bLpPYe6PK0NRPE1Dpde0pVIT1rStF
t2m7KK3fWt6GlPUVb3Z/w6sRNfbmmUlj40mLdhu1jcKHphgbkfVUl8NFS0a/OmXr
QplSDBBVujv4KvPfyGzWkS3iyRYUw/mXhKtp/3cyxtcep8g4uBDDotwPtydoslWw
UbAG42wSQDyOBot4DZ6nTztsROWxtHeg3bmRqYHK3fErj4jIE+jEm/ydrjvFP6B+
pEU8DLIFy3imGblH5wQh8WCTCKos8ni7nh9LyUb7xNK2Xx4rlq/1DXzDqmjEvc9f
d2wkOKYniOAW4BAqRPv0j43opjbNVexJrY4sRamifAyYI7NPu78mtSvshv5Uen5d
dOEnt5DpPFl9Ekv2VvT5SQeU5y5SCeMxoGZo7FADugScwiDMDZGsi+3u7TufYd+e
6ukAcnS10qwZpXcQGufitxNJF0dpXbiXnyt1KwFL9htoqVtYPBn5S5jggJ+Tzi3/
j3yNN+TdiqBMUTbb6lXbP6QMTxUkY1qko6M2Uyfe4PVZoRJFCNcpj0e3YYU36LAe
600ZkpGkJYDY5sOXYEChv6dKPfL423DH6fMTD01Mr5SM5p1hK8ozi3cpgaNJxvnk
k9/Nq2s9mLYwL33tK4M0CUMaCmSdfe9YUr1HDxUw878o8gSutePE+NDkSypbq0EN
uAKtx066lb8CtdLxiNNhgRRJm1OPCNBeB14+nVvK8olMph++h1DYzJHmmnsUYa4S
sktTH/qzaVSo3rOfaYAK6yEyqdHMj7W7gF6KlqieusYpP4SpXOcCcMkJl30My4b6
V3aW0C59jlCzUUmtC8qK8nF3gc89AgzfPlK9668ek4vCd8v5VkplWYPLlkdFZH/h
aBr5OVAhU8k9to4u1TP9ethmvfrJeAxvhDUt/6uo2kBkclSFxI7+sWpBONetrino
qTccB+5BxRJokkNAKEo7eRQNfQELr74eMfyIFONJUjuKrFDJ33x+ULAT0K1Juj/O
Hq65V81S1Zg5826xg/zMb00eyLikJl6ciE+wPNqSI6Etb1mzcboAQS/RqENBkKTB
sKwGI4u0WdGe7xuhEjvrj6il2TeA5DurVhI9+TLcvRzEd5d3bg9S8g4kbosr9/6D
C/V0n9dQrbH09Oz+4KO6JRBEXMC28qOtGvFkGmFl7LRQxdgOpB/rh3pA/xI9iZxo
Ua8kBtqxJa362ZF3Fkh6IcUpxJPATUVODfNeLMWh+Nxmr/WcdmbbneTn5Tz313z6
Jz7+EcMtaEMtjc32p28NdRkVwK6GPhi21KCRyVI/zhyaXiGJYBb0Q1LeErrwYMo1
nsabNI00c9MVumF/pV1G001CWLQYu9UnsRd7ugKvHa0raIbT7dkn6mmCXjNVIbFH
/Af8p1SfnTNs6NjdDNgDGztrZfRunOTC56iJSyRg8hUtAjGWQo7JZE7vxW+wKt9s
wg2k4hthR+tzkSSiV3cofiSUfwSv8pP7nTRE3g4pFwAzAe4SCyuCCwX3dceap0Xb
/8fph+4p/CQ6boIfEBnFGtkTIDVwtX5UDtqXZLig/AhNDzNBgzOdDa8wBjmvrEWi
sV7OrR06X5SmK0uR+l5QUZfG4w227MRw56FoUWsusd5yYp+kiK8d63s+MVGnNwF/
UF14EqLyvmzB8zQeuTEgHen/xzUwK8yuNU2dyxhq8Qss7/3NruCu6I6B806x0Qce
mjtzTgMViTo6xrcWbas7AMNFTnbVCA49gJ0e/YWfyDICzAGIb7TztKeHt+isV9M7
laQJ7RzcbPRgZZjThk+95V7shgWzK4STf0mEYLcjOAaOzAcUYZ9IWKXfZi8EhIX0
LLUicMXbJ4kObEqLmed9VPbkauftkj1H4VhS+87AiK1HbIBQzcBsetlJmnZjUNqg
rkAM98y8h39vXMaHM+l7Ks++/o7qFA0Szh3hhyfPwoM/BeRH1/V+ru9iKusfQ5W7
I6YnQKlZ9Y/cTqj11pu/1w+R1BL9G3ylf5t2P9wTNIkhkf4hteseBEckRZlnUUIE
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iw6xjojN/zhgoo449rDPkKs0eGz2j4IbQx0BJFd3ezvI007I4a91MNfnHXznORSx
xbLqEP3S/WxKYcqJGkfeU1CDPAHDq1t+9MN3rF/d2gmYkzsRo8f3gMLVcnHYe5NG
2G8uG6dptN3pS1J0AXFc+PJQUSVxZqmTIBGR6WE29wDMZjDOa1dQAxZ/1JgsgAHI
qPSKNvFLywk2qtXP6B/Zl16CmW1yKMNyreSvO5FaekQJd3mdDCcoe2mlL/ADCjcy
rV8r/6C+S/txsd/MxIC9XZizSBswE20ee03Z2q6+TAOvO3iMSkj2ljiFdUlhhuY8
30pUzUJbWDi8KeS7N/x6bPbQ7xLkqiPAIKbL0diWV9GG4mQRtNUHh9OzXWnuaP5M
repmRXqZdq31IoKxUR0g8bDeypq5FYYKGy+QqZnebIM+NIGxazRYrL7BMb2zUSQH
33XWoWRrkyfyjsREwR9NlnoOjMCwtiju3/q+B+polA2thPOFF1eEfL4eu5xsPko2
3JQn/77gyUbVL6KhT+dCyNzVB2rNmJEg0jCNJXkMuj4SuhnuDRY+kns62AUPn55F
xNv/QEbj5P7U5OsZv2jro9vrjmXQsvKCb6/FZUX/gWXQHYKfJk4HHbSBvKTz0RpU
GLtVe+vxjV434trFXw5cLskoM8IAH7Lp/1yelClNzR1zAB7xRoI+aZualLDEFdLE
eE/ViJw3QEYlIJJvNUyncLCRTWAtNaTxiKkpthGcQXkMQyXFX1dbChqYt5pZpKrT
2BtOUqwCN6AIiz0uZU/RVe7muXfWf2ibu1G6tJdk6RiMQJ5/BTg22WuV/smpk4on
MPEytSEsXEoaWCsZJT6f9sBkfmNi5ijm+sdIWZNjleYE7CEGRmFMDV0btNuPaOZb
YtQXIgSUX32NBu8vW4ZKmemqJkPuNgoLkeP6UesCAWTWp5/EzYUP82zle15NHbbs
/+2vQ8On0iBip2IslOGGrOdngaqDU0e2U/me9CL/tcgvptfFy0uPtUXCCGlFINRv
CVoSRt7UJYISAain7cr1BRIrU/N478brm0jtTb8f2XGvqQHK9r0P/dTZ0wEygnsb
`protect END_PROTECTED

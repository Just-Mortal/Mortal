`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZKIu2WCByP7wqyOdWNGzG/JshY7W9MhicI/SJCQXaD7jnXe7mNiYXpy1AAi1ZD4
UZRp1qlmqk64VvQEQEtAKv2KmE+MMLKzMBKHzY2tQRi9Cmi0sUxRSLreZ9m8DNS7
awZDluC5ipvcOGQbJFeXUI8/7ySgYMCuxR3UzAedK7jwmZGkhUz4hYBvbQ0RwZeh
T/0QyWzvIJaThSG7nT+lvzfwDP7jMEx3kfFDchpevPhjkBIlHMcvhDERjGsEN/IM
DlBIGhjQZEyMvLSQqE4JJBqWeShUk9niadlx/HSd/77RAL4DZelhCh6/UPVBYPCH
KcAHmXvExzhLDHOE68cDGm6IM+7+LQ9RCMh7ojddxXf2YDQ2nK2BCJ7vIk118fRc
MuFyS96s44leI+RFcM7E/6YRiF1X58OFqzEKIVQXDRd82P7VuH01/LxL5GTHNI27
CLHjjTXZOB05va0WhmDebs/vX+HMWyJcGao2hKI4zGGjdJIZXgVf7+fVrjKXLtWR
1Z7ogfzEQxo3oakOY1+3/39BIGSd6/EIs6b7zaYRypxEKF8TF4cRWfYJrIHCYZ9h
0VGVHzLODWU9pewa2W9CDm9Vz+54wb5nbM0/3F3vqPcsoy6tZ5tKtmWbKoDjVfYe
ISkq8kJZT7VPFtscrY8K9CNohfxpaElh7oYYUbMZUiS+ioaXLMNCwnNPwrhuLizW
sDprM78O+g93Gao5Dub4rB1qVaT0gdaZT/Tysp4Dddvk4BPX0Fym19X0Unj0wDgJ
iJWdQItOpToL2LbRwbOz+H5dV8P+Ei2jCgJHSuHJssJQ8mKh03y78/MsGgt0zgvo
uS5WnB8uzw3HJp3D+JZ2nKx4buvJsekkR/d+1dhyquuaZhgzYujfAx2cnWxkcHc7
edWj8Ps8h9x1SIUXv4aagqnmLrdH9nfvRsnxBVqjLR182q+j0v7KX0d9G7a2DF1Z
CUYG+mDt+eQUJhg2MTSM6cuH3TKC/4T0CDB1UUAe5cdagB7omgSKDKTkdEcLVk9m
NeX8TBnjZF4KnBFL/gKTQbviksFfeeZ4XLOHnbhiRjT/RO6SanWfBgnJIDxJvvSH
w4UEbgRwrbiChCZ+TbeH5runukQf6E0emdA3glDUJIM=
`protect END_PROTECTED

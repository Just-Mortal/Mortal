`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPQ8exbpCs2Hwe+qwbG06JEZ7RiMZpLoEF97G9YfqusZfNAiXxtSTv74vVRMpNKK
1PhYl0SgtgcwNu7iSfRPJ3PtqmwEHMArsrxA9ORuRTosz1nFuXC8Ed875/vCIlXM
xRKb436fpeQ3PgtRShoipoyRy2PM8fwFAyLYwpBamazCChFuXcnWehUXfaGUwY52
/LpT8uV1QEupnuQyU7XB3766aj8/VyRHd93hYMGNrqfkeV897qEsw/iaRIb5CPNr
q6O8mvgoqaC/jALUfXMZKFjRxg/HYYz/VkSfOE/GZqwx7FSa4xjcimhdEjdiiK/F
WwDo7tkEbWF4u+hU7u1qq8umLn7Hj8+G0eZ014iK7TowPQ4kScthKwU4xDaSCqof
BewjW9RdAKs6fISlXdWTYimSLCuXghxjT8nSUrNnc85HYXz51mQweD8MYMvmoL5i
0kL0DpEu9jczV7CE9oFH0WKCPMwR3V/qqO6xikCCtxs6LO6CxzxaMQVBvAy0N+SZ
xyBvbtZhcJJWR5NlxWFFT2X1Yv981bdXdLfvvh+uUK9icy+QGTPCTgB0uNa38Bsy
4X81K5ViuKdN4nQmcoS6nKmKbgMTaHOvrjAgHoaqC13eRmBz4JvbPP5DZrB2umDk
3WoFstzKTAuYrQFGQoROkxOwkI61pRLf5MXuiMqvpQpJI0v6vq1G8CM4aeAntOqR
SqiD/MpBf2Y4PbBNovHlKo5u1tD4d/bwoz42B6B2X+NmMtBK2gl6C6K3Gk1p5mj9
+QlBnDit6G1ethxbUiYs8xu1/CDMcKq2qhbBUeukn5lfENGQkHblnm/FZFDR0RX1
pNooXWC9R5YwLemK0HTVAm1zvk3wBP9Uou1mTA2qyPB14hDOjcQRjJsFdbMXmNc3
l+TjNbADMI04xrTHIkUQwVndQla8rPqMbz29GBZ9ngDxLH0WKC/MR5DR43fl8iYy
VKT+lTR30QrmF1XNYlWy0DMWqNUWIPp773/o013ICaPkaB2u4PZBOdi/0Vdp7Ssg
iLmIDxIWKg/a/995LYT+JC/NLoIPoD8RTq6wYLLHPlDsN+Rvpxqe4Zv6DlxeQsj5
KSLL6M1MRVOl/TCYJBrRbnw1cHoshScUKSZq3ya17t4vyUngAvP+DThkoq82SUjq
zh54+FeQJNAzorvsSnv5nHvzim48BeSWLh2nXA83lqWRIm9afeGXn8cwg5Z7paB0
8m+m0DnPQPBWX/IQmu+MQCQLvJUd5uFHGvMetswteL7U8iO0cJFyTk+PMi2BGhRo
Pn7Mve1jENs8B0+ieCbKlLqOsdXgnyIJGvq6/zi7eGTeHAA8Vi3gU1jSMi9FdgP+
jaZUVWSYw2rVtneSaDWFBBisDYSKsVxDhFDSUFg3bYN9mNZdSveXm6bsJjoz9g26
v848Cdru/EQxdLfNsNH4yYrJI0PWHXOU0f/f4zaIPIQg7HEdvFw9Ck7a+IGB0Pea
flyx30Z3P/HKeAAhQw6crOeRJsl0kdlKnGQj2O3Vn4kANEWRaMKbks5otGYANxhz
oVzlsgsdT4U8leaZ7j2DbvZzcAvNJMS6J7uzgu/t9lQ/SffEzCN191WKl+lGRyxy
RRoIn/l30EvdjEq3Miaas7ybq0u2FpRqByCWksg4n+R6pnNBzID/0xH8p8Udw5u9
w4mzAAVqTuaxDfIQ3Bl1NLAVj02BUejaeWAb7oKs4+gyct0P7xsCAPErHr17ue3W
dLe/ksSYWf32DtSCeH4vWM6LceFflGRrxyBTaCdCxULNqkAh7DktchEppZGnLPq3
NUPasnM1f79pDZr8sUk7q0Kv6brnDdoF5lBxyv6Xgj1IvFbsh98NYqY9WLJZQLOZ
sMq6g5Flv4cy2p+bGCo7ZrxI/k41dlkunRBJRuCNWq6UHSgILlR3jDbsH4EQw8qF
KwE7GhNCYHgISEoaNOYXdMJdUxrPnyfpFUImGQ9LqHM2IqQymUetMskyq/HWdzVe
76c+TMgtFxdPLAFvgjYSiQ9zUve9hl3+BZ/bNpsGPNy6hm3yejUIf2GWLIKQPcWL
2QgqLOboaywbJf2f5Tp5TqaFTd2o89frRWEksaspNCPn8eIMl16XGk6Y4wynpxRz
1IF3x1V9DFTD33f4Xv+NQVTPiky9Darn/RzhjiQCspZyPZWfzCLJmIPQTH97Brqo
AxdG79sbv2zAF2+kwCjwvhgoqOjHn1l7vHUQlzDSUsEfWD/UFVM8kBEX/kjnVT3/
bMs4KSfMaxLZB+fuoiiwL/tF9HGZfhOSAR6ywfKnr9KmS008xKqCM2y5yFhI+zu+
GQxbI4ISX/3fYOWtyU0oZj9TVz1twXsO780HxyyWlZV/ozwQ/dix0Rm1Gd/6bZ+/
Tnd8wqqHlWwgZqdbVwJAnNSXMY7ZWl+QSOwSbnK4KF/hodJeTkOM5fFDgu6JmUPP
6tiZ04Bw579pHoY3N2fZivzfqvokIV3I66qVXjDr37WSs5LwZ/5rQpbQyRIOLSgM
uRvi7M0/9lcN6EUm5xcODJPKVLpLofAwQOoqcGh/F+ceMsGhOthiKLppIOeeWxzZ
ARJr7Ak+V3yRHJC+ctonTLARiKHngFYdbo6ZIqAYqaEfN1u+Yw4q+wfLGACQW+8U
OgiYK+L4r8YcHJTWuQdyA8P6/t7bXwPLafmru24UY6cCvU0gOO+6AztF95YfcsjX
X4ibt0+P97X/feeeLe068W94Wu7IEdQXxgahffPj8iA14yY14ExyfXwtzAjoLe8m
dO7otYebH1rlCPVcR02lNdnI0y3LU+YJvsNc3T1AnxFzcL5X1mFzIFFwYZPNZEgU
cXmX8iGUx2R3zz2LAlrKNog/uFIpG2IvcDnVBHFn5EOgdf55rBb3WRLOkDVupbL8
Lu4XmhzGGz0w31Td34KqoUg4bT1EZGIHBxTc2Q6RCh8skFcSN+pXsAm4D3FY3BN+
092mSLPJ9Up5SBQvY4XKCXFdPvP+D5rFG7NIqj4RBGX/QGPYOeEBBOneISXYieBT
SUHTftpwkremBTotgcDLOx1qDdhIvYsqE2eC/pfqeGc+0CIuCFz9je70hCml0KK9
jy0z423C6MCDHcOO06ROidpw/DfR2hM9dgiW8a/IaPQ4ES6AJb+eqIiwEJlvq/XF
CxjH46TCBRhtFn02NfsZ2q/usvVuucj0t8/XzqQ+q/7/yVG2U4l5i6AV2AmzbH1V
0kw0rccJMm8KHkZsKSfh4a4Cgcf1v65nD3zyWuNmejAkixqN5Xths8WZ42gHCwiN
6sJtsE7rrpTAUUZKLipzXnq9Ix2ZcrAUoTn7zgRycYWOfD0bvMowhDR9Rx1y3oJg
cZPnrpP911XOxqrUP/FUmU7ouZBlvffe1u9C4HYz7w+6KGRAAKQtc5frJMEEwERX
nvrk88+3sY59zpbS7iTnsZnfGmp1mtm+G3TuefFYFr0OpTjW/A2Eovcykyaa1C9B
skRahN7QkYuUTpqU3xQtJwJ2nMPb5UKrcWCnb4FScR176Mv0eUwcbQxeu0d0YRPS
Uop+DBPyEqw6o5zUe/S/1Bc+pKVi3/9/Zz07Um3Zt/AUCQ43Q8hFS8nw0P2DVTKH
h6BVIsCHAA7XbyfHIwAa3+uq2AvsERC8tHCxwZAs3rAaHpydmpDhLu60iRRvtDHn
W7d4hFhcdf0Kfn8lmwoaacs5n4+jF8po/IcT+EqjU8c+nUtDWL1cmqfnEnzPJCEf
DpQ7jSrkF5PJgsjfpUHsxj5laybk0q46TnJizbyyABoWqBUAVfGtoo4mjL/292Ug
F7ntePwgOXEfubRw+/vGGctsNm/mZSqaRTCOV8Ik/c8t4cPdvs2OcfexmtG3Mf1Z
xrbXjL/7WdX7P+RWOrV+59E+fx3tlKaX26pksr3J6XSWIDO0bn4rYIh353isCal7
etVR7dYRckEoDaritqvsQgwhCRST8LsWZh+0AZpRmHcMvncnn6337t72iWSSbn/p
YNSFIWhu1zdsOoOY4KKPM0huqtD1NVfg4/p2iIezCm5C23y7QlnvBIkuQHRwTTCw
FmxAsirNxGqN53LMGVikHnbIQJ784Qq3EWLo/9YvHDUoyLbWZuojz+xTALGG6WMF
WHOYJ274X05XxIHbq9ybxEyNTlVAtbEY+u25qDU09mAKmq73bTUfptJz8UF4ZUF9
dzWS25UNaMd1BgnyqHh/lEGPTloJiKLszGEWglELGsX6jUl6Y6JLga0ZZ/pdHk7z
/qFOepxq1LIDrui3yA/NFzhYw1sEDmAaiuII7P/+Tu5owRd4QrPrxW1uSrWZXxPd
ZiQgFep/ihAtO3rLZ855zmz9f+3CRQl/7r2c28mbg3M/m+719P+q2w26c9IpA158
DGQYbOymfSITNllx1bd74driVlbC60UmrFdOn9vxh5SBUZ+Pb0Jl2wi2KKmj+yg3
Np3VClPO/T974NSH/BiLAQ0OY0hIufPHGRF77J1RuYJ8UoSmciCFgevVwigat+8G
Tii7dV50VsNzvBGrm+TCGcCUZr5wBP2lMLU5ZaMbjaPsQJSZDyYnddUneb1JZlwE
lwAMjqkJU/0D2315mOGh6fmjgXWbPCPcuJ+oe+KGkwxnMFIzprxFjbITKl65WEE2
jMXiAbsWAoPqsyxnzh374aVQtkkv4aKmE3sE99vb0cKazy6Ex/OjQ1Cic63zxVkg
uSpZPQXrdQYZ5y+CJN/V2ilkbIrUA7WLKsbK/dsALXDs4ebtQc8z2j3mVPXvr67p
fytZV12dczBUs9Vk7+txlxf24SYb5Ub0YAceVzMZ3R4X0aCBYCKU4t8Owm9H4bIx
5O2H0KcsNLzVID6Yy2QDLX7/GScUjWlCxgme9KhOyXIPNiBNuzkSlQLj9pqEQkMV
sa2CpEi2zB/rjlLWCc0GlcZ1JkvPisIoi22DCUMi3y5rbQIhhz/rVr96IKVfr+vF
uglQAzsiEhLA3E358FF3aBw+4/mIcNyowcbMzVCIk5mgvI+Izy0R6uIIM6Jm2RWU
d17HzhYGngWlwZqnmJO/bmRlPZWwOfpGIOjN8f+yjTTdj5bCvp02wxqjC100SF9p
brR1zYkrXIjZ3pB40Hod/i8shTOlf0mD2eWxral0nX12cZN3RCVSJuqNrFMrfU0l
8E29c/bDkbY4hqof6uSOtM1aeBJF02dAdvX+y5kBD9L6msnc2tDwzOsdwH95zcc9
DsVfGLvfzZf2+Aj6+C6aF2srOYG3HSpGXzIvf9wJ3xrv3MD4jPjn1zsEIbGYfPyw
ZgWoKdj0SBvZewHN5KLdLLwR7ka/22SPfnhJfw2vlnowhLYCOUetuxrf5EOTGLR9
HbKe54wSB+0k8Z5cZJvJvMBYmtaDu5KpprkLB0oGpXEYBQGXZU+U2dXFYGKDqXtd
QsDoE778ovJfsIVRw5PVCwiqTQJiJ5Gl4G59SEZ55jqOzaqP6Z47UP2IjRTbhAgC
1diPNVbfeDD/qFn8zCEhTiFsJeR5DVde/iynyY2ShRHUARkbO59S3uSdf/xC+Kqd
9cMz5JBAobB9ZkdHbl/hm+U5/hNnHDqb2tEFZxz1cFIiADa9ukSrxQX3IM/CTsvR
nk2qoPcBQKO3eLoIu18Dwv58Iv20wK1W4SrdIRbwTSgus/aT1lRoCpusibLIyI6G
lyhKTTSNjz7rW+CDti0uuQphHj7gXX5BdmTOAJVmCrIX61oMaoyjLwRXt3gKjBoG
2VLo60E0eYCEqqyw9RoiDm788tvmyokphtjr5o8phbN6kVdv5JF/z5vIOJzHM5VX
NdQBOuCrVQsBo3UIzXfSazUWlb0qrisEIoKrZYb1K/qr9VncJPJL4SGQIqTyDlPD
90KAHu4vn7yH4G3yUO0WAph35QndeR2xdlFlXmNodZG/+KPREeCOX/PPu6xxqD7/
sR9Ej5qB9wsaXvSo9+4cmOcsfWdtNy94vQjN1nUAmw4Z/VUHchbvX/IQuQT27DBO
Ky8g2k9jXmz2ipEQRYJw0nYPcpkspvlG4fAdoIXbazUkw1YbAm81KUxJlDgY4oIZ
24GY55Lhh1jlRbQzwXwOejdlP6iUXlbWHoN2WZZCVagVxbRZZf6fs0inpwBe+NJQ
V6dowP1KeZxfIqpQPGoUHVo6HFvyptcWqWKeVgBYIfXxP8oiBEzZJAQD42vwGEFB
CsrLljjrAEdigreTsAwybazHMrWruwE8zE82EyfG/aZFjtRH4RDX2eM/SMJGK/Dv
e42i6cFrwI3KulyvGLOjYdF9rbnjnc/RW8pqw7dFz03cnpbgzyOA2/++LXH/wF0m
FO+zL/Sfw2TKArdr1i4RzOq7Gu3eDasFw2o/51c3qhkN4DfOR+mnbavndZKS1oXc
uTgOdwG4juN21XP0a66jMLvUp0VmfOHWHwDPyGfHKgWs8WHKFAC5HXXnvm/f+NPJ
eTis5jP1veMDY7A+oCZyyAfLwGUODTcuTFbBbP97wqOkhT7qG+JkX6Zf7LD9r1Yz
9f7Yuidz8X3FnAfgrLwgsVykr34oCYDWkgfhNGq0OAXJblIvYGHSzBwf9Jv3eB5T
vlgbIPOmrB97nGL4eoh8fuQZFA9JgEJ+Sj7isLl6vajQJfQeBBxXgEMG0lcfxSqe
rnrSqKWSkLhKgF8CtRxnMVH8XBatbKH9KLcXocTzxXDro5YZLGd0OqY0PfuHe1J1
JxYR79NJ9ABZ6sN9rP6ylhjfh+4rqIm5yqSHlllxb3A8ArOo9rCSmG7DvA1IDGTO
nhINC/sFk9CcPDjuk2qf5owP5yiSZT82VOtnqYY8ikOFzplNYGYDCZTjywnzSRnr
5t0PtQfigXEF4pSl8u/cYmP6obLO4mNIO5QKfcGFbDcZONTBwtaZMwDT+lXYEbVn
ASwYxCugwrN3uBd+5aA5duMYLxczOBJdm+XROUhM2e0y4PxC7DY1avAN1SgOZrW2
lI0WfgBp+vM1BoZP5KhSGMbEVmOV+Y4MBcKOogaVnRcH6acUPdbnywvqK4qoG7+i
gF0yyvj13nCTLW5WWws/Str9zV2SW6jYPP45OY+gm58u3EEiMzYx4IdKQo3XwftC
k+0qKE/FvoQlmy/4/gr/783xbRR3pVGjgEw72S2H0MjdT+2umNgSO2wwYXJCdBPa
uddZR9IAil9anTODrhGl8BPjsbJl8f0MswuHUIHk72iO6wS9DNG8N0e17NiINQYM
CHGMR5+TU1qkfuXTRHOrqMh5A/koL7QUi8Rs40p/XCjyVIbd9Ng7wQWt4x012hfN
lTMYslsxPg1mfteR5iZUGgZPS0PqkLqBThMF+Iho4dM5d2BNqRuUNkfM6tkIQH2S
w2xsjT6HYKvEbXh84qjx/g8J/MxsxYUMrwUYZVpQvIxrZMDM9V/f3lXoTU7Rlp+i
E5/zXrzq74x8xlK4IC+UfBvQ0CYX5mS9X7I0DyIAyMLjjRj51ZJ/KDZWu+Emglpj
XWrm2ilqR2x2wU+Ao98/e7P2Wan+CKiNeq3nZCHzEKI/YQkg8GRNPEczcIfj/O8p
InHlDYI839h8Dvozmjg5jVXWwIfEna+ugb2BLW6kVAE/W1b5+5BZhcG2d4KKZMDV
1ovQ2kiDyP2e9M93Ga+gylfpyG54lH9Aj9WCS60CcTDVb4Q0G03zP5c2MPlQxT1s
PRkmAghZWX9d9kylead4PDQp329qpmnICArB9H+GnxTk7FPeyJVnDumsS6pKqmDQ
9axo9pQmOVDo3eAI7QxkUxKrk16F/I13rd5uhtJk7VkF5C4ryc7syyUXzGWqsm2A
IqGrkaDWiGB+2zO5RacT+kvfaQW6ovLQbhKDYqie+4WbDm+Mxd83hslaW2x9jmN/
VlSVpsItJ9Ghi3U7mgmb7W9PUJ4cQBWbveV0GXDfEKYnyqM4LCuzoyh/kp+qbeui
nPWDA5rAse+ZTQ2z1QWM+SwIs66WT0MMsmt/UbPvbGEH/YuBqF4XwmfxjUkfUTFP
hHt94n8UGY/IQIePlmlnfEkxR7bXQRu3rxs0ahB0PYBmlotq1cDDV5/r6l3ZkLBb
5iWKK0nYdZJeFXRSTvHBBzqIB3yvwjT3LHw5TGoRqUc=
`protect END_PROTECTED

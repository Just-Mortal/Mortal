`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7lZAOXvfsCRyrUXnkSIVqNkHtb4sc8JMx2ZdrjeduYP/5QMsU0RC+f3tNuIhV4wE
IvTKFoVV8csHDzuN6CxnRB6GpIoih2xNttNfGHMEiarhy4yZVsKiehzGrFW+1ZX6
ncYCN2iiB6SCx0FnHBMjZbRE9uRbhnY4VTrOgulxFFTgK8H6lQawcMVkrGfQgRTu
Y63Kc42qWWC3wyzJxQsWrvcUmPMtq0+pU9yR5l3ItgH40N1SZaos8hzReDrtga2i
dZGG0Pmt/slx+AHQxhZUKd2CHigFUJDSqKkphc+vpyIhXC6sTrJaf5CAq4VRjavy
jzzIwcM7J+rI6rLNv3s9kinCaV2DFoFffLzNA6R70ot7NicuGBK7BYaEWLLMF2Qc
Ttvamcr82dbJmNbTAxMACrDkpqGNHjZuH8tNitUTXld9/gZNm3/zLMCmqxi9zsx9
+qi5HDn8TJsVo6PkxDpuT0KfXiYczC5geqbZeni5eeozbC79ogVKoqMWq77kl49o
vuXVOb5ZoGoszckyXIRgAgiaD/lF0ZuWYtEchxgMmgLVooNNQY6nyJKYCsuOHbU1
qxW9L1VsBdH5Sk1PvTd9HM7eRmJy0/oPKUBLw4HxYuAU4kGn2cM5iXQ8/UBREXHX
KtbPZrIknQ4gxfdLexshpxubl7SrrGbzEKdavKesHbvBy6nGAKg0jMnMrXqM3H2o
JsnOdjkg/BM7mF2R+ht1fHuSBeZDiKytUMpIvkF5gOGXoob/g9zkyfntLk3B4hzX
Xj2jzISYOANH4wIFy4U40oQ15nhXHkBP/rH1uKR+mnr6DOYfqKDcnpg4XoOp8PVE
Xbi3JrQh4HdBQc0d3ypLzXp4wxULpRDXCuqtMsZOgRoi8xdONYCxKJn/68whFIwy
g2IVuaQWO5UVU0HF//JITcpnP+nWM7DgNaMeD7Gfjjg=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2/CL3E80INODuSbwaFT+0buC/p5Vmymoq69F6qq1SAHVu/PRWtAxrAqc55FNc0d
tBRq28OXE+lDycdOBtvkfmMzU2O/Abj4jk+9sfki9VZHcmRFAkk18C+4OF4olUrV
rBeYVOtdMzxN/dTHP53MQz5y1uqaSq/LsIWQe10cuvmLADWTsHAX5evq7IVhe6Bv
b4lZ9P+ItDtYH/UUXI7uY2AJlHBmQmhTE+fs05OG9ScZn0SpZuRCAFS0OVjUXMFm
bV4WjxDW1wl+YUgh3exXn7jFh4SnJShuX4ZTadfIZwTSMkteJa5McYPVKJeL4KUf
hjCTS2/8bmTdh+vknipbmoTn0M8xnUiWmo7KrzsCk5QQQxO1qlTFamk3K+3FlZZH
n5/zF5e/azm62Rv9q1H4vWF5vdkBjGSANf6oVcUdCf1r2xMbTc3wYDmnje+tQMHe
zvsWkFhvvpLBpwWuBgdBhKAlS+CmG71pXK0HI7keDc9PznOK4br/uuUHPNLXWS8t
AlzYjRifpbNfZ+RdCqp/zPmVoAIZIIr07YDfuWFAzJiNdS/QYVwmRt68eJ9ayICf
JqoCo5ubFNR+aWnZFPHve03gvIL8siZiDDqdmbU8M3XuG221m3pbblaRlHTTj2Y7
0rugbyzpmQOzwB5vB+WrV5IO7jXhXkjX1jRp5ixqNwSS/ZRluiu2WSSRREvyi3mc
F+FjtRsA06epo42VDhdk8gN6bWLx1uLwaQVoRofL5NmoJ/BiUtiZbgf3/WQzujbo
QUG+goMJYbfKdeKG0KqvZKOAlduavPmuVzM8Q0dUQWzmMf87kXyDfrbqtur21kbm
IxsAkAs8Dvrkvrf0hA6hsw==
`protect END_PROTECTED

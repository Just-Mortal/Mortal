`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wt1eP5D9RBqAS64dtuwGkBN2s0eXNMHOkBXE6QmG3hdiBllsZkRxnZs0IFpIssu8
nsKsf6ReZaxVnWsIslx9ZkUCpm0zu3e3xSLffNLPGqWN41ZslDQix+ral5tLKYYE
TFZjkG3sXQX7IAKudntK3i+77dZx8h+7Xq002M/JQi++pGsqtHvYtFHLyRP4kEy1
cwsuhqgk2X4VMfHAGv2FTI4tI6umJU127zxytY4/NhZ+9lhfrvzgAUuj+jh3KDlD
z+bh2I4pbdXCb9bzgOBt3e2YDOVoquvIvebVyZIxSKdXErHBaCV8c3MAFoJUD4x9
6QVh212BdB1z7C2SCn4vj+wHmfZT4vPduue+fb3d3SOg8eMYy+fuXPoVPoLat48j
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
um2xGEYcgV7Sk//6vvWjlsdjYsmYvCfq1tSlGiFOcfv4l2XHPJ8ckSqiy0rDbsa/
fTJecle9gV2qz1kXDe16XMMZlSzlECY4YKSX4bcfs9tAomC4ed1EiDFNpo9i9ONq
kIX42omUYMUpaI7VgvU8Pdzj1NdsQ3bQTngxekh5khiU+uxT1XeyaWa47BcwQfQw
NND3BPQorurxVjgg0O8ErVMZAzAd0NKEgSD4wt9gw9uotKb/6uy7MrTLSfs6sP13
006li6hLRyfG4XW43tpv0OxVUtEz1upIxBFuRmC4vAet85xU+T1MHEFLIrifFI9D
k4L5pgEi0byT/wweJEbV3LEsL/TBk/wyWozTEsuZLltpt57F/M4k7OsHfy5awu6s
igX6axOqOHVO+QsyQf8bWmjPIsq0nDiFcD4iyxLTmTFEq1wVatbTq0BFfg0+TzMJ
/nst9x0wBwPP3OJgMPtt+klmysTHGWQTMb7KouWLq9UNHnIg3YcqwTYRnrKDbsLy
L/L0OomKeazOFRXVwhKUyU3wY+ayI6scKq4zOgqMvlCjD6EG3+omxpBnRaaAKegc
9T+h9wUAsp3+YVdcTyVxqGlhFsSwzYULwrlFKrk+Yvklt4NZrZ3g51ZsOLprGSXd
ubrxRMJ7h3P0NG1gcxhN9B1D4dkB+EGzCUyebKp+3nLzFtRH1zylStLI+F1kRDB9
Zb3IrNhUIR7k8GG6cg43WQtxjsVEtkpcxpsslUOvcx/pLh9nN0SGSPj2D8Jgm10e
6xVwUNjmN7Ce0dUbn5knwQ1mmI0PrmVeXfJRxmzh/BgYO3DqQ8S3hiBApiTpfMZQ
DhGT8MZ2NWbN49D4yEASnqyGw6LyuCfMtLg/HAxVAdyRiCGoIdkufpouPnY/FffA
Vb8fU9+Zc8L2OFbCfxqTzMzYZWJ4T8VnBTholLMWmQx2LNj5qHeUibcMxc1WLWVp
sBoxef30yXmTieGQPZNuwLfG8uDpkd1cCviwmU8O3y5Tmzhz0ln5wrNvbCeJGwfh
r3rC7F/Y45Wnp1Cts39NW1qsiEd1H9OF/A+f95wzsv4KyycvguSonp3rq3QixHao
zF0oqD0Tb9nqRd6Cih3HaAiKjcypsLNCt6OC9iCaN/sGz01zJo/C4yGNedk/eZ71
zkHXEtKXERX73vLIEIEkDg2XZgZfDs1ghelPmJbkaAfJlIyK89epISirTVL2jGSo
ymlI25VuMYRpEFFCPgsmcu6OhpL2mTwfsKFptOYL0Tp5rGC8ubSZrPptuCZpNqzg
NAaqQkr4Vi0YR0Eemn3Mh99BnP9mBHS1M3vdNACcvqZofS+w9rIFszI7cejgP86j
e5E9+EiHlHbj9S+lUTO9yfTWR14815OKjS6IJhZHyimIRIrASYMs2mGjBM9DZ3CF
EyMXq2hWiXj4ZQXM9nD33VXOwH6PnhMBD2VgNUKyKiESxQjZJJ6IZd2QeuNqrsk2
ILGKE9npv7g8wctEFqcAFmCZRHy9rZw+/3VJpF+Xy3P+FdPOUhh8lExPNs9YTe2+
acT60/jAZWoSe+fmauUA7x4Vi+4AS6bzihgPNV+Ap7HX8TT93JE9EGOfWif0NQOb
7NjTg/inajMWFl91/VbWsq9zqordSFv+tbYFCvrj2MRoA6XNJXxdg4lylrVdNZG1
ji8zD6BKEMQHnWB+PmgEvmVwsKNuhQMSlCvUa1QzOBCM/5FXzmUwWVoq7IbXjFB9
PjSBx46PplrP0PwczmDhM10jEaloTmedXx0//vYVZ0VgFM4yIId5YKZl4irMennt
ZTMXAfrcag54SwAjrd1B+/QVqU/zgW6erIrBfEkJL0pRMpXXOP27+2qsn+7wqVZ2
EsJ19ev3TPf13P/iO/wa1zCH/ZQzZoXmlogky7RqndmTi01DeuN8ctd3x4SinK46
eC0cmO6pF5p8xq07ucgIHETJd2Dtm6LtYk6pSEulHDg4Fa8w1zsye0NDpxkFNcgY
yFMy0KlX/Tl0LwFSXbA/YlrAfA9SWEgvB6fazQzz/LQ84p6EYQ+N2zz40k6sreEm
Tx5Hrdb59YPPAE9bBaO/dg/CcU2CMwNFisQkKLimEOK8DMdGvoluu2YN/3fitUlI
I1cFx+6ztJc1kO3bXdh5WpD/b8JnKDxK3oaV0SWCL2UKuTY9/wzWGeB+1dQ78Fda
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5eGWhMGR8skwzf4xhestOrzZzF9MMdQnq4rES8vAzpcCR5KU5uRE9IrpXw3WDDAF
ZVdwQspD/0mlw8ATaedV/jynzT2p0T+Nicp5uWiEQsoWEu/uHfMCQlvhmd7PCB9D
LFb0G73Oh19G2vjAoEN4kPHTjpbNtdbvc4JKtrWrw2myRNCmXsTN0rliiXYbO3t0
HfuO1MKBJVW2XLIdjJsoqcMb97t1IAchBW+k/IpdQPI9hx9cdct+2dVC+6Tbmfq5
taRXwr5ePzb14zne0k/d2mlaJWwDmrbynrY2mnwZfUmmrEepAhzJhovRZbho4XRm
52v9T4fAo0+T4MJPf58EzJrJHdNtmPE8YssxCLfTO03Rlg4zS8BuKnphqecQOhUx
mzGcJ1zBJRApsVs7sNNDZOeflUhuxjJ4t8KZ7diUUc0UgSA/5ikSFC3OIl1uDqmS
i45hhF+actx6ARC367BFQWHn4JgnwybAUrWeag/JMyI=
`protect END_PROTECTED

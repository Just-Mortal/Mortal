`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sJCh9YB9xFK0NlvtDDjOxkD5ZcAtYtUsCRWUv5djuMLZbIUcGtGrfusrnwA21njN
z072T3drdF7t7eBwVSflAc42hgnpifFiIG1T+asUvkApnH7hkEbWwA3wvlEzhA8U
lBy5M89HzhOzFpnWplNXOApNsvyPWGxEI7FvOCPcVj7w7lVA+vTTLtAwFmXOuMee
w6AXbSGqJMu83lKD5X/MEbmlrHU49J0FACAfN7BdM50Kjuh2Sw0W/GbNFFdYgcex
DuXAy92djFyk3aYOw19TibdRyUZEgYue7/hgc/YNjfhAsrpUWuPzap/L7JucPeMk
myCzOXKC8PM9q+Mbug7uPxDEHbYmIYXg99iEspCLHKK0kYDGUizGNQGX2brUog9R
umgywxF/Ehrde5Eh/Jki0a+0TQZPCNIIngCIZI9MHNNIHrcrrqUBDIu/KhXTXfa4
dpaX5GQOGGHAa/NoaiFom5vQYc722Sai/g/Qe9sPaSZ0l8sAzCUwm4kRHRsz46ai
zFeG63Pp+oCx7PM4UxaaF7FcqX+KOyessjFOzNtR7RmTjN6Av4R9aQsyRV19I15/
gCypTalqV3fGPXtBdNXnm35ByPLmHT+TJ4agZy1dRzQ+9CaXhV/NgPrdWHo8f2dM
BC09bqteOU2HzMS3URZcsVEd/Yp2AlC8PSlsS/XJI5Xieo9tNbJzu/DCTSg2e5fl
MeFJOqT4zReA5EvsEuDpUnGvj4Njo840l1hDouGiTjBwSWAP8qT1aXeGF9Foq1jh
Xq92l8+ovViuy9qMC5BIo/9w13wJZ1VX9wxu8FoMmRcDFzqu9mgVRKEilSX4ZLq9
yuyZSpIAoothSVJ3nZpcWhyeeCjsFiLiKGWIaTu//4Xts3MALzW+4NSdEJO34S80
L07CEMtWxjAEuX8nLQD/fE2bDj2bAJAVdOTeuUm1QEWqI4CdHNPObzkdTAxvuU0c
lsyRbCcKfj1AiJPaBT7MRwKipqRe/wcOE2jTOIh7e3eZogbX7fkE66UPWZ45ouK5
q0lUCrDNcHX3xNxslWH7K0v47l9MV0jTMyqdYEXwcX4tUU9GrU/nGxCya/Bv0tfb
JV7IjqGNAXvEAPi7wk91yTxDuAumGTEG3Va0DGzOlybPekQA04VfXtPSnIcT5owh
kKJ+5XbBbpBlwfkyMpUvN8NCtScAPk8lLZbg6exUiIW279rz2TU3i55rNmOXdCpS
TYvhp7x0ZSAJ7ElxyWhbp6nt2vt7exGCmrPb3MXXPfrvYOiau9ylwsf6GoyUID4V
ix99HhPRVBuST0uN025Q0wKB8pnSCNg5eIWcQvhMRPfcBDeUrfasbli8bX945+eq
7LkMjRzPTkH7GKWAIrmxFDk9k08IKMmjfCRnEyvqVFMRpv1UpuxS6ql4uYLXPCJs
TtskyviVUh3hW3cJ6T78KJW9xxaQ7RaDB/s099Z8ji/ZKGz61HWOpsAm4qNuoxcG
AGo30OnxLIBcpKAf0EvnOBASXdJxb/6AwSzfxldwDE0ID6bnisSISiLblJt5npqr
ur1aN1Yczt396eBpo+oi9JmKFtiU52jjSArKQggr0PaX2Se4JicaGapSHsk4AOCE
Atn+ccH08x6rGak/eFIWiJD3IAQvgxuhNuGyDwW4unNH4Yvkg/4Z2QcGhoKxVbAv
6s6vmm8/ofHazFkuFXZg2e0b97tEvJo6m4/T5lfx3zofS8ys6Axt8nTJT0kMIdB4
S4h6vA3xeioXwB03yiYO6ijImU66SNPja+foHdWjbUC2d6TrbMVTQCycbArtZs0p
LFVOnFatMs0kBmAPd+25ciCsJHtiNBpZTT+Dz1yiek7ACZOBi9ywmZOGFuErj+np
KPggiaZIyrggcmZ0S9bcAvN3W7NKujQT2KTtGIGJqxW65u+uN96U6jQaddVQ0tJu
kUHXtmSzCcQpCZfuKrzjEMUcIs4lYv0n17PDrQuDI0/yX6DkTv2zCc1S5Y6a1H5Y
jSqnz0FNTIGEhFRLThv7UVJHpLDXqxDFNm42m1hC9QCpuFSYZMfLDAtacl7JpQWM
FuXTKSsAIeIbbXyeWEquFC0EQbplwqm9wDb8TI7qsTlbDduvBcV/p6McbSAUztjK
0k+CYbaKzWDQD96d491vl0wgkVHKBUW1pklqvrdSW5G9cpckXPZAJT55TaC4P/YH
SJJvx7wfFPEzIE/k9fnS/VRNfPLiiRUNqNtkpVJMK3TPuIQFGXhFMXfT6Bf1Sgr7
7dtUnyPu4XVLFL1WoXdlbHDcUQNOXkGbp6HW//KknEeoF6AELq4pTH08cB+WDHzN
ApW2VvO+yxpbCrVZ87Lev9bcPzovE01PpVdloYexnszFEzGE2VIwIvzytOvtcBsy
Oa6GwRiAZRfzb+ij4JIaotrc4OFeQCPH4A2ucg2goq/VKSKYa+U/ozRJYA7oRV9u
Lidzi4tuqp050b5++VQ4efDxLbdYApDsI6LPqJdufVgrYwmbdPwV6cbGQhsrQRbx
5aQKmAmNz+WXzbP8K0XPSBvNKo8zue9FLdXt6ttrkfaMuVbxpoX1sJQnkNuTzsZ9
8yaznmY9r+Kh5Ij008VrqfYQaD7RKPUIHpnOT4G0MFTtecRa/ZHifJx2iR1Vi11+
jnQMr+kX60dhP5wutXTc9iVmu1I5Qv+LPIkFmsj3rxUsfaSNgEE9487H+XtFxiKO
4cC4CWdM9dFsIj7eupkKSnnl6x3El4diDFuNX4xxJL2YQbbHJ35NBDvUhquBZzFD
k7AB8aHmqb4qYKQc6wkBTeJvPtqbqMGAxchCaFvloMHEWdEVaLPQmRGCaTdbQVkB
86kE714oFIqBGjZyuQLa0xk/osv13s7svprGFeWJ0Z2pgmiIzy/wtDrn7m37Pd1B
k6iVzuGLTS6+loDbIzZbv7O1pb/L17l1/2Ai4hnzrBZdT9UYRPt3p1IvgbiueH0+
odmdU8o98QjraqWLxrElELWavJROGZkI/Yb7jOzQpcaKRSLYPuIc+2FEbKMNbw2U
aJcLe/PhZ5ouhPRqq5o+3BwaurEPKVKNLrKdo1sqeIY4HM0q6swKS9DdheSFBCgM
ijFv2kp/KJKQrQ3pzyvDADgVOHPdBv3wx22kPf0cdNslvCEHBePJM3nTjmap1ftj
aa21Mu3isPVo//mQtiGRaIj+V/zguwRw2ZYuxr2fxo/kIkYjYkBCHYnXvqIMCigM
ybhBgvVlfjjnkqnAqwyIy2zNUXCMKI9EaYVuOIHQpxK+PwtPvSl9O+azT38iEH/1
HszPguW++wLK6UktShKs+x03QWtHz9yOcBxl+KkOTbEU7olkTNSgv0PdYWFWKc7c
OKwyq9DLJkhCZOCq4TtRf5iOE+w0cO2IHPEhlEC/nJcXLBYhB1zCIEglsGEs2yyG
9MXmwPQ5Z+6pu+pSxTlemynF0HVraMqiMvbhuM4Cbgf1rA1Ry+g+zrAqlVlO2LcI
0q+BklOL1mQsH2/nPJly22bMwoLQgTlnuiboFyLKxvcvRKSCnftq6XH1sd3NcWjD
kn+CyqjjyQfng3hkfjsXygwwoM6G+M1gAiSGBD74g0J5PC63NxsLQ2CyLJeVobAC
HJ3ag1MLHxSBjFYm3ot9yvWsiZNtxOTiHRu/PwYzEBLiEiDicI7ZEocn1nkU/F3d
ZwTc0D9+W2hRbFvXqjMRJiYFBGogQJBNs3HakzuNuAglGe+xc8aKkxSVpxeA+Tos
WsxC4gM9LBr+Rjj8sdTh3gM3sPZDCc2zNWYsqSTb4/6v9dvLVOIPC1OJSy1ZHNCH
NB1YIQ2ctqk14ODZLGrzez2b6XgrSji9V5rGMBFahi+kL2U3244EcNCUesshk+ZV
BdHEwxMU/0rCi3w7B1V8sOhhKBNCL/55ELGm6+eKXTcNF5xsluBfQsrVZdgBqRzJ
mvxby3sfYPxAY3ZYNNGXBdmcDHUOVTQC4ormsf+00+Wbmb7TTl5t2xF+V6JwH+Hm
n2JElP8a/ZazXKTlmCR+sVP8MT4JV34UYj95LMz3PDuxWqbRdKSdrXym4w+HwF/j
7QknP4i5g3EM1BZMusKZjzjpI41sFJfLR2F6Gqjx/B4YKk/jrDkKhUK+aUcLCOoD
HeIPkDBFqFByrhhnvhuzY6ZgHFJwqH1si4fuLH59LnBffDwiriD5tJTInsdLAym4
tFfW4mTI6gKYAR5tbFcTA9k/ojoodgegMQazrxpZWc3HEQRW+JQPxZdwslDffj+O
m8K8Vo88rVxaP91eZ6LSXD7EQ3xvBUaj0Hsg0ANNt2P8vdW9MVowbG91G+9aMfU3
ZwBrI4aRSl7crvdv677a8XLswD3pyN263z0/lJiXpQf2aV6HNr/+htk+9qDQhv90
xqiHwFHtxAP6BRYTKyWVOr6jEKWOxGJ+HQ0baDhoA1HlIPEyCqRyg8XVF6I335HW
mWuAoaRWvW8cs7mbLn33gDBIZ0aPrf9TPL/fkja6sDlocxGX8U++9ppCJXS/s5tG
1f3xxlN/Uy6Hbyu7sGK2xYCLK2v98ADB5cvZga3ago5oiHDqFYKM6Um4/v+7pZIg
zyOWM2AiIOAeYbE+rOqXGECGqDEK900PIOUcynCBxsE1eHVKTHS0TC+KYCik/myh
VoSGiBg/qidmWpyKAoDfsSmgqwNmPBiDrOPzlW66FaYppYPKrEDrAZ08K2hRxrmP
dmd4fQiUaOZq09ii49sZ6CsQmOWgig8r1QVe5IMs+3hU+dEW3ZcnFoZkl+omSAoo
o67ZQZxhUutQlrT/ln/S6dOjyu3jbRY0z9QI4Ri7deFNk4Uhl9QzaGakQPrk+yok
bpniu4yMXZOyooB4rpZqNRdlA7kKD3DpIDk5MLXia102J/ZlTtcWiUI03w+gOe5F
5WXSUhamkGMc9UjnMyupPkSvZtFDw17LroPsiT9jQKvCZzEFvxYC7skbpuTYaSX3
5M2htg40smPFZYylgnWEaPF1oTgoxLRBNVd7WcRVCuu+O5/LzMaaPosPxS2t2eDH
+5RueBl5XVySM271aLxsCAMUO8uLISqHSooEt+pGtnqmw07w64KiliqSfBe1+Gyy
leqtTSFvgveR37bLvI/8NHiIIdoTRXpbCXkMs968ytudiPVCf5vB9XAZvk0iY3Kj
R8MXQh/JM3nd6NakSOhpouLfe6+qVHjPRY89YjnGtdNdRRy0ztUbin1fBviMCglN
k8KDVvXYRZ0Nj0ANF5MhccjSnrq7ZqPGxAlE8/w4j+8TCgT+Z9Nz1DtAwehuxc1e
NwLQXep3RS9riF9CufS3MzPIbe8se1qZVzKrd5B9+Eye0aLtdcqNd0Qe64RDpkuj
niHcFmDfZ6bOfaRbZWnMRojVlw4dPyR22nFveqiQHLsSw8Rpp+P0qeVKmNO3okyr
kXfvE/71/yXKgM8oTN0wB/AnyV5JtmEpwDb/d+LosVNm1EQZJXAjBmDxirebvXJi
YzDIbLgU/2Jr0BrnaZDmuG3nybRV7nyfj3PC56iX2JZbxtUeu0Rx9C/LtN10MWmv
MPRHuMxcOdxKWBuhP/mHcY115mPEgwK4MaK35JCTjd7veQD7wnIj6OK1ZgVnLEKM
ArL4XiwvgYqdaBNJkIq8wEkDkiWIH2r3e0pcoNDJlwBT7WKhnZ+bi++aU1l2Dzmp
sIfVgk6QAZLa8yEEcGdVZp0RifCshGMmZQOV2QbRjqIkZweVcaUmctV5xiVAdP8X
N3o6z2eIpnPWrH80Ia3oYjRF414JS1L/iLIy9f+RBy2rt/LSasCLGDS5wAK6vjbe
2hmrit6itMCy/M4kkP1z2rHO1PY5VigERy4sGB+fEEAYW7cXe4yjnpf2JuuFqHd/
hNp0kATweO8TWW44aFS9LfciPPHBnfoRu6vGaa3vltsmWNQloDg6EeVpjSwlTHFU
AgyKupxgYu6PnEGQlDOPsQb9adlwh7MtlvibUNmXBRhEI7UsGkKJ7XE+SLNkw+Kx
PJF99aYLcpR2/D4MAWcwVnORWydk6KQyb9Dy29ApWpVkJzA+qpqI4fvjQsV0Nvlk
DQqlYqwXlRnTExGK8tFdoOSnXlAoKwa9txwsztG9FSJcQ2jQduUoWmKijupWGTQK
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fN25dPOQffHavSKVAbMbH7udeSyDhj+pdO+kbo9rMSfx6LChlAGV6RKjMxXSPtXv
FzzDQKPhSOtgshsMEXMOhzf8AtLWouoCp94t+Mlxm+jY8BLE2ldzYC+l2iSGDBwM
ymgqHqYu3UL7frtEuthozVkBn63Ttl6Ymch0GXciGYQ27O6ySz1yUhDK4HKDnrbK
72MTLHEDg7+bRIXR6DOo/Q347iT63Ls+VwsvOZDxetrkzEGLJUyH0VXQuAZCf/qO
9Xh23jNXeh0WvwHWFZTdVFRz7Qss7JdtVlHn2YGpqE3273tJwhMlwrdyxV2gEyjh
Y52Ir7AIOPclwjqZWr/XBHVDsuo0WqaQ2ikZJ0xF6HdwBCtW91O6uapKedoZX2zP
eD5Ixy+cKp4l2ixAHsANzY30BLZcGQRaAK+yeVntpp1CGpZuU8BYREtvYG/Oug9o
3m+C2K9gQkSw8END73xlQ9lXIrYJY4S0n7en2w/XOdat8TwgbA9r/o/TApfFtu0H
vuq4yvaaFu+JZl9U2HlC6Z/fatG8CNsxBUvCbLrEZrf/z+23IYsygSX4jEqkqoqI
ua/a+LzlzIQmNXZCiVGgFNRi20kLt9rMyEscSRsDE+Mg5e8MgTCM9MZNitk6F1p2
XZvrvKCQAMGPzxmtaPezAbRzKqr7wQjx6RyeMNOqtI1ttZVnn8Mzfuou6OpEvdLU
RGiD58HMzF3nTnueQj0ppnXPdzUi7Z9ds/3eo0nAO1Aso+kNspe15kdNldlKifux
QSXBb2Rg8/ZL7RfHBod+qq6I/PLy84ARp40ROsb2TTOvWCToZK7/PM2H7KWzxgAJ
yzc6VTT6XBFvPYV9AKX1qEaOx1dR2SX+WGlmqNn2rg22OjkPcvYzTOKoXDehlcLx
YnxDV0369hFwc2GYJPNsOCrRqwlovmB8cbd3sLHCMGDBpSCD9C+1Phc2YUiicB5j
r9CO4g6o5oi1+v5dK4amHlWLLqhC83EODgCbZyiwaVnA6Gpc635FQ6UmDLs/WOUi
JtEy6btyvf49g+510HNVqOSrOJmuorA6VSudDLEo3Z89QrA644c7cF443HoNlkS0
5ZhOtDCXqOAnz9ZsHgePVsYqwVwWH0ovL4pMPqbnTfCF8CJFEOb8AaBk4+z8do+l
2C/2BBIK7ws8RucHV+CUKr+iFChWX8nESy2jai/xiD0Qdo2bu/zmrNo9ejy6X0j7
UMvlUjEWFDI+HNGjprdflBuQ051f4ntjzXVEEZ3lRIhClmQus+xDswtS1QmSgODW
5jKlN6mAqc9Nw/4frTLakM/19qLjs26rWccHT7zrgKgsOcKpNxCRNmFQU18lbLkp
q1MRUcvbxzCQTiFtuCO/CZP/wyIczb9tqZcmcB9F0GAyrmC8/4nML7CDRvPQoDga
ewV6/QD4RNlDBwVwQZvld1oRRMsdZHTuT1gJJ48DjaErG3DuA733r9lDlA+VwdpN
V1epIfJGaoxSZ1KqyBjUiCELybTeOiCNbxnKu8z1OQ5Ie//6l1Jtm5DoK9xlU8Y1
b71xaQ5KOD0MYnU9p5C/9X7pkIMRu+QDG3UKo8CppzJX4xWISEXmHbHUHvd0/Xf0
cd0hnB/ldGZSvc1OEfDg+yOPGNkc5zkhWQapLHeRgjz/2lx2aD+0TdQai/+o7COi
DCwpVBUdefEWkre/xceDsBTxPckzL/4KvALIChPYRrIXTv6atUHUkhr3UQCnYJHa
2gziscW4vn4qOcmbPdWVP8jCfs26kzCIzV7cja4iZL2HZ8noTmf46IqRtmODqAqn
8Ave6g7iT2gC/eqdXisErHxhChm6DgTAg7bfsB3IoDBv1+IUhMQ7okwCTEy0/Lc6
LNlCHuIKYCDugatAI+kEz1tF6Upk+LZ+R4KDFGuhmWG8EJ7NNJx0KTGE9xqLUZBk
fmIqE3iRJ/Ekl/1bLmxmehZcrCK3+PU7g8xeMAOU5+p5zQU1YKQg9mceM5LFIYt5
5+Hz90ZPe/jVO/vwnHiZ49K0UJsW2I0blC1AZGPfqH+S1pDNjduxlRhyPyw8Myj1
3UEEpiIBqeliL9nkM/Na5F1jPXu9ZHG3SxyDK0jDJWMlZ2OP16Nu8puSI6TUpicI
Ro+qohfV6bqQtKVBr0hlrFbL9vb4caSmGekXHi/3p/1fF69+YPlOfURywXOdx8xI
Fiw8LfRLyxaJVsmJO8LoQ/JrUik2/G8Psjfdx5gw26yi5L3WiVlR8RuaE2hmVLc3
i31g+ruZJ1S/qVeLx8nlb5q7rPQ+D/mPBKgg0/ysPN9HM5Cv3NJ6OR72ORH8hJWu
qpzytq0W7h6Sw5U8u20L+84ajMXo6Bak0aGQnasUGRjoN5UDIKw2BplwaVztg3ZG
rV8K1PaRlRr8dEYG3TIpE1i9DUW8pU/D/B4jL+aW5GDPIB0jQ2URPq3Ajudw0Jv4
4Qft4ybJZS7izUZLJy3lZEz61w9kr5uhIealkq7PyC6XqkvZOArbYfN320L71ZZA
fOx2Z6Xf2P7Zifvx1h6nxrgBa0W49o2bAIw72pFzL7To0MDBdWxLcs4F8sB46mZy
0W57isAjYMVSlo2a9dWKM2e0qxNZdNFEcV5QDGnhyVXAhgnJUHI78LlQKlmKIjmc
vH5O/L+cxnYqAswori6XmDrUU8pyPLmv6o5qYu0EX75bf3j7vnzW/abtW2nUBs/O
yyanRoxiRxdXWwAcWgaP+J+Y2IrnfPSWUu4q+LmTMO6yacJ+qXDIGDmIBZNQ0OxQ
B1JK2F9aNIRXImx/dRAkt5naunjoJotwSu4g3RMVk88eAtkcxOKYk/nR99q2H1Zl
gqvJRgjlB0WoU7v/WJiuZwY6IKaW2NpEG7+xSLyNG/3QI6oCVsiqRUBz8+dowowv
jZt7BPgCqsUUjPPwf8w79uTkNbMI+CEICt+HiWfF0XDggU4Q5m/OrIA3O6swsc5x
eFAI4S/ld0f6ntG/LMz5GeCXhKC/ZiX5bTW0eiFgxvGJBYGuMkqtgIgVpBFcVb4Q
8A/wt6o/nTEIBiw9ZCQNOrKNaBXGd6M97pvCQfXfx/V8WL8J4uAw1ZJTR1sHb3DB
WmFGJA/GCUSfafvt+TYFyazDbX4b6M836bqOha8oCAC/FNbH5faurvnt9Bla4qTJ
7MsldzqMHOduM9vcTm8KO0ljTDNKcLKdxdOsgNsLeIj0obnpiwFnn0V7RY06F61I
B+h4RO8/7pRt5DJ1neMtSSxl+CPuaaBz1S0M0k3EH4FCFZGntNgIE9l8QaIxIAiK
QwnICoIaKJfY7hQ3YIUDFmqUi3IxuUf/YscioXLNq4oTaEq+KJLQvRl8s1c0Ggdk
s1FrOlbal+5sSp/dUCtgIXEU7EkSuMw+17XemwmaIB18tGpnCQL2LPmxh4ww4EFc
weQtarbjv2PJewS3yJE/L0485Kd8CDEdxeOqETfZdf4StztL8BA+R0K5NjtUg4fB
QjvmfaOIWjZa/BOYVZvd5AJnym3knNoY9yrXY1XSyu6dggvMr8nuS7xFKjj/rQie
/Pm/VFwX7fUj3A2OfCZ0PO8mTic6hNSOnnKyn4cNaVJFohnpyDN49N/tOP/7QrQZ
EJzppFpGFk0SzcGzwlFkX0RjLbefxeudhG176H8dGv7qLO66Y6+N8dJyCYIJ74om
RYlzJws2wk4+Q0y4uevYdIx0wQ/ZQeNT9CwfKf9v8pHQvO+tusoc83HHJQo4kaQp
FXlmQyncvKdq5KqXkeoRG2YP6ELkB2svDKyXXdOKSbVuUTZDtborSImgow3N3uaF
inP2au5JooyiJsWOparN94I/s96IG2YGg+G04zaRKWzPN8X3iPJvZ5TlfKiVYAg6
uZRGz8GWnKxHGNJB61Gfg1Kz4hjDU9QRRRzqJMGNRAsmbb7CF0HIUeNkbWwGE2Yb
nXSrMS1sx8XFzG0nQeYMvEqMPFyKYvrO0hnIdfaiz+CNGkgJONYpgajJTFcHKy7t
uza73qY3lty2Ur+548N0aCiYc+ZRsrt8FmLcqXhFNKUyifR5Enc4eWjgoNW8455B
Ykz24LOhwx7UzEmm+X89Y+YoyNBX/jWn5Z2DhcV3KdmhRSch0czhb2vCz8oWOtl4
xRRHpYFH/9nteWCRQXyvA84XoqXVctaR2Am8ArPXDoO5w0gHke4Omqg7K2fQb9yp
koVEwNfDH5wDewvyQ/X0IcDAOpJA3KeVjVHtcKiBnE1wym7puj0oTE0x3oXAd1VB
EIItWoUt0VR+9xf4TcHZ1n4IvJv/CqhqpmzYVF3x7muhqndroCpIV7ymOl7ebMFK
yCcmpMxhU6wjwCEa7rh9EmvEjW1qREkdRCgeo+NsjPGOwtz/G7Z7iGNbSzSoqbLM
mREQ8x01nG0KAu+v0IeQnhSTqWphTtGXqqVCyAt2eDA/wR/YHdocEiHDoBjGN5cc
etPn09+Y1Po5ZpMdwzJVoFOHiefvxvb2E0atGBGV822m4l5ROJXkxxUhAxf5Zw2T
4SmU0TAiZWN2KeXY+fXnRT3bQdOTtKPsFd30D/BbOxSnPw0Wk9yS8C4M8uiHF39r
5gh0WxOKW9tSA3kPkIHvAXRkPSQLNMuEhAY+v9c0N36e9WQp6mjfs/ELNj2m/ZLr
Qi9O1AliH+afy75IlXg39itQrXVk80PmbOswVuNN1nagOCQqi5pqow8a/RPbArWq
YDU9VyCUmpb3N5MTliwczpAjoGOg+Ir6WyM0r0rslGyU85sMZ3i/21ERvUeBIcij
tBPvHCCXeInNmkUY3nZnr4Soo3mcKew6q1htKl7vs8264SKwRrG5sdOy2nyQ33JK
1E9DUcbfoS/++0Flvc7xgeyy1qH589VEaDevFl+C4jLoyeOgQXU2dMzAvpOHFcfe
3BbpgoYM31TBt/2Jbgvw9f7XYo/YTQz3xKSYPy6a/IwoxgIWzOqE9N01qctyM/pa
X6Li3HHaQyO6mwKIgOwfX3uUl4DqQxw8HJwMioDiQHmXsT2MZJKOLQCVq1IVQnzu
mCx+qKk/vUJvICnWkvQ6jM9CpRg1GZ3uOByLu3V52b7elggzrCPAlRciEdl5tIvU
X4nP5MsLS7lXhphxMZiubg5qlT5TQ+5bUG0bCoAQRB7oXELAbrOI76RbOlSm4MxZ
P9l/BIjk8F0CqPhcaW3n3wcSE9DwMXn6alk8HeNbk9kGzVt6vtwNg2jZqnbtfmgn
75xGwUIoQR9pjwLOZINoE0fqiFUBsQlBP0ajGXbGt73TJmk9bFA0OZQ7Z6q7F7NI
uw1O++9bCfO6brUORYpbVGaVHtX9sp8B/g0xrbzbn2HMqEQ5jAZUOS+9X6OhqSff
nFHEFOYklanBzUH+Ynklkb6aypYX9aXt8goUHBItv5yzLqPTIaHahtfqkEKrsYfE
0GGxPSML2R8XMzWvUKVmJwRqi1L9gt0pV1DDwo/YS8DT/ZKTbg1mRu0m3UKxqi7n
ZMFU2nrAkfZHMo/BbiIA7DTn0L3UsIuUJw6BYzDAqDxte/tS0mIuUD3tSHyHlcoO
SbyinZMo/KDQEP5ewnf/kQ5S/aydK05tKC/L8z0JNbzavrgBxG4MMzkO/LwsfWf3
YJEoDDC5iSmlTtTAqig7rUdt5qGsFKVrGMcPvAGgDp9YMglqp91w0Ti1fftQJKnI
/qWECLb7b7NKrmb3P+2ldhxuNRIKvTmmu/6EEGjj/ozRpPURvZ7SUhe3xTqXuUZl
pciMauR4ZXrPyYhY1wR1FlOpO3SEba2l6baWDz6RLL1ZzUwgPJs8dO65IyfBpbIM
7YvZRg5fAmdC1xboPD4ikmLL39b4BQE9I49Idj+Gm9gVGg/6IzCf2Wc07rmBd1M6
vWcK28NCn5C+uLFAQQgCY6inJs1bAeKFiC8X/Ii6YAm71iGhzhncpZJWElcsUmGI
QriCDOBqPoVKPanN1Uw4AZJGTwvqi8iloooLbxSPauLRWLR0asvk+nqnTT0kSp/6
rDkKoNreqHLBZYwP6uqlCuluBTixuw4rBFcqfQYO3Eo6lIw9JWN5QSCVJfZXEJvv
rEbh44+Dzboc45GXA5Ann46uZ+QQLTgF6R+XW9a7ulsykHBLebDSVOA7aIVdIcf1
oMCWTNv1uA22eZqb2MGon0BEhHvb+dg1gfNaRiSHBoHJGrTfkgPyA65xuqD5EDzf
QVMXhkhymNMVDAu4lNgSO9gxENLPKsQj+PDtr+r8GIFtBUogFsdlehBllnvs2mLy
vw/TeK0TjST92KY4EvW/l+nfWFx+qKhCBo6QNj5uDoRWHlhXFKO2cSjT6/HsuROw
S5i8s4yaZsvXq40udNZRppocI2H6FrCxyka+I1E5G/+HoLps6YufN70Q2JOkqP3k
zNmlH/HtWbxOzg8HyYjz0TzpqA1/pdnV9VMSuzXsigrSbXmbyp1y+Ik/RsbzwFJ3
Ov3OW6sF7i3K6alTS6SPcUYPf5FyEP8YY01QjBCH0TTgPp6ajQh/fTXizgJFrKVM
17DdLpYw+dPWuVSdWFkrl2LXC4HzCEYb+uv25NbDyPu2zDVcspu1Ut0SbEFGaFb/
spyAnXRsSj0DINDVp3CG0rtLhjZWJcKVLNJorZqRNv9wPwAyeHC7ydsas0oVLD1m
A0aFWAeePmMn7WCYjRHrti+JCV/8oY/uSEWvcOW6cYEs2u25X5aRe74XZ5BLjxzO
v/p8o2qLg/a2pyeZDJM2DGIrxUxox+LyU949aw2k7gkGC49rOxtwsFRzAu7fTKUq
JfYn2gOUZBcBIw/Y2UdeT+WOKVqMDYAjqMCFUB9cKFbxjv8GmL986i6UN8FjKHVd
GPtIEEI4Ivdw76f1n3NLdKqdEeyUG2zeZHmH5wyZC3nud5BORTk01hcx1/p6w17o
8EZnE24rJrbIu//6GCBS0ocBxyeJPwvXL6Ay659oYAYsUk8MmUko8FRUiKScRG5y
rqBkJGi9A6AQs4tjB5ELe2x6rWFbtosmbU9wdQZW4xMsDganPTTthnvuOL/ODCQI
EuBEjWb+6Axi5mYbBsAJ61gIHohpUvibQFAvKgoMX5MHEKx6jAQkfwTuPTqyelUt
7+Kjt71zfZgB6NGcIInF00+CgPKywx6GELFcyS8963ZI+amHZK1GA6H2cUhD7vV/
5ZL6mOqWzDLP5NOv3Uuym86fkWH6j9u6nr8NZRN+AlZucccuI+K5bcPafKgXKXVi
noeuwCgyOSle4CxoyakmU0iAbdgsrEmAj+LNQtttrM/emKDv80hFGCP9GU0uSTte
MZdt8Mwcv7H0v2zfKAZnbI4kKb/zp6LhMWEHBdyIMiDpHVVyNY+c++vEGmaHZLds
NqTtf88wmbMwx+TInv8O2zl8U/7znjHK7E+mYOB16zMrAJC7liiVYZ0fzN5C2PTE
ngyb/vQbaqd0fuRsZrnoT6aMsH9b5XpvnlRVDCpjO8PgYQHMNFpT+J938H7IivdU
Tsf5sPDEkkwZ/ZZ08/NwE7VgwpBh/dcAZhT3hP1r9RHpg6E5C9FvhUaxp0ESMIVG
bnkEp27C7bDy4LicOE14nr9QNSrDuMmwHTV2ztOzcbS0mZ1je4ALcNam2F34VvxS
0PWP6lXLS3kVISC64/rloXM1v7jUjZn08EFcS0OVEX/h5RsBsnj/YGRCdF4fjZBT
RbJRULR0Pm5T+bd0jgU342IWbHsJu0+OwHZZ9ZdI/L3yBoW+ZGevlxAHJV2uJjSq
4qFj8CCsJJK+oslPElT1sJx0OkzseWNN475mBcCnaioLKTW4ScLSUm++UcMYeSFO
+CHrHps90gtob9qNNu+F896+wLqI9ssYC5vic6oQya4O+pQnIOEz6Jl8Z0aIHd9R
QXPtD0AY2+k35cFJaCEjHIrjidcUmttTIQBBNkKdPKiaAUOJ9X2dqR4njPfocl8a
EqfucYXafys3zQDJ3CdVhGVV/ZfAXFv475WpVc0esjlVGHrxsCdZN5uwYg3KO88B
QHjfH5354169BCFZqEjeE6SnbuFZXZ6lQe77RQATMZaf0n8OT2oCv32+O6NVB5Or
0y7Db1aFa293xe+sW9nIPrRHDobaMUYadjE8mtJJGlF7ohHkGgwRhv0Mr9QN9+GR
NkRuYdxrhuUj3He/C6LP2Ww93rCaoVT+px2L/dOeg8QSC+YLwqI9kq/br1pXmS96
N4EcsicRnyyH364m8CZBd85a1dfpGTGXieBeUuuN4BKkxnjd/PogT4VizJSP9uid
1IcYzJLscdVfTwrdjRhH+244FLV5BZvMdgbcAjpgNFTyspxtf1mrkIHR6bmqE95b
ILb/ky/aQL/hDZQqculpEMyYkL+KGSnxOUI0SaWq3IVDyongQLU4GnCYNd+/MIVY
phWGXDNiB5MYI3kqRnfqfmdYdz1r4VwdCEO6f5xoj86vW0sxiYStHCOizGtxiXCB
tHfMKIFbJ2DPw/dH9JSxFluJztBw6jdKgdAWYYdaTU4ho2S5eGb3Ea67HldHDYXa
EWkigvDn03Z/dgwezejV2w/kofybo5Qf5mrNLEnxE9/uMcUtSv9hh7fjq20tApuU
dgNeM1ukvtR8bLvxCXYQNJECD9G8UqoTadibGNYX9qm1mHO4PvXrlDr3s7eTvFwH
eKE7o0JBrDQvUDuVP/GoEyttvkmJpDpuaHkmwO1/Zs0SohNZSrmKXQywpkgEljwf
VXSSrpGjkRWJu5qlIs0a7JAsURM32l4mADITezUYomPR5D1637p02nlL5LVi6yQw
6ZeRWNdRja8LbqEXpnAlfZ83UhGfqH9xj+j+ZZVQ+7MB3FJhmLv4jfq7Am0998C7
WW5wdh8MWa1NGHtfwnrOZQ45BYNzyQi86vxx/RRoFZdhfVj0HkzuapQDuwlHjObu
t4hNaN3vNM/pz6eQgUuBOHuZyY1xk0ZrNw9cKuCB7s91flKnI26PPAKBSWz0NQWH
Whb3rTSmObvOBuqfeqceywPEIwPKpVbo9p+zk6cJOZn4iq82Z1Fx2IGp4djhVE7o
5kET+MtlgMudZv+7c0PzF9jrqMONXBddY76vKlKU5fC1+N7r0QTmFI0861IuXj+o
iqUYyZBes1plydCy8xlFTADxsxlYAe7yyb0I70Kb8m1WogCCWABAoAVY3Egu3gIj
/H7zT0608YzJqv/RxIewk0z+nUsLtd8+BwFSFTq8WREMbSHTSLPwA1Aewhc6O8iZ
2p1u/va2mu7pdJd6QrxJVxVI4JyWaPS67tiIa+hTbVUAA3H6RUIiIZpqJ01qGACK
2WLoXYYkFyhhOZGvTHyajl879VtKFx9QjMHB/0ycR7mJa08I0pax0sb4jNNf05TX
WFqYQWVEmAQmEIIOJOuhXs3nlfOJgS+soWmwlHjhp+KzCHxizx8VSO+LJG/kyGm7
CmI0dlYbw1DQxqx0UGp17sNo4rp4F+bd3lfwmLLNMQCLeEpvt78A4v6OKITwMxR3
pK0W8t8xEZXFzgTznIkhLiXyKx73kGjQ3ka6oos295Ezz4kMlNjSicO6TOLhsixV
CirSss8D2raDB20ocUJqViJLoqXzPk7qahQcSi0TKSGYgQn7hFm8i8IKoA95V+ky
65yqDQswCmyfWwDatTrBk/+vdO5S8xY3xHiLYdfojEts+FCIqZyKc921texc0RCH
5hcNxEu2iwXe9fVe328f8im09RgFWHEZqxKg7I05P5P3xbBkyWLRWUoYs5SLF/Px
VgQHlM0PL/Vkden5HAGvrXJYXcdnlsZIdGPhSRcI7CGKav+KSrbZT9tDwZCqIM24
sdjxQI8d37O2Ay/iiCqBjedIR2p0jjSdTkUTtVEeICgD5qag/TZ/zIWGn5kNLhYX
Bt8MVeEJOSqQ2bjCHUxPsy0INJMnNjD3YDiSYocPZG3fRkTovsQG0GgK4ieiZ97c
pPEOlDuC2FIrIicO6zHh12yzauUZLg3v4RJTj7LX4rVN3e5iIZdQ48iQQBNDa8tX
vdBdaVj8CUrLmHV1EYqqdmhI8Y0bZX2C7WURtDN1xNYqm2sm6gtJr1M30VKg33WL
uswQJPZkJ8Ff2K7o/yJrJuDSZ8n4rq7rw1BM55j4dt8PeJd+AmdHftLOWJ0M+uC6
6KPrPShFA8gkN3/aovcsA1hevxJVx3tEH+lnhsvSgMDSdhFZMH7qu7YfvMTmqmAa
1RgmGbLy+5cAvAXZVV99X4Agf8UWvKo8VXOJ6Tzbr+IhVHyk60+5silrUuii/2AD
MYUvPsEWKhsmF/PMihqsTHr7e9cgQZq0mvI939koRYZlf5AfncsRrpt2qS3N44Tz
Ed8r9SB4E5CL7iMZbSqrneB5JfOIbAbEY3fmRVN6uEhW4UAbR8Gh5CSwymEwj3Xo
NJp1iLSoOFp6eBtRbOCSWtgev/CkWhbmUU3tYD0sq3BC2Hn2lnL8q+4JfkzCASax
Rq/iftf5eGwbU8hns+S0zDnT29iIrYF3Skyccm3uCSHSSLUpFdtRvQxRcn4HRfhP
dY7Cdfz0k6f/0TvuRmS+si1ab31yNi6VB5eYWTO9G/0CUyYAkzelDkz8doiiBDOt
han/kGnGbengim697F9w53HM/xp/SGR/Nk8OEn7YIW3FjmOKPklgrcDzPsMnXbkE
Fd1T4B91QhBOQqQ7Taq1cJ2svbCjB6mdxVwRUf1+h7guc+ECZ+jo40PVXSsPfpF5
d9YKP4fhREAyFL6AVM3Mx/WhNhcmSqpmCtrRUXEKvdMKMZ1Vw5faD/uMkghVrC+Z
3/zv0bKGckdvjiAGHb7g1bjtoo6XiTAgWrYodNkWBSdAZyj+DreUjcQh7LbuGQZx
+FbQeI0cu8F1/Gm37A+/dWOybwfDE3GpftA2N95GbJHlTXpOB17Omkh2QTt88iR9
QRnINmi/82Sac8JHbafzvi/QEFd7dS0chL06W4Yn2h5zORwAzCFEKjcDxhN/fdlq
c6865oyYaAlgaLvleYBro5p3NFhNJ2ufYX8h9sUQ23Uc50loSYj+UnAbN89TAFr9
jyNQuJBHUJTPFG+/ogW26uAq30sN3u2zZXUyet4BQvRHDzDBu/Wc3Qtu67JDwwDG
Kw+8/RxP+vh2ccPohiIXHzpfA8A5nh630pyRyFdPH+wlcGjaqp/7XAXwiYqiALja
9LfwM6MjLGLY970UdTbdkfnOV2r0EPETro0jyYNPJ9O5oNi8de30+OJW7UdFsbzb
3C1K2oJ4nrkewjHJM/h4XurIN1cSNzPAZkGn1WMfCKxpJktn1zjBivs97OQUArRf
FbLtG56cbvMp3h6hpqZajndVe/mkD4PQ1L9aNRQHqaEqPlT807hPD9sAHPq38u30
6n4qooQGvpjhsDhY6vgFnJXTMbywL4ckhRG1MpefXWWcYoKcLu0aYh+DT5EQL8SV
BVk5cj+0U2fLuD6LfOoCfMCbsaeNtIOPdUy5HB9VwCIasikcrI457jVcIRkwnU72
DIn3LiE/N9ebgHEOjy+T9QER9uAAmVU1VYzujToUmS8c45PgtFh8+24M21Yorq/U
0Wyh8zrOV56iCBzbmn/HQkCDYiHLU+W9lhAfi2X3foeqCB+qhtDrIf/sK1nQ8bcb
V4cdT9pZ1Iwu4ljuXTKUsL6VqxAp2LMjHaS5/l5RkR0u1R1+DwE4V0kh1/3iayKB
czsl9WbPE56TGBqQiwfJIKokSefbWoapIfHIcm+tGia6x6Q6YXqM001C6Alq8Ua3
47ecFaamQzJkTQ7zns5aX3VZG0FGmfyugJVepgXxuBWhB2ml7Psl9w+4hFhXSESJ
lGiXUoXrFvyWx1EgMwV7mWidZvS5+Ixksar8v8at0Khq8hxO5is9qgSiARfEJm7b
+ta8DjXA+/FwGzVtYcY4VAuM9COkEgCaUHIzzROPbutBvK3g3dp6VE3SLzEKtvpF
vXmdZyWBFT2s0CJDrtuj3MOwovIosQTnlrYDiYIVEcugskQrmoim+JVl+P2boVHi
m2o/DQnORnA+oaMA06esvCfqjtz5mpSbsQpmTF0AktL3aWOikc+UdVZ9s6u7rwwi
h7/cuTRa3J6qGAJ4nnbeI/z9kGx+/A5bF0uBznrEW27DXUrk1tYEnwa4GuH7t4WY
3lnzyptGkooM+jl3Bq+sgqCmXBz2/XGDdyJjq/jGVUKAuAlVDQzkynVvhmUA7O6F
VCXwWuPLWnnRdLgx3eEHCvUiJEMZGnJJk0ogpKoJEdf65oKmNc/djkj0LKPoeP9f
+WncdxqG+jJR0bA/6YiXHZ//SOy4vy78vHZC6lzp3dFUx8Wmo3K0D1t7tXJIBFid
6aliVfk0+0Pt6yV34y/HRVmJsq6KGtiIiFEt3I3uCJWeEU33cvujMk2W0Awd4gxX
6unK5ouWyJ1srl5JxI5qMGQKVQe9A1EgUuytYFAYQwIS3p3yDiV3YU9NoutoSdK8
T552csx8Y6lyTuvV76x7wIEaEKvh094mPL+jrBbr2sMF0P/1AP8GfWbuBKtLs6CN
f9o0+TlwJEvAwt3GniWTL/ahwIa4/cx2zCNmQtCTwc9cwdZM3y40KTsTznKd9y8+
ePBFlU5pjkx1DPXZIjypF3PAMOS7MzRp81SVGTy/gZ82e0KuKKLSnGSbHzzeV8SM
modvYVIIj4ayQbSGW3Czi84O0GR8Wcg00zxAsyxETNfPV+6gjss21oBQeMRWB9Xp
/+cwzJmXKqQgzGJhTbrY3dFVTzgO9kHxTmPCxpDdyJLxagut/q5e+gKO+JRcyUn/
2LOQAdl0AtqZl5kuM0au34BI2dZTJN/xdH5mLgKpj42V6WCXcytFwZ25+a9VlK2s
kQWu5ZbI4XLGmmqdhoG8h027NKX7gSnR1Vf0pNVJqwlggQSI2ZMiqLu0bmrCU9+8
w/jNy0ZZjSBuiskSm+nHH96JazpdsniJMAYrK7+45KUv7FoMIr4TjzaUbFMoSflH
UwY6LAs9U3NIh/XwkNG5wMab4Qt9vtW1JkivYMLqCcx6fV9m4oMJRfcvZzU/edO/
eAEo1Uv8dWZAut+aCHa8yXOio0uZ40pF4VQl72KOUUIYNG8uSjdYPC0vmYZeL5tW
07yZQobEBIsy6O8VHv49Na4Ni3Qa+MnlcfS6Gvy43qWcmUoYrKVnP5s/qfFFBBbI
iR0N1yh83yZwQ9COTZC8zXoh3VeA90zlYrlrz/LlORKpbPFLAQAfVvwDiX4GrBQI
BMQVFM739vxbSAK8nHLEzAGSoK3OAe3svsL2ih54a3VtWzx4PA/u531QmIZq6wSX
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5rGR+vaArvR601eF5DJKQd8YvR2uMy76fSf9noIw6e1G2PN7BknDP/o9tkn0sao
S1SX9EDMVkF+W2jKEsGn/Wlkpvi6M65mkijshOGe/0cMtF3lpknrHoMJxTWChkf+
RJm27xYizzsWdjnzxLBdVYsJY14ILDYiLWyn3KzMRCI91Ht8C2Y8wmGsyxUEFCAk
A8+5zsr3DircOF5cHD7oCVgZE/T8Yk8YnT2jhFq7v124qSaa8pwbL/CUXgl0aVTu
1fg0aW7Xg9iY9pzSYeNEBgMmX3BVUbNE7qgpTkwtBetIT3wbigX3+GJIrM0BIu/J
7ScMZxVtbSVAfBJA4EW/4NjtGFdOxUzoyyqzeMNFg5R2Yj7/4HRsoU63oA4pBPTu
kY+YYHlKuwkI3MaKXAg0ZYIAv/nXYH1FqGqvc0C7czVSefXAzw+VQYLkIYEKUz/A
zYCzca/H3gpdFimMctHXGWrIIcjhuB1fORCglUoXTzeaghtHlbOanD8n4dkq0aJ9
oX9zu44ihbDhtbVvdmbkIeONuSOIBNE0w/ntyhcIg/64wWK785q9WGjDUfkp1LZe
4ycCM2G0rucH9gW7LOEiiGPZU2zz0TH7vmNAoQEUYSuUf5ycZdj7ap7rOWPCiLY2
3+/gQGGMvjabWULP034+3ku5KHKWULn7qbm/kFXPoYTPWq4cUTMbC8zhm+06Hfsl
WXyFQgVDmBOvdv3foT+XpXWSk5y8GRInwN1lt1kpScdDL3Av1gNeAFK7SlQ9hOl1
RmEE6+srCNmcgCWy9fWG41J6mf0/6UG4Vy69zMe4psigof6uaHf6GonXNRupV7BA
49Bn5PPmtBJfcfjAv94CIuWbiEURwcjacvILSDZRKv7LuADBACriRxMvRiBCGFVb
K/60/QLz0Uc65QulkrzCsc9JbuxZhEXoXHqGhS4IQNHK79w8pBwoZ3cW5Pab1MnK
kW2absDwLOCjb4esHC7TBDSgUY2Ll4VIZcTZjhWBV/LrM2YP4t+NNCl6XLNBFEez
/QC7GI2TMz06l5GhkeUSDMuERvBqgNQqYI9SOt7yENgpTUzRJxRomSpUudwLnuaU
yRf/4ftqTDK+S0ocswYPHsqmGHltUB1ohreVsxrFNR1JXwHLvHM4OJYgpfm1Gpze
zdP8mLh+mo8Y3I8E6ZsKk7cXDiWO2QBUyiGzigrx+8oeXRbi7nwsIcJvW79hUxgc
DQfGhEVW+W5np5pN9EUs1zc+dGTGLBfGVZO6t86jJ2kQHhSQ9S4aOIyFSR5F764S
jZGAEh8nX0D4rLwSs1Zz3v1tLbX0bbYhKFslWGZ0/b1jLoDRakQPV0Sv9zZ0dZZH
bpVmhUedAaDJMz8XOT5K79tdsyt47nHB2uQOOJzcDmFpxPbP3GXA+w6Wkyfddpnb
sRU/YTQlzdRGIPYBzBcDGuWpk4YDnnnPCV7BwJ1yOt5wJrnTd65RzelPh3+GYEbF
KE/tddU75h8RfwXDdxJZ2UlGUTNvH7z60zzbbDtSbc3e0vU5jIL3/BU+pggcCV4T
5Yfbx/mrynzndobOCt5g9M9Ix98Itz4RD64dJ9w7JHT32/oKnERPFV6YCw0i1+/X
/BabkDKjYfqfp86dhm3HFEh4LjtzxR7iQWJyrkafEAm/Jow4Vm8rWsQ8WVmSZ0KT
yC3pNiS1vjsngU9vfnkT3nYAYBsRUwjlMGBPm3ea0YG/u2EHtJNeUWRd7UtFy7UD
f13zbZjQulgWvRQYIy8XVBUfX6INyCnZwb2iE3X7PINQHeG7EFk5aShUlh64ZXjo
sIYgqzmDCeCZI8ZlzszMYsTgxKmSAi7sEn13RkkrIhkNtcqKQ03ec3L6L6IynjoT
oCPwa9NBGMmRnGCFT1DyD2Mlz+ycIz91IZvWePdhQM2lj2l/6YQMtC26uLIfDGhV
A/P+2h40zSO+KCxvvlChYZREhV4DCrZGtV79kn9Nv7VBUPsQqhNb8fUpm7CEZd0y
QnD7CI/f5fpWhQx7yfbN+bX77U6VT5rlsB1ktmlVruYm7umoICvHutWcbmE48xc9
+9fCo2OxC1MYfXooQCP8HCw3pU7/4G2fb55SDHGs4cJFPaD13eMyhaVSFEahrvDJ
Pyj0+Pvp2R6ktDYu5gr4NyPkIzzeSsRWQ43SeKM+/oph5HqLErU/CojNcGvH/7dE
It1q1Gq9ybCPaZQGtXJOhsSQWdhMTrrtrZchDdeTxynbHWwVUk0K1f5aDWyZT7uk
OaRnBIySqKif58EUhkmdN/tsEfVGcFm8bEQASAspIWAzWLPJ9ET8S+BbMeYRaCnm
yx4U3wSJzXVUxo/eLZ1g3D3Ts8pXu0T50z4aQW8W5e0qiTNXo9m/zH9+Yq95T8lO
+ndIRY6JtwSh5tcLGPZmOWXu8N7UcdVvYHm2pc4Hl8yZmCdgwypgI1uMLZGXhzj2
d5bm8xQWI2S18EuvaigqejPyUTqldQEGrDQaeJRTSnjNo+jD3OCJDmqoN68qvw+S
nM+cNXGrNk9yzfKSVeIW476i5u9VP43S+iTV3r3kxXMKXqouyawSlhbzezKv8gDB
pQQCrLXlEP6hMj8q4B180uFg/z0/m4Vsz8jftFVyhgIcijSNNtf9O9mhEten+7i0
ezYmtIA1f21zzHEWkieYphYvamCnc0J3/kIn22PaxGIhEG9UWAF9tnoXWO3VpjAb
Y31G3UJztrlBTMlIQX3BTwdYhcKLhaejv8uNYioFxhtZ7Zk2kW14rpqC8zBWoVHC
GYU00FhnD6U7snk33kXxAVQr3zc8s1UFeHkQZJCM2KxOXARQ0qesz31nnQnahzgL
H5lIYtpnJOHBbYR24KnCrinFRD/maDKukKx84EXjioWEM2lO+H9gEkP6GDkjjE5c
zTIBs40UiF3QtpkK+wVyT8tOc/JyWjF+BQn3QFQq4KpLSbgiM5mqLFLhbItUvSvp
zoaXc1+tyvbyTKXVVhEr2sDn8387/Q/x3KB+y22JvUoibfD1nAAbZkL4g3euqUtR
b8vcpWRrkRFKCjPH3uNLvZGWZYTGxykV2/q6tkqRHB2gTpxs8ePSSDF6h1Vt71c6
t02pb5YxfO37oCFJUQzkZJgV2NE22NORT/kNLn4CDq3/rwIuwSK1KqyqPC48FQb1
KGKocYMh2FRy1bMaMTbdAv2LJce6vw6XBgjBr9Wke2iHGwBDvAYJgVuPvm+WsU6M
I4lQjF3W1+IzzGWhtY2a/JA3KTNxSDeUsEG/34IWwjJHGpXpngORo7Q1J1A0e7A4
EHdS/qeRwy4qfC4n2eY6F2+2aabX+A7XzVX5FEoiWpW3UPEHIP0LWpXGJCs9hiiy
KkI7xyntGbJ6IB+47t90RVkTBan4zY/I5e8DKuiOSnb4GZX5cRdZzaLPzdVfKUD1
7qqlW7OlWvw6wSOUrFTLFeAkMNIRa8PBrAo2fwAaq/2tx+Juq9lx4SCwe3QaByro
IS5tA2zNhtYnT2eTPjQ+fD4i9l0eLZVJdDuTPUKikkRvAGMp0yjTuChda98orf+G
TySv0FM4fcdUP1znjAc2TpSAfBPCiF1vmiVsVxR/ozQBlFPt1SEwaTUOtLnTAKu4
LEpNi0tx+B3FycDeYkqdRlXfqcRXCHWMBy5BML50xDZBuav0jk7h+3kL8AOXxzbF
nmEzU9NDxsP1APJFFI36krJN9xWrqDk0B7kPOca0HdxAL7BiiYBSPb1G/Hzu0FPs
vyAWRiV8aF5Om2C/x5iiZvl1fo02IIWao6eyl1QZ7hCS/cGSRzneTiBIq36GwN3n
4HO0pRZcWqaiOAMAeJhtNgofpzPlOBIT+6ZO294FEqIuoOlg3i1LXCxJrTryhp3m
WOm8K8e25L+UskOL9GFn2RbsbmnMd9J/QTeA34NoRKZxImhQxTtXY5/L58GarNwO
tfP5GfDCR1+zDToYxv5/f5wKcoYU5r0D5lxGZUIQOMzsvRyLBP0qaOP0tZXOtZnQ
JJ+NbUU6GFaLsDR3x7Y4aFZ2zzrcmr9QGpYEwkX40keTkdufVlcpT+wJGmboWlnu
VIjFhQlodjJmdpvPORklYGKPyA1V2aqDysHnHNPN9Dt3nr6JQGV89Z82Fzck+Zrt
eGRtGI+ql7AxsZ9683ZOLS/b27Ck51p8PM0b/EglrCbzyGBWAFO8tc0CTW1YVuO2
lDlKAh8N1AvQ+zuuTc/kY8Jg1LAKvAle4qTaI87xQSMt93DHmqCcgrpOw7vbJPzP
cR7Ryszg/hq/ETs3GyEoLt/mXbKI6Ngt8oQseH6bEpDu0dClJUNSE+7vkRkv2DOY
sQ51s7FCqEpwttwjtMhpre+RcRIV+wW7ApZxK0lG73p5MWo8iHI6HlbbduKBABsz
8d20HmCFJ34dKu28PVZTbSHPMJIhrX+ga2p3qoei0DaowILFqw4jcr1y7ZtYWRNG
/ESlCG5fNRLUGcQ3A0baU9a6cC1yQ1VK4+C6w4oRMrTNNBhwWLE8FuWl9HSuca/7
Z71kf5cdKmhx/Ybm5hB0Q+oXwzKSv/fymVNH0rQVpyKpobsI0/wkPm0Gn91WzTVl
hfqiFOxPLmMfG1LD64rcoTQ3n7sJ9AJ/f8hpZI3gwgXH4gDV+6YVSNie7YzKG70t
o9pDKGWEp2mdNMMu+ILiwdfLfmTLyM4mDJ1IjK7fJOb0nlbvNvg71l4eWtbuea3N
2/4biUrfI3dUnYgRsBZf3NvV5opEAiiML5g3XvSXr+96jTfX1bAFJe+WKLvyK+V+
S2w8ztAzDY+IShKKrr080FktLf8YqKSVB5ColEYYqA3sB5PO9vBbdoS7jvjpjdjB
/3JQoz7OaR8vVhipapmohVmJNAJuQS4UeeFP/G2X+UTKZFZePjUIOGwsXg7Xhp1h
qnWh6um2jg6vm3W1+nrK5uxWLtdV/k/aXmfO9QMyMH0zTaEWIGvyGfoyFVdJ6GnT
6CZLRAp+EHX1pE++ryDybL65atdHk+Zw3LfvTgGpVnRcy7f6CSkuqWBjRXVT5l1L
6Z9HvIrj2l+J32y26rwdtyk+1aZpvlZBYWrK0HOuEy7RCnZYDq0rVveTtApBXl4U
W2SNw2ha4XpS0IUXLg/0DDxXNX3GbCvc0nQ6NNqCdwb8ryvvGoJXidg283JEuf+M
M6Q84dauM7yotVTLfY8npa6Xl01OIZTZyYqekg9cSByfdLqKD7DTjFkag6nQURPp
YdzEp70agkxS/l0qY/Y6J8jXHBmFq+ouJkNKT+zp9eu/5u5LK4+zH+honmumtCpY
3JXQkbH5U+7vuBdF0H+bZr+hCxbM1/uNGLs8sFxyb0M05vIgc4AdlAFr0pT0nsU0
axNia+SDlDwH4Le6eRbslcWJClGHVOYBvb4Yb6+7kSvssXNBvMxC4hY0ONSk5ypp
5dpPVWJE6Xsz1utaWYVzFUjRMJlByctv2mCM2vHZf9h99KAnPxwC3rl46zfi+HmF
WZ8I0Ygr2Rv2PpqS5fEz4AEU8xFtJwzEPfqlk16S5J6WTOXoZiCj+pE1N+SFv4nH
tddnrCDI5iuTvZ/WZ3Jvi9VPK75/AjoMCtuJ8f5lSrg7MqIJalhWJ8lnUS4KryEU
LcFxC76x0M0tXxWFFozGjSc1n9p/D4cwZcfbGpgFxV4gx9dccyXUAwpRu7qVU5ZP
3kIYl4HNLGScUcX2ahi/su4ye61Wx1EqXuqgjFYuVEl2Cbg9RV8ABe6tsAkMSxpa
HmWk0n2pGG/gTgwvW1AgksTRXFejbZ3yYF8Py0RQ7+t67FbJZFQZEfer+hozn3mR
ECE6LLBLQUufxDKvczaJRnwhRAPu2lLR4fEPLR7UTF7BvXywBQRop3jCvLuCarNt
V3fh7acM8c1hqt1PDnfRk/goCa60NUVaisw5pivVRkkXe9oAVfwj+/zsnTfE+QNj
qUfdsUccy0V1gzVkWutzAKqhytqRDBfcf3gZmpJEZHwHp8hmBElTLXnMeDyi4CEd
PB2XJx1D3Ac3cNq1crc6GVMp8fSXhBSZK0+VhSfLi75G/OqEBo2C1cs/2uWo2ETQ
T4hmp1owkBwmyDu/g31/bBdFAiXOPpbaLzOVYYwrWTpg6UnE3GQbj+FaqST7riwE
oyNOvmIXlS5MLh9LWhOgfN938z02QJpB8rucGE9fUYRosE9whOMkwHiL7iFQQCXF
EljdrhVDU9041UPpAeZHLanEKfZZ+l8sgqJxdlIy7ieZgvMWtA8tY34/658PL0B0
HSb3eK2O3klwouRIgWd4zizk+mH/ag+Tuu+wNMsADKvEweLTubblG9OOSypsttGT
CZ76dAttKRsi/bHBtbVgp/GkjhHdhK+9tCIb4C18FlLYtljC/PAIH8f894AxOzJa
UsjUDlemVQCUQSsW+Ad7CNxX97PXtGgAT8crXkk4ZKMqAgxtlxFyVbjd3Q4OCsg/
lyTwzfdJKuV1OMeDhe/hgXudkPt4FZROYezhYdbDDHZxk6L8tGIbZFweXGdKkBPL
ryA/9kuSLyCUYowmJA3wYbifF4BC2EE/DyQj+ZLJ1CRyzTn+xxflXSOAhbWsezvb
4KfIqZ8c9mTjLK3W8qH6CLQUmKttBUguQk8pk3Hj6rW5pp4dS0cA5V+zWWVeoaVL
cJob2JRaIBAmh2BsFo2JuOmc8hoYlGPwBQ9UIU5XfGk0+SqczK0NFnKKe/i5gwUF
+JrR5KJuUZDAtVTK3RSHpQ7i7+nt8Hs73L0B/Tq9Rf14kWEefLzRF3AEJnqm5RgF
reVmlv49fUX7Tey9LIGXSBBWFOOcwkSm0MQRXK2UhhftDW+emB3Zn5fRjlfE7GZR
SzuEYWrAFkdpLFQ7mjpfNGNbx77oID79uaPtJSGKXXuq/K8uB0g8I8j3XLKTSNm5
b8fVpnl49yrRbj7KTwVqeeWrXaGNXYZrXmKvGG9tsK/uNrh+29y0NcYZW40SxC3N
4mFhy37UGbPZfIq+PRQ4WxKCtgplBxzL5OLphHM/0jI0dCvL5SOFT+s8Cx7Oqo0K
fzX8xr46afn7qZ7zIrcW0628WuoFdOfvL6I6XFT5OYKQamHJvtAu1foCBXbWuaFv
WqDUHF0J/SM0RmMItVYQMYgtgl7/hgY3hCK/KNTkQOknbmNFcLuSEi/oIcre9P4x
CDman+WN3ntnqFF0+lSiaT4y6r4Zj0Jq+V7Ir0AQTAs0X+JKdxC4UDDGjekFKd5L
VLD8RK5KVtKWw2oqPsfxfisaDoB8o3SKZ8+1q9cAaDLFnInSdivJyuuve2O+wsyI
NOGX56DnJ+39fsibFhmLCcpVkqs/CKYtkKl1ocD5GExSQnDkTZvkZ4oE6W65Cw9W
yvsmrPtUnh9XJy6hd3WWlliwdJWSkgBgbUBwlkl0b/KCJoR000NtauQyQnFV/ZRP
eUa2FJvbEJYDLjWNV8svgTd3SX8Xv4b0fyEgwFBU8jErXSP2Viq4KaK5O1LWC7Yv
4IkMVbnCLbei9NXV9AQtqhWeOsizi4+BPaiEeUXMbDeqlPrpUx5RhUMSzzZ68/1L
WNE16q9PwgeSUAHUPB0slLLr81Rvin+LDQh3M1kpcodGU+UGC2XHn3uToKEWBYku
P6LYcW7UvALzan1sRDJQhrz9UuOZmjhjXbKzaCe8SP78gOMkOUmgjJ0DjqZJhF7L
6XaZg7qC+KYb06vUYw73NblBiGj/OOGBzBReYuCwUxPtQJ6aNoxrIh9nidTfXovH
AzDrZuFSdi3S+cK/w0mtlaHfQuXLRA2KjYiMBDnd45ZyeYUtPGWbG/t/GDawEyrX
DLfts9DFzt56rql4q0gxS/4Aviw9zAMGYasvFrp86clt5Z/abRXFh2l/bxY7EnkC
60V6fcfMrbQB+cHCEd//89XiHextSaPu/YAZf3OBK+GmQrpzJbsoKtzx7JW/e5ZC
WvJEZzXPgVhDjLU7u5LRY5HRtDMB0Wfypl6UcsW1hsHGEcg9DPfbu+9qplvcRkK9
f/i1wBfmb3TIfDEJYXOLOW+VWim2W3nxJsWF+Ib6tyaRZWQpNIstP0GZr7qghU40
Kab5DZ5ZewRjZxoHMLjv/q9PETP5pt68RToVz6akobTiVw/5qtNlHI6R6PreRRU2
srH9+pfUWNpkD6BJ8oL5jc8BFg3OMq2pkcfnjWu9GqxLaS6FVlF+6hp225JWlFc0
M9Q5/KDMsJkfLkTb6o88tAw51Upi+esw5d8ofSN8GciHhjALOJciHepOSy9oVbLE
XPVJLZti4I1ME8aGERZvM0KQKzc8fHeL+xy3ULFDfITK1Xp3WJk+WT6Z/LfghukV
63DnbwDYqeUh1ZQ7JA41/hEuTAM0W36Si0sRLKO57CZv/kDPBOWh6BN0HY9nJzlH
3BaL1+mO9gZt5o06fLor/Rmn2QkVvAPbHu2myCCo0oXFSkkkSuZixB3RAPTpSCBO
MUWwhSfqiQFAoQMT9TiRXIG66nbotk0n9hegFnrsFWJ7v80SzOM2TJEddo1j3LJa
LPeZgm9QdiJYgydOSkh9A/3I+Z+JLmn9LPfed0aYuXxWYfUfIq6+kJjiLjbYU1Qb
AVoi+rKY3jghqKJCOMzXWZgGpagNFogng8iHEDLkljiK9nxYSv1W9P/3RMvD4UKt
QeRBGOpEOxcDwB4sS8hcnyyEt1sIlqy1jXuQKK5fkpbkNN52sHFn4mitFEC6MUsN
NQhfV1mZABpA78FjwmFgJmpY1AeeumK60+Bxv4DwHZYxcNf3hhbxjxtcdXVY3EpJ
w94hd5s13aCzcDNMP64LYlMxVPLvl05N4ZlLbG+uKjWMGjd5IpQObuI+5g2SjrQ6
8n/XXCNAhmA1p4sRJsGjPGLF7i54rrS+lRkHE766Gbsg3Rb1hwKwII0PZsO8TqcP
EUINhv9nkbUFYiYEq51mvoFlOmehMlarg971zxL104nIL7C36MH0I1gLBmdomZdf
johR1vW9CzhxvZBilTRnK2cVIrLKA4T6+124VqXoqYXWO8auXj7ZrNnq9RegWZzh
pTPoJYQ+gRLmVviAo2LqkmhSDrokUW2sJzE0L/cVfCArBq5nvdwC3XpkqEFJaFmL
3uVgNJ1oS+zCIMd4QlMJsAroy4PPpt+iSxlwZ0xx1+EUrA8tWbBfUNjs3oJ6pbLX
9fTFGEiozASKaMi/4oSLcRzmfnj7stJFsP3UhPI6OLnYBd/Mp8HLVIPR8sY76y/G
JnrpEIVQjf9dNhkJLDJ7K3Iii+dLRK+edwJFj5q8aymJeeLRVS7ba8TweKbYorZc
jgG0uWGXbhidr1P4tbp3mBOqe/gKz545fIuAq3miKBbGLJymKN0Gt6UEOAdEa5yn
oHxaVsYf+JgBhHQeTdvhddj8G24QQ01CF7QOhKjTfhFbSxQVrasMlmZaAuAY7ufY
HwUOooDi6TJQ6xDeVEBKz+NoW3f66XOa4GSTW2SuELQU0ADtaDfs6GKOAlIYqj5F
aoFb3Ukeb1T26z6y7djsP2DQDnteIHdaHp2StzFutw4GkBy5ZJ69tTCCD2w4QwP0
YFK4VHIc95B7JqBoheMeQ1n/pNVmGCCbSf5WUDH5B8VjcEQTdkGNo/Ic0WKeFIMm
WikRkTryxIZatjCVYVIphUnDiXZov1hBU6y4buXwkowXAjJqNLupNocLBG579FSi
SNgqgmTGrOv2qNIw95xF/y8AWcVLLyQElnGzieQrxHS6Mez6ReXxu9qxn2bNmbrO
`protect END_PROTECTED

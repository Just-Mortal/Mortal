`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4gE1JAo8fZ67YdmucL4DtDPQB6GjN44XutThSqdhknOch9HI5Dn/32na4yQiH/L
ot0cbR8BNxkqQc1+4EXwaLF+qfPZrm/+Tyw/k0FFajwufDbyJ2VaEPVpi04mrcBF
rIyqWF8GWBQWnb+XshAWjvZMTv6jNSnIjy0S/WMRLD6tPHeiViHbVupXBfeGSZrR
iyRCBDWhx5BxdvSYFCAB1p2ZI1JxCsQAWnvo4UmPz0ddRjswCxuMUpxsKy+Y+Kcc
1Z7W/ujEHiHOvC/qIr1m/q97DcQEKYdAGkcekHlzWEmm0CJzdE62ijO51N/jAPof
W1HR5YrlPppdWCFJqKND1Jkgboo5XfliiQdFY9NJ2g7kxx1Tu1rzJEB0XaKenGfF
/+BTWlu6dIprtuPMj0VTHulNQc0BtzZ0y/0oPFq0mls57CG+zMOzBihKLhwZ+k7U
Ju8/qfdjBd5C36Tc9YosPrknFtJlsjURHkdUc/ZYaz8a0N53G/TkR5jhS3p/I63h
/gyoPrrEdX/aFpvVvQXTFSxYP9IU9DCnnT8xgfksHWa1C9rb+ZO3D+s82YKJuzog
D7Zd5ADZcWATf13z/SSxwtxsVhZR67VT8nWJ0y+JhhNIWLCaPlNuQJwZbGz9uC46
INHXMf/IEi4YopPtWXGZ9K2FTsJsRwYcwV5TflIOvYfgKitSPd/D1Oj35R7SEQ8Y
J8zV8JknuP8Rsow418RREGKu48yGvSA6kQWiA6YiQFClRc5viAEiW+PqexBSyfoe
Qc1hNmLWv9nj1lXE3S+eNXK/hsgc+rPVwP1HjqgJQHrKsHZ5iRr5DCgeKApsNU/o
NvGSNUTWKjKbXhW4ySPnhmyUiRKJ34qV5H7vuoBNXpePE6oCr4cd/SfqtptzjArA
bIqRxBGG7KCbL43vlT6MrnnNb6BP4uA55pNNpYr3XDgL8ml4M1+NovxGsoIDs7A9
h0dKQLWWLO0rZX3I0nu+dpYzEN9NEsUYOaltdgSC8wW/hA9rcAirOSMIh+bz/Gan
jM8tjKecUAzrDUWk3Q86FyuTUvtD2ujNVRhIW8ROJDoqwjHl/SJ1TGe4cpwBthxO
Yak3hezS8gIUXGElPCdpauf2sE0FX0fw6PAGJA4OivRAITrDZqzd+XgcTwKuHetU
oLUMxiEHvhaV+V4o4ZswbRSHle3Bu7kkxR8GnjDDsxN6d26p/mzBf4jbHUMpFE1j
rl3t0/96F8sT8bKsG7YIDnBr7EiZNFDy0LwbZzLgTAD8PLbkAzUS7zCfSOZWUDV1
c+iifBly5SVW7AMyeWk+REwYhEh8156/bNn1Oc+BT0jhTjQbR1Xp2ZcujqP6I7OK
BjAv0enBoOEJ1DewvPBAN7VMtb5wT/gyuzhZ22kh9cL2pHMkhHLRnj0027aUBcAS
it6Yoz161qJv+etG+ZtmGXRfGTmweO7fv3+thXX8wwRVsqXJpMU85+4Zz3k7R9u3
qPOWKvi3NTc5x+t8qouk2SnzCgW9+Nxw/c9jvXt9sxOy63gDX+lFmIrLuXmBhSLv
Uh6T7/lYOEjPbx2vx+9EbsUtCtZw2OiT5oHezA0rK27yoX1WJCTwDLJjzKR6DNf2
YyyOPu4zLg3LEwKDzJVsg/0fnYfhdZq4hjbxGYRF1uA1m8CUCKI9pFrKGQd/bAp0
2NWhzO/9ihwt3bl5Z0s8q8efcdspcbqHbVloXZ6EQ/22ZpfIU1282nxxxVAMOtb2
mWULsPCLsrAnS5XygeBBJZFDypPYIhO0KlqfJkmnS7Mw9a203tmyBCfVcrhL4inK
tRqktvHCCSgWojHlBQVZiK+tWJkDCA6JUgijLEE5x+VpLAh/SF+34ZsAcIK5Y1Qj
Se+1h3t3ky7l+jx7uj/CLDCgkrC5wBwLiGX5uQECRhRwZcjPVPb2u6C7migSzs8w
kgWUniTQBfhUMJLj2O8r87KFCI2ncfIeMiMFFNySfnCauEXNLh+D+jItkv40/ZMl
/7zgE2ahRvPdEmMvIUB9+A+WaRxhU+1sn5JzCJOxwLDSKGi5gdj+tr/Vmbjnomhc
0NYuZNOG5AMmqWNM8lzd6gBmvC/udgKHz31VEONzUByhzQOhOhoKNJypjOmsO5dQ
12ckF1Q9DWDwlMaSM5Mkq1bz3vFCCzBHJaGtPSAYM/Ci2854LbSvh2BacEGSK7u+
inpEE1hGV2HR7M1mbAlw6uXJ2hUU2HC2TbFXyMbD9t33wqX4b0t0G3edFsysVRDh
sGMscZqLtP/n3SXO0xhBNvod34sEwAAYlXMznTomWIeAunVtwA71MYlnAdpVBzxa
yimFLVZBK1DMgO0PB/zE0uFTJMdfLUDAxNv28DQLPdCjV0NIeXkVtq1IbdAeUQz0
ibAR+mbKHs4W6jz+hTs0AdNx/QXHj6z+G9r5Z5f/EEsD5pSKzdW5MlolOkmR0ZvH
PkE7Qo8RQfYuam+kXe8cAXsPMSleTE7BMSB8vEHQxM8TS7UgizKYP+p/w6h7rcwm
rOY2gPNesq1b5POykWqmWStIFB6ZGv6t42VK30iOW4AQCn9p+UtfAmTFKHK+YN5r
SLYssKg+FdX9M7cLshq6t71CVPyBkg1wyhLaBKFmAzNgXEQt+uE18Cu34iczJcpM
0t6OkaEbKlZlyyd+flXF5VC3Nt+D/Z+T0iLSneS52ocEDOzltm85TcZBX1YTUv3V
duJ58hjJkFieQCLLlDCOouHcsPNiLbBXSUaUtETxB0G7T9e1TeIOjCkpF3UVHULA
1LLJK2qyFrjH48OuWscoc27Q5tduetfl/syQtGb091/i49c9mqSIndItwXFpz6xH
/rO9yOr1/ChokJxYU8Zc67nfzgRAc0rgpPY+6V85jVNAA+mJ7hEHRTdkYnAuupCZ
TI9D3PBibBNi3fSAqIoua8ro6PUd2xNp51zP7t2LALcMVPVQu+uF0e9S14J8Q2sf
NgjBCSgogJWBC7FkxgLb5Xquoc+xUagvslZV3/fp67ZqeHbHClU+nSsBiSXNTMMy
uG6jqBeL5GlPrnohVhDVUzVCY6EkdbHtlKx6pGmBNkJBLXvQARgM4Hqf4Qh37XCc
gLI0lKwYimnUByFznxxPIq83s+p/oMuwZt7ydZ7TCX+pH6AL89PIzCYKdMjFCXJe
8Bntes1B4PZQ6KDa08+f+r5nxFYCkkJlz8rFvM6vVOcEmOfySZBclZPDYFRHru+a
uErFlvCQNxjAiGZ6zyNTi3HrIvM7m+oEfXItXoM9UmrHItQywqExqKPu2tEbwhI4
/hYvg4Pn1C7/9FJ6rtrKkG7zn/nq7q1pUvixjoSXMl6n1+KKv7FLRnoWavE8e7XJ
kjgtakNf7/Xk0/tnC3HQvwOjBysB3wDIDCBYj367VuABpuDFotjHeMFFXhYjn+1E
oRJj1dEUC6pj0160hZeNHzkENNP+2zDVByk1BYO1Pdi0Z55By+g3so/t7rmRVX3Q
TJAp03dpISVNnPwu1ex0c7Mg0muNEBvqWcUJZ0LcS8jxRmgcCTNLIc2NFM3rUCAi
VwWdoLU2PyTAqBSvT1DceIqW1CZwZEjRyCMChdoqVUbr21+Ej5kTaxrqYzoCfY+n
aevXWyi6qphEgzzvbB8EHg00GUGiEYtoXKRbJFCYk9UYItMF8HU87HeDLs4e+HAw
dvGenAI8jpdSBAkGEGVHP2Jl77mi42g21PrOgrY1qOarUPEvByib975dV7dw3dIS
8KN3ps7X/pHplAGlYTlTc4pKiRPXDaeqyPWHGJ0zIBbANBow+1PSaYSZ8hStXNNG
CdS05jifNrk9F3IUtW0Rd945Dp2LVKhID93LVz2UXYjAUvYgkt5FBFmJsmD0wALz
M1GbQXNnIvvlZxynbltY/B+UeWK3/1JblxKs0yHp8j/kHSW0bAeFmBYZfYuzPFQQ
PtmK1iqtvROIfi07wiZIRJx3zdqJGqW7RfuKDvCRUcHInodpaTZmrjiSC7BMhzgM
TMXll1AXEqudcEMAFE2ST0dZh4hMe9Y4WRrhfME0r1zC0hmL+PU7u8oa/Ayi6Ofl
TK/S+dnLw736R97kJvwJO2JxKjlUMSPg4ojdBLSvnyy7djy9K3mj2GD8leLpQcaR
klzUOD+9jNd87cKyyJlGhES8avPCnzVM3dcOfy5Y7jdfVHAPvsXQIPjXkVp+aKWL
ow4ZmSxDQ52ov1BcEXPhOuKdlXlWg8gxWgcOExltKnapl7b1ZUVBeTtG09jMYyTl
bIDAdy8EzIVmiSRsxlhANeHw1wUo/4eMxdxpyxWzafT+kWFaUCpt+7ccExm64upJ
qn3meyPSERsnMwfYCU9IW3dmw4Lb3YBj8zMBzcFck5g3sHnk3kuMBp7ZS770Nwqn
oZILHdk9nZzwcqFjEYAmTaY/e7zb8M7gSHUa/yd/a64pT1POLF3G/ogFG1JO7kBn
INBQKFE5zrE/yL/O6eEJ5U6kKPsASKn80ngR5pEAOqTZ/D0R6Ge3ua8Pd/o0964q
jjPGQoJkA/Q5M9crR+mFw/lVRabcKXZ51LxC/5o0j6wLDsaLDrgGCYUWKTUvlVvn
5WX4pthVqDKpezAeiAYM4zlpOzi7P3I43W4pSlZKuWTE/f/CeunFKBlHO5OQKMEP
MXONd3iQyPcpfZAVAcv4DNAB65UuY1gSF/wgZVIPdJ/LEylggLZifVlaxo4jZ0Vy
DbPZ2rh5pv3LiVy1QTUglmpBX2nsZFNQuG4dmBL5Mko+ORikW7+EhSEXMEeyYsLn
TKgRwD8kmCtyy/YBmp2CkWyQOHGV65b1vPjvPoL7PRIVvLaYQ7qeOAZ6r8KkACiW
Lx2XRxGhVQzoq/Ff3h8Fw34dKtocdzfhUJ6ZlCHfAsZBqMbGwaSlZt0U5Bica6My
Da7somrEWg9tXWBs84kDG6pQAf+PYAzdgEsnRPK8kS+WP24UHHNp+RBr1TDuqP9y
5x0QZyrwQtskSnRsV5uHVIBPbKg/ljivoYtFRJ2P+wbY6+KGz4CIbRTSKe8EMdhg
lalHuVqUoslc+ZKJ8C2SeaI2n3Y/m1NcLpFg4pRdNhDA5EkJE2t+04xuxi2V0O/9
Q9bLSz8fpHXLucKoaMdioPxEFkMDa72aqv3YpKkTjVOXMlbnoumwFIUE/LkvJGeX
xR/Rip6m28h2ZeKohVGIyD9tSvigtWb3XRs1/KhjVq78BIko2Uf9HMSF/NKdOMEs
EqupRbz6qvcy9DvhwQTDBS6V81VaGrqZGKZoiYXmF/HRol+jXHyQJHg54XSoMgGp
c15//Hq3yiBGlPCqC7epJoUW82/2gcBgCCTAbsG7QbZPVFbIYAdMQzA2D1Qms83g
tAxYqJlmjQ8+3Z+oXCrhZ41ujXHf8p+ggX4monv+XrtknzQ2UiqM9GVCTv39vqZC
glkd6ndkrVoRWXFjh+vOM8Bg15/TEbzyDU9jEOiuKfnzsFkGA+A097VhjEvFu8Bj
WS83H1z4i+TS9DZ7MWO60zy1LmVUUQb7Tj9D/Qesdd0GRzdR5y+6SBJ8QQQMGmIw
4Xyukfp+HCPXOUbos2Y5o3GFtHLbglwofRlBI0FV4PxCVWRvGYlyrSJeXE7imI9O
ldlKd5jXaDP7CQy9cr7ikg6uLjDaZNLMNt/EYlLUPKXo9jrRWF8Sjc2eVoFg/u9d
m2Vx0lqYspV4w+GGPqhNm6lXczDrmS4Dwiyy5LKg/07sxBEoSD7UOEjLz5u3tmX+
ioci05sFvWyYoo3oLZAgb1v4McZB4G8YAJamHB+Vdhq+3+/b+oPZ0+w5/oE1RhJM
tPg4FZjWzElIGcpm7KXBOH7gwyyZCf3tteU4ttfLejTIvFStoUFl9xB1DZzomDVR
I/0ByANA6IViay7dk9pn4kMvs+kNpv+D44p3oYjg5BmrpVtB0JmWNv0Vkr2U86Qi
qnEovHegdGCnkK94YkU+XaKexOqqOBjgbNW1og1JREMQbQrWchy1QxWGn3h6H/kD
m8Wx1P49JfPZ6D2h1Q1xCZhjCRKqBoL5I3FLBk1Pjyr6EnY35ujZqsN/mtwVhSG4
TncBSjKjCsbEAqCltlbtH6O32cb0u+Muf8wn5UEM03FCkoWDzD6HrXWesNcSE7TN
y+UwoTj46W5L5Tk2szcQGaZ2zEzWHVzJG+CJijKdonis/vO+IeWtUkO8c1aTipzW
N2lAbIHv6AKBj9+R6f+JciuXzf23wFxw/xUudwCKPDmN6e7hAPTLsHriPweAXcfi
S2fBGmi+BepNQueEhwE+vNqtTJKRnduEBljFG02NMX1LzaYhAyQa2kdgGsQ4dIbz
JnPFlsemzSRVWWz8G0qng+FFKb6dFxj0vP5gfpzeUp1/5rsQ8egEBfSdNqnrNU2D
scrsm4Or5obWNbEEBCjpPvd2FzSczTA+qiyKilKxnItecprr2ZHrf0smxmXswiIn
/Xe0JyQpq9lwF50SYieGo/p70OLm8TNiWQzel1DfByEG748LgiVtDOtIyJgKVTLD
y/unQG4o5D0wayDwziHt1zpQnV6w1OGZ0W/WdC2wmrQFyG0PkDWnLvOvg/b8fLAW
JeyyJ48oFNLg9s2/PxhZMwxDRdz1rdr04KLOSzjEm+KMgxUbawY3+dbgw55r6Mc/
pFODumYjnhgfgjOF+XR26UQltAXdVrV5eyTWncEGmWxBDM9u/VIs8yF8w95ENewL
fTTkFnzCw1mPU+nN5Ufvoaf8vHiJeVpQPq+JebnyI5dFRosB4atx2VD2BZ+HuJrY
0TJT4sa2AbpkPjB0NWArPevUerQIGBJMg0cG9cAaZLTiXTbo36HMQ32Pn+WQ1D1q
/YWQazf6vmjW8plnY2h7hqG29o1vQnNC2EG5zehioppIjRYsVOzMuvtRt3vKBLVt
ssyHSaxp8MYZhytEd4zj1Uu7DJDhuKaryw15eh5PFirae5mo45OeseKYTYWJm10R
pXyvSQo2JRdgHnIYX3J96K1iR3IIKzezJCnn/GaBVamnxuJUPe9JWq0ZYOQ7dW2V
7bizzOXMgRrxlFDcwkvBpWy2d1ej6xpKHSW4PIGicyoTPQrBxLtxqgZr+DjrZeyL
oVqZPMqF+nNTNtbRvj5IGZWZQXIlFze0UizPhe37+VRweWYbcjWaEd8QKYxkCQV+
7uj2ablj5HyAfgO8J34M2fO8sg1F3BVOWh6x7/mt5NWJeEeUY4tNvGMG+40yfFNl
7ag6g0LYacv5HLGzs78R+c1B34SB9u2ktMXT0x9eZNQeGOdodqS12Rfq0Pk42g+w
6GXeJyvgQJx5oTDODFOTp43ev4bYeacxyhyX32mRgAa25nLCWYYhUJ5FE8pMnKV3
5QJwkN33YllsjJWG82OAKbMS3aL2QpxKU8cntW2ppA+aXc2kjM1LFVEsTQf7adme
EO7saz8y4r4mzX07TBLpeOGhYkuyPVUd+5dVb2AWBlljz2oxXpBqWRDLpXw3e0DC
VcpI69q5NmZx4+duPhbKZ3Q9JkZIvodH+mGWO0e7MoLc00DCF4V6DGRphf7p5kAD
RzkjpxZjV92FCfeZzMy7JLIUP0dCvUlxEa0Q4iNHwmOaJzWWjwLxwGNN+VK7JCAa
4m0YkuGhtRtmbG6BLR8XvJxQQASAa7sq53Tzy3cKWU7D2DBm6MoO+92o35cRJDJP
AkVXNeyT2vLH8ftGZ0Z5nXEw80+H2YvEQtIkjctomD73HgqMJ5f6ORFHjIy/6MQp
WRih78AAM969EjNFdJc1bhnkEDybE6XkRrHTP1NlcMx2KiqEh8W58tHRJBa/eNGW
6rW6u//RgpgjJ3N38pM3xA==
`protect END_PROTECTED

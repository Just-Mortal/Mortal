`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcMDbhF1YzYjFCgQbLlSu65Et2J/N4HjErLLDxg4r5zzqyJrWYLYgPhfXrXB5HdQ
oipS5zi/oCXrw59mqtGMwfdtDDmcHbFPwJPDCXZ2kISeeJa4WpsqQ3NW9S3BqKY7
xs0Izsn+0Ras165GUDGAeRZZS54Ruz0e2luUXnpipCug3UOAATng3zXWVt+m6/jN
q27EYx3mV5URBZiXm7ffPMMYRiAwuMF38WBP9D1IHgOI5N7bq/ngwy8F/EXhGEoA
cn1L3RQENeApTnYIcZ2Isd+qsW/QVB27B2tk9BGzyPEzy8ugmkFj463EPp8nWAt7
FHoohaVD/lI57E7f2zPLctc43Ynzl+uG21icT3upwLbvzi6V3waU/2c/CJOY/pjt
Yg6DfzAZW0XUcYDa4W7hcud0w9gOwxPDAtEixgRQl8fbW5QFlQcqorz+m5qcIxFE
/p60OWO50hI+y+uBZFYXNINeXEuDg9kdb+9TQHlJlLIgnnyetzDSzADOXLGARsf+
0S4meW3UaJdPXx5nA7cygjA8U5YmHs3J/vrrt8+qWLAZqAeVJQLQohp0m7j/llms
LEiQb+ZkMFzFvau9HdGjonRSQCXFYBX7XgdxEKMY5oWQD7oJPvZgBjHfa4vq/7bb
zj92F57CbI7UKZPy8SC9s+5/KZPB1BSVDhWoQ7jZ/T0up/7A2N7ZT1ORalLFLBsi
uIm9bR+x07yln+GQnfL0GgVhMIlS6zjg5PST/F6o+GC0o3AsjrRKCukpk3j2xEo4
n2dJzmFOtmsONyCtRCSQuinZtAGsfip6AHuYhIKaB7StqcVdMzfWOttL+dCgOI8D
OO0omAgwjQT0rjOoRZQAemhJJbO/oOo3OaLknvGCQTJcDecc4PxfMJ9TOJzkwzSu
c/CV+iabPkjatik8KBauiVl1OlnIg8k64x8kDOFucvm23fU+WLev5GkNiFIaIa02
oAkNpJXBV+34vcRq4OxoePR2a17bpKuD5AJynKMlGxGcunSm1lTbrCI69dXPXULv
n3KljfCCsqnundnHRIGZZefC5GUE0n2Fip3vDl6AuX3sJxDF08zEf9ejl4Iup9Bi
VEnFXNeXiL4950uVghnBvZx4gENPyeIrfCITZMRgt45/jcWQcMi0rJC2olTy1ML+
n2gfVBLRwMU09+BsGD7PYaenx003Ib+TSVZ012ggI9QOvr+4X3qX86PkZwtSoLuo
xMtUbFk3hL1LjO6PlpAjbKja7wzqC8egmb38bgeUP0dgE0yrvhVhjhf+i9z3/ls1
VhFw8mbmXoUer7WG2XJUDQGkNnJ6yL/L++30SyU51nOQElza8XzOW/JjS0HlHQ0t
0bFfBU/hbi8RRNi14FlMox5sV51EEMs7nl5bA5QW8gU7SJXr4CXGBtwBSXZEi04g
L2wNrxX4Ijc2D31pSMYPQY/7ziiuWmp8CIEvdc5Uq9+A/eOL+/0JDvylRWnLXatp
VKgpXi0k8cJ4L7uMtdIpNHdzZqnqhFb4XcWCKnXTN0wpcmQ1Z3Wic6oPXtu1I2rk
97Hx/h3Wc5bDNIxkR8ebSXyt623JA7e9NszDm0QmVigb11qaAPz2zLcyv1PWRzIb
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9D7fhvLYWJTXjGw9ouiCS+51+nQumj5YtOsOQoeR2Sf9y3ygglk7/P0Ak8bSW6X
+5ZLMz+GGQzTXJJIw7Jx7sRhNNC4xocdqlBjfztHPKLbxEZD6YTeiHAdhXmpKbLi
9Xqq+Z9CSqnL4bsBy8Gdqj9kZI51y6kPpR8LkIXB05L9+D6WVf6pF86DyTWawBg0
jDlr4S4nWC2w2QewF/SqIJrybj1EwivlyfHoIYvtEs1ghAwbUsrWNr1O1LdY2HDM
0GNBJb/tcgdDd1eknO32CmViVltm7JJtLKW3tJ7+2wZzouSghoa8ir9frReX46Y5
LdUB92Vm+aSWih6bvAxkChEliMlmYnCVgPLwiD1oaZG4bcDlslho67AvaA6f8/91
XgEk/q9cm2gyvjKDJdDpg5f1xI4zUkjqWI2rPKIG0HqH526EBJmmqgKrPAfKEdMB
qgRgqrOcWZvZAfqifpK9qMG8p4HxI1WbgiZeVw+Xe9KTWhVf3PxMBmVkUAUB0WLE
98KkMUF8GqLjMMi6UZUg7nJOpSv5fJPU2bP3vaXDzH7PZTkC1YZNCHkmjB4Ap7CN
/GyoBXni6vRjH5T9ROdVYN6YjpCYD6YOQ+ymO39dszfDvl8UpNOihGOu/FEMr7XY
7zBhQI/4NGWAuss81IQlz2+U7LdVCjFDHgLWxli6eV5Ba095Rsy6YioQY0JhfQc6
nwSki4mNp+tpW66MrSHFIvuNV4LlbhVxvJLiyhLHnXsX0Yks5/yYghwvTnU9v+St
v4U/PzhN7wlgrxv5CMoLBOlHkGVIwYocaAxHXf7Ng1zuSmxGDR8seJtXaP9Oqakd
OHy5oaOO3SnvtCNmfriR3j73etiqTeHDtgzy+c9RqzhBZQwKyngkeEHqnW9CBV2i
kK3OXOJ3CU4RJlbncdWgvrGo8Tg41amu8Ok+Z5WeOOA=
`protect END_PROTECTED

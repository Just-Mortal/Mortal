`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xoBjxn/zrnptmDz0Uhq4AAsN37s/vASQ7jSZpIZ34vgsXMd29KzL/Vp9AmKTmc3B
Axl/2/j1DPCAv6Fsr83Q+7EMo/NxauYeDhz8gRtpBVC/ofzUOaOH5hRYpkY0LF3/
YjePAu8cvYlGRPCUXFdF0+EiVdEc/V+EVgIvwWmJZAZQtnt/jgHwMqqmUCza88lB
B8gOzFL/Fhm5rfeb/UkFEjIREs2I0cq8xRr5UF4l5X6n9QHyB8oMNT4P6ooiNisa
CefH+WkgnnO2HGGxEg//f2Rcm1xaAyfrEHNTE2tw2X5I9RNcDPV47BXJMU/81/gD
Iq1FuIawbDYGHvvjqVX8dmQE8O+bSEPHibzt/H+Uw0p38Kjsc9nTSiYKnXfO/xUR
AGY/EcMaiBwr3uk5inHPdU8ELJVup+IosbjHUCndxcs1N416sQmGmJ46vSuNrri9
DarbbuVyl+emH4zp/ocHSvYvR57h7C9O957zjUcwC/1/NM8Mbhpk5P57zWdNhCkO
RrdUL21jGPRGB8DnU3oiU6amD7MqD0iKdXuxGYK7zZ1ZWuwAOBLZXY8DQVj12Gsy
hcMF8r5aqMDx9IairS+vW804V/50xxFPPxpMe7pGEbom+ydIB9w9rUasi1++7q7h
kZ9gY/ZnG8ZPK91PiRu8i6IVQiCdI79yAbSBGYmkU5A/SUKIMxhkuwhHRrFvIV+m
5Y6BcLcOEyRLnKx1hBUD83T0opetZHE6eRTj6BAarbspea90LTCpG/5YVSmvIfwI
kakLqiqB+04Gfv372O+8ij8+WpQzYdxtagITZFw/nSDQhzxzoLhu5geMWF64L8VU
NNVQE+VeEGq0tYJLlZhoxTrFOq4YsnW0qXIrDUzf9hpUYCRUDKZP+1mPyhQyp889
+YWeKT8yrBX+2JuhsqlCnyX7w/CqWErg6LlxdU5/igG9NBTJ7j5K7NjOid6sAWjC
E8ic6tNwS1rQKDDZLZcn19b/x4t6ajX7vgyY11xQTp14blk4zRx0Qxm2pu//bn48
j95LLPPytPcW2GSSmtXn0NbLLoBlnNsbiUJzffietQpPMbHuvrT71wDJYTXLAGfT
zgicx/PCoPlXTa0+GQUQEIRSZnnQVQkpL5N32Hx5K0svyVJ9mQVnMwMuzLZuWUsK
fKzwJsVCV5NPXDyfo3m3YvAqaYHnRyml//jxRtsF1o04k9EBwtvQpMmUTkCQJJbV
PJOZNDc3NIC0G2P8ot6wfEPJYhgX/YHLipavjJ2MMYZS6gIx+17F69iHAOWnk7SY
zQzcIgE05gswWswULSzUwEX/VtOKKnnLHWkvdcPccqKGJaPWOKQ3eQA+2DWTPXnu
Za25zBIPE/WQ1MxpX876hfFbjYPG0n/mLRONIGjofv4CKPfEIcgPD5FsIs87oIgZ
3WaMB1UKq6PXYKMIz0HrZBF3pV2/tRz91EIKAo8i6h3f4/scuFDlU/HDxA1JA6T9
+Io7kcH59yQquV+B2t+WGOxM1BEBIIGdUfL0Qcr885fSEjtyEZfVbafXstXG8ozj
RlhNsk1DbGBScPNP4w8DsXM/7BmJnQSbyuU9eZUDsZ4CNjlcHQ1tEY3OigPw3jLU
IJC/zhlHra07AgKLrseMVQWhWKYMsrl0PenHdRCqW/b4ajrv8FA/4jnw8ea9AwTr
VjLoaBoAO9HdxSHaJdFG2H3Or6XiIgmx2pImq3LegaZ0pnfapO+8FjmotxnDCR4D
cI0rSxL7JqututsUUS0aBgLgRg48SQCIR6vGMC2vqpsnejxJEyHw/sLzmjqpdgls
KZa80Unk8OT/3bi2sS/xjLfSD3u0HSYV5oWxmdnUG9h0D9sYCl09e1w3wgY8rEjD
aT6AxVCBWl7cyvTl8K4Wx2E+wQL2SWtGNeON1cykeZ7Sgv8qtrbQkKQ7HDNcQ/uJ
f4+TUrLsxFmSreTALehtUc4iiK48rTeDVMG9SvcQTZ8Xoy9RcEn4No7KGUoI5hX0
l68trI/SppPjyku5I5/idndBF4gz1Pad5SGaFRsy9c8zTxXZLGhpC3toXzcNGFWi
MtxOQ6LtJ9mWFAg/fmQu40CdmkJ5v8io0j/CMwWNAeAMXBnKo/GIS1/soXrB6dmc
kswGLBJx3/fSG2RGCAQLHeZt/M8+uunrl00lEsP1FHu1Q2p05P1+8+gTUjEIWzra
Smlu2dpvEXmCAJOvpJZh9Rvtsym7p5NJ/mc+mVETuzHwuNT7uDsgkTjtFTUJU55Q
VlL3nPHYUIEnDXRyafI4XA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QyaY9m2uFv6TlEQFQE4cA573DCdPBhGYddZU4M2Cg9MsGyFQqwREuzpCJ5edUpvG
dpyDMAo0yd5x4+QuLLsQI5hsJNAcKRfbQDiBE8+EYY4W2ljrLGRgUSZFMc8CSqom
bW9YkM4GtGOmTzxLtBd/AyGUHCzsveZ55Yw2DJVE1o85DzcJ3vpPvCqSDqahKU3J
ePWnfwz3PUp3EesVtwWK2PKn2Ffp89iGRWVqeqU7vyEdWIjotxZJ4ZfSIAS56Xf8
TJAnWj90mrpPRiU8JnagP/4/txtPRXAA5QcpzL4QwfGKkhbZBOw7e23cuWzJMd+h
vNUnTLDgRb0/tiQk3u3PeZLmlGN+JlYmP4xEjLoYsgJx9mzfeTLVCYlMoVagDFU3
/AilNEYUnvqBJNT9YIhwNtr3hnIZXi4Wgem2kIeUC/S+K2HsAwiOOAg6IZNpC/J3
/XSowh9Wjag25GJNc2x0aXzjv7762B40ZzwP1s1j3dtiv2Ia8feDbwEWOmO38Hc8
7ND8JOxRLEnsMLNhycmXX6UEhlkO9OWKpFFNTye3DEfHfjYpU695/xhlwbZcqPQf
jTVfRIFhMuEDA50MjKw8jFMHIpafgRqmpS/Y+GkTzSjpj+URLoJNu8WR+YQwSvf+
3X0FxNrYpopRJVhbjYGY6Qf6tB6gWglKi0bdmc+wAf8gdapWZDu6Lv3oc1K8T4D6
2dUgJBjxhxyIinFinDtz9pOLsTNXLAMNq2yXFx7W0SweHSio7SlUGF3nGuBzTTwS
SBk4HIeCgx5HqEn04aAVxw==
`protect END_PROTECTED

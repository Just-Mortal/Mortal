`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OP+SSxAG8aA2YRBH6e8eO/8501Vgksay+1l6b+ppeqNCdHlybj7An19QjL4UrDB3
16SVvvbk1+wvq8iqF/5Wy5ud3Y7Ew5KQb5KPO8Gwa+a528vy2BquInl5PhIc+WIK
nhdZcigZVY2nm8vsBfC2PvD++a+OSiF+QUKvLfj9sLjEN/zlxOr2N/CaxU7q/nxN
WHW1SWRlsD82cQ0A0xS3YXI6Oyf2sSlNc+5wTKC9a+6PNjCUCVFO8w6GVhEqpsKr
c/2nRbt4K4LX4EqW5K5oh8rYmnpb+62DpDR/qw4RJee6z4Dx/H1rRRsfaoveexSx
g0QX1HkmKdiDQpDsGHnWtOoWiiw/9LR58xohXiRULuZbtJgQB0UabfynlqMZRM2s
MVP/nkFLQ2iyudKzh3K9y0KCLFPxSs4TFEgx8SURbJj7m4PkL5gyvGkaziAvWoxX
LbdFY55Pbv9zP2ZpregpA/T0Ul2jXZpWaReTw5fJdrlju/xKlHmu58LDiLeDAtC5
FX7EHBHwVqxFg5Nm6GJ8d43RauSk4smwenyrfNJJ9hAROn5xY5RbhLWGZuIWrFyw
VD20pv21ahs6XGVt9Gv0qdIDb+4J9UY96P03cwHjsfVcevCRHjPAqDiAbQ6kC39Q
9wdCPNDviRE6EvSymyxTOHjov7l28qn32qUbpJB7Ueom3+6M00fj2LefGWDDxW0z
PRpbJ/KHxgVUi0Fss5jEJymteQJhWsFtGad+tqQJWcuYLimob597iefYdbaCNAZe
40/fR7oe1tnQniYF2FXAPIN9nlH1YQq25hmPNiBAun+33C5KbRClJFTocaBhrrx/
pREkHKooKfVB7hkMENSwNyZx9BZReg8vhGo0kACr7ZfeBapUWnYRJydiZVAYtmMF
mSOV6fR4G/hxs5sw1oGau5m7MKD15blkpIKYkUnxMDQAqc4BCxtrCuvpdg2ZrP89
VoxecFc4lF4kNs2b3fsHlw1EtF1IIloJtBQsooUmb4ax151UNA+BuCOUPKHuHO2q
7kpnWIYSXeoSp2FDTaSOOIODrpw4wHPqZSd3EThc7hrKCEDj4OtvVAqgTKzJGEX+
CNydnHPWhCBr9znJ4+iI51Cg/BFfiQY9QEq7tWEWa812zhIBYe3YRMD7CKKjFkBq
ztxLe5+BqtLEM8soCIp0wyzZQsQ50npccQqMVKegFi2zW1a07lfyB7Lr7jb458bn
mLqF0LAECTaKhT43HXt16AvE6tMREx/GCgmXwOUfdr72hAtRpAW8GZKlqUUGx4JH
dTcb6tv+hOPukpkfvTC6Pr2U47wj37Vnf/CRgI8CeDnziyLIevfb5aYbr0S+1zd2
dvDZl9andr1jB+d91bgf8GcrI5w8RpVuMXM5VoTVuSYwXuvsGfbAafhpzJpX4LVx
xiEkEOsf+CXzleBnTf5i74Jrws0Cx43HcqRKEAK772cUFBtpT2AMcY/IV83Y488b
aykBcPuWNVLl5QcT+gPFY5DknOGMDsq9dAoND4Aw8ZhmtHzHHySf6vKxMT3JHIGE
NPnRXqfCjwjzpJ++qT+UpzcCHkbwvgVY3JkLkqYFhCvysfYvRKGhYZmFGf1e5zK/
KxmDqdJSOu/Zub+SPCUhrurudOzQUQhTDvEefVH+GflhU9tWfwaAWGsCEB6yudxu
8EZ3RvlIavNBwmBkQ0+ZHld7oez4YdeYRbTaff4LRmF8cgk6gmWMjYBUfIXxUFlw
Fxzi67Lf5n/H0yH1oTfDX41+awoKoog40pQ9/Zdx3V6ZZvZHY6Z3fD7yS2uR9s4R
0LpHz3GuP3xL1tu/bmhiLz0QZX1l8ETe7Eu6yAIPnmEI1JoTtklMNVHDS4wzjbpC
vXkyiQxfGPettFiCNS5uDhDkbVojdPLPR9Pz3IMLlMxiEJjdcloll1Zpa0/HPvLv
AOLjvMXRaBCRGAYjYpHfYkg5uf0mHxku/mKpqm9CZfTDQh67gNbk+fX0JwCPWBLa
8OGbrWv1WMBANEiOaPNL2VLW2jcvXZacHakZge8ioHahT+OjvLe7jw+c4yGcBp6N
vZ3VnR/UFn/7yYqyypEbDCGrXVcxTnZJBtHIyRsCgbnQpzUvXNjfUK2JPFFGJnJy
EQ61uhesfyWN7np8N+IWxUkRxispPnBMQX1tA/L40Td63842iSASUptwjiS1iSTA
vluGdf8x++c9Wr/AHkPcS+XZC7LkyM4ib+OCOebyv4ODAorGr1QkzKWxENRMpcpG
eszu5NhdoeemP09zbZ9CL1aJpqkLbXG4+7PbvmN3/toJtJZx+g8zEOIDfKBGYEDY
q39KNlNTcTNOlSroYZUvNTD+4mOgOWUQOerqci0XeYxWCQt5WseHeqUx1lTNu8Qv
+YaAuaLYG9zSTVQRJNX4hqqEpUe2FB6+g1vHMjTMARr3eqGx/k0R24nFpabge/hZ
V+phyjz/Ayel9kI/xPZD+/G4HEB/t/xYMZIUPsFOP8/viYEq1ARjzbT6UopAcsfg
STvwaUGhjuySt4jd8qcE5yGlvs6y10n3IE2cLldAhpsSZ1EPYH50gz1ysFpGAcwO
vCh+/m1uJUvFBXqRWS0n1BQ8HRb+nyXvNQC2N/eh57O+ZqV1fc4TPnSqGrrik7dE
hE++thRWJNH2lYYbxO+4oAN3qsstRi13mPAV0hBK5HPePN0kqAtDRASBdVodLRd7
E9GQgcIRlnixfy9fDSsDX4YuzwxZh1i6GeFPYSiL4dFGtBzq3C+0w1nHMyDl7mOV
pQ0IgIEc0nRgVDL0ZWIe9v30SBgliYHwFNJc6VHLgqlhNo+g6J95F0FcnBjcs1Y3
dvEGqIB8i7KvNAUOMg0pIK1FM0oy4obotkvzbIualo3TXmYuEDMh2BPFMJlO8DMa
mmF91yX96ULrFw+3Wv6ezby5GISM7AbuoCunCrrr5v3W8GabR2lQE93vgyJGFD9k
ZkDCJwl8me7At+DmXdxAPOHog50umYaXtlNBR+/IM9mTWcPO+vqnNy2O3eyhGy7m
HwPNgBsnY+YygeFjWDhVh87P02ykPVotWRAtDqDY9kAcADgezXMyU1ZcNT1pOCe7
N1LfJUkSEA3kAHBxYdj/V5NcQWVBqmJRkW+6hANF0n/4yaaXFvTeGwcclciMbiHq
/pdHnmO//xiOCA27zp9Lt5ZhUljbljE+Y1rI8Q8CCrK4zY4c6tg31kB6+eK6M9Qv
69lCtZMhYmS/Ky8nD6DF5QPIngqSGhvnfmHfMhK+Qxrb3NZEJQfOlH6RmO22mUQZ
DggBBsK+BF4fQxkVe8ewUD6ed0aup/vzMyM1LMAtjKjozhdhy/7dVvP+GmkxD2AE
tJo+tnBjC+SGFAeptajatCQiwsV9bd33cbZv1dlklBmSPEl5DvGqwk2SVeuv/aAu
BtGfOGO/AK6TlXgGErQ7PCJkgrtS8ayQlNM7Re937ORPRdHs5PTUNZ2dLPynNxcx
DQCUMfZdLl8FzjeFzoXE6BOjWWK+QrdorjLB22sLvN70pBj5lTjKXldrI0odiISG
H7cuQsILZGM/IC4CD3xRrMBLegNoECyOljp2kWn6LHWtDynMgKpaFAxZmvBG66oo
Ls9LrAMLEPYfpJ1PybaQAkQeKjX8nZWqSzXBZkJqz621UXaDBXhza3cCuy9uLB4B
raL9dlPaZquPYEafd65ukOQt6/4Cb0bLm5Te3sRRSTkihtWZG1SBZKBu6XzL/BwD
jaaf8fbcl4x73mDaJresyxjCGfh5YdIIsl8O0/9/q0tId5resS9tAkJ01X6eppUn
rUIVtflveOJwG0KxP51t7wIduPDzumhf5he7l4oxzDYZZl4HIhVV0MNbCYlGPTpX
2MTP1ORCnwQVadoD+6xBchsp2N7BcSMPs9XdA0MKF/TMfYQpTGOpsVuXZI7Mh4o1
VIg81Y8hmMyA3u9HaK1jM6qmxc1IqVhu9/o4AEt+RNpLttvGxmM7ujRAIvDIJ+PN
2k3xARQ4nn5djxqgzpiX6cPUcqx7pgAdsqV+Fa5Gk74AtzE730BCGsA/dGgu78En
Q1j1waSSDT/RfynwdkLzQEotXutPkHSFR/8u34YVsATrFN8JWNQjX9zbUvO5W53d
nQ+Jil0d+ib5hcxUZUQ54+C/3WkEyZVQPZtduTydgC5vOgtLZmnqFiYZzpDPiYb0
6p2qBaxq2ZeMfYDe7uYn9QYW6gwC//pwZps2P1Opi27jDW78Enj9fcti4Te02UBv
d9QcwzOUUXwR9mGer9NT2rSAs1WxkHhN96TBZ2ckUqWR9dpje9X2gipIZEqgI140
mBa+43SLsa/ymvABTKAtuEG6wbfL2+20WIoqHV7JCkF9Jqs0C2UBRw0jm1TCS4WO
kGjCgit1t67tDJaut8LmJLo3XcSX8zxX2KhylyEudBRH1ImJdlGJnzJk1pawtym2
/HKaP029njOyTx0ZZlko4k8xTNnNhk00D9fs4DxzgASfR1FZv34wkXU+MnmZbaJt
qXSxkNV8t9AvK/8p7E+U3ZIcVoKqTO19uA/aH68RzykJjy3WibtSqRymUf8OHzdo
CbG+6x/ofG72NIIDMYVmVVOvYxUaa5N9UNOfLJDHYJ7pXZHViuw7zrWzKh9R+dcH
kD43TBbMhqbCZlcPRVKL0a35UXjkNjy6fgZWmaeWg5Jcn/utZnGp4cNa52MvQ1ir
0UklGV/NZH6XKtGXSuDh14aN4/y5TF29///c633+RB6YTm9rQa8Ex3A3FeUkvT24
qk3GMXmFMfZnhNpStmn/xQoT+QZFX9J3mOZw5n8FyJK+aWqSWEBLH1/nosg0dRKw
EC8vuQ6c9y86qcYgKU9mIteWPxR6TXVnW8awrhgCEh5kERYwaIC/9+UMbYoqG8g5
9nZAH6umJHOaejGBJZwqq1f7jToV3v65bUDS5/D84C25KOm0a071PqYphdmIyQKr
EEjGKOp1ACkerau8mwFyu1m56QFbC5QIENWIDfbGyR6bNF6xvdsr5lVUGzFkBpoq
oksoxQqP+MCn//erv0nZYa/reuQSPspvWKhWBFcgzfvMTjaeXx6bVBbE2W/jWka2
15Wkja9L0VUStQOE9o4M24dmXKP1Wmrt0XMzhCkwi36zSgK7d7WC4SkeHoXN5/FW
q5y5JK3iRJgFqxqJyDKCP970TTnOOzU01ceUhMGItNvkqntOXiD1hIzqJitkkk1Q
og1pLmPPmbEdkKe7mO7uEPz4vMuoNIVJZ1fogKmWe9KnJrxDeVeOY2UQrllguZQy
sscMDrMTSDgKMVk0QtbdVrcr+ijKuuf9GndzoVa/PWByjatTgIN48Hgjx1MOihjx
VajASg8TY36sUEo2znFn041yBqquOiwi/bd9/sFo9D4YjhdbkDPFU9J8WlEUs9gG
VaekSORCx06tvZ20pQIvrncPqgN1+5juvwnUaNCgnTop0PFPgaf9+OlDlbZsgFIo
+2xv4W5eGu9211BoaNw8FqgA7IfDxQInN78jbr9K9aUjF611hBkCQpLNr3ZDLtut
/gZj9d2n1zdYtr9sC1L3GlkLignDogquJr4lDkchP74R1wrYvhokJrXGNyVEMgvR
YkmJ2P2wnUmRA9x9kVseAgfaG0qvpvSuxlzA5z1oAVy/q+o7bLSSPrtlAwhpyXV0
+NVBiZMbe2m0usob6zs9xTZwduNHAYt0ViblL3ZrI6+bSF7KKmb9OpMeXnU6YHL4
08tXks5KgWD3dFSBr3yc6+JtDmnhVXi4mbaOkAerEers+QU1Cs2R52roPW7ckIP8
fzRoqToP23Uedxvoh+uFv7Cf0WJV0rP124UCaCQi4mJFJXBTAFfeVkKnr+fTAHeY
PULyWcm8MnXyrjaXWJw5pWmJfxP7jP7l1aIm+uFHgKFef4sGh3atojl5yjzzMsuy
HJkltGpjqWXCc4teo18XM32vu+RLaxwkNfz2dyd5m+jozYg3oFewJJjS4YG4AQC6
qhZf4aeDALnZqS0oPVNu0GL0CqNW7Qiea16GsHVojweGIdsUC9EzyR8VMIl7s17E
oqqBmTNT4bamBaiQ1MHwC+Zq1v7H8zfbwMBrSKm5Mb00cst7oz0pzPwqsd9Ee0p8
fcsR06XLYIetUkDLOa1D+tTEvbKcMGV8d8QPvpAgY/xkL2Xd9WKMFcPi3AfVE0S/
w7LBNWeZvuNrWDnv5khB9WaVBVfnboU/M6QNG/4FMzvszyMIdYfGTn02vFBrHHys
xWMYq4BViOjOuVT68xRh2niACrNPKUPCCPP1L7ocLrsHWb6zHM6M4Q13FsH6ajle
zC2m7iqiqLgPjVu7eS/isswET3r6ERnFWuw1z9+2NB9IvfP46dJKRZuE8eYmYeEB
4N26GiXVYwj72d7qFhTEfSHcdxa8hCuzNsliapm7tG3QSbfS05pSw/21lmuntUM2
s462rTneO/ZchMUDx9bSGDDf2M/a7zk8VoyP4EZF4XssuxD8sdl0o4EvwDiTD48m
ivWTG2lTBg9VpDU7mIhbebEOno2Wm3zepyb76FrNdcNKBJ430bJNrWxpEtB7aSz7
HAxrOo3DUvd+Sm8BM3PMvt6FSsTonfv3uJQ44NftH62IUStySaqJqLY1l4lCJPeA
KviLDo8bS7R3gZtvM7qxSY71kX5LQqKFY/au/lRm/SU1CO1x5zHmgxzPpTDRnwaG
jgYCD37pIj771YRsaWwPVgxZcC0r6D0gfccwjgD8nAaaUj0fEYoH4b1d1cxgSZPI
OBEYnTLNHiJ7aOWLcHOdblcR4eyZq/Epxx7GmSR/89vn+67mcO9+wVUhE+f2Hf+m
8fCO6zl01xwSO1nEc38j6vRrPPTSvUweCLOhxxqrD1ZsC1QKM1nxIl+7xGcJDNso
sM0ld73wx+ZVa6vkpD+UPvfAFH3c4A2yzRBZZjn7A7eAyidumlgbvfpyODjeUnjd
Fjxz/wPxxnFh5kkK4AJFJET2MTgMklJ5BIh/j1FtS81JbNRRQ8KuCEdkL4fM2zgR
rQQGWTM8+jaNxAL+1ndmw8f6RIA5T7dZmArdfJV7PLOOyFwNW6nfpslA7P4TxbzM
t5PgiSOMpAXqJzBBEm8sE/O3l14ATgkXdyvlku4QDE1gmtVMiCBDzDuCi5i4ce4B
1eaN05g/CMxixKJM5AffXEbbpuTrdsD1pX/Iv/0w0+SFSeWeeVB5HXP6B6oytfYp
KUW3DhKMBVphKa3coh3db77YYUdrwnBSVr1iIw4FTmazqbNo2ZneWJ57PWT7sueS
/aM1zHfsYVwVQFEOP3bDiNPf0NEUPI97qeKzMyEIhvNDYKrj6CiFOZ9blE7Aytsw
vYxp67oMkccHi435pT3AveuUfqpiI1X8/vsAHqQd5RYGad6kppZlMI/37Td4cZbC
sJO+cAoMLVVulG9UKyt64nfR7mBqKo4iPeED/sd16c/9Gu0BSJna1+hU20kpOf2/
FSxYPH6zBAdn3pU2Ov0J7ZHC32/x/DL1CP/h5OfO3WjRluhdO/JoXBILmnbvT1bT
EDGJs6c2pDDXo/QNL7E+lVwczzg0e1ZRmuG3tN+IXPbzDYJ8Sbn0D6c820aS/2sF
tAyQx2DSZEB7PFYVXrBXQ6nwp5qxsb0CQYZ9j3e7YGYwFGUjij2DBGxJ/P6LhbNB
PjC/GUuYvmrLbbjdDaI/rfYI66liayzB2AYBeIcad49NSM07TGgT901HPJ1k7ZET
yDyrPJfOHxVzclC926Zp4pfwoFlw9NqNZj4QyZGZgD4M1CK0F+9JOtHKgbIILfi2
0q6Y8d9vrzfCPhmAVF4l8N6MvabxcsQajj0FiorJ2t3qhu1b2vanFYKnfz2Mrm9e
tBJFge/QKnClFYFQYXipFLWhWMFEW4p/G6Ye9+rOZueXzRDj/hJlgxO3GeoYJqUm
VbfcvoS6ei/t1oMPTJzlZhDoAO3qXqTnT8umaxGAKQ1qXz8y7MOsnCYblT3YNy89
eY4nXR6IzdGG238yLO6ECzo4ddgbiNrzuZqe0Eob0KfZ85m7EOskhABDowt4LEJu
ZdompIF8JzP5fYmSNNR8wWopIIlUPxHstucMhpittLciQZzT2ED6KaGi4p78bqRg
AmY0RQdS79nky6WZj6MdhrnyLHzaEIHaa/cjCQpbKbKa4dtaQHGaiGz96nCJREOu
pJIfV/EYz66GhA1OoC69xD8QX71VsQlqKbiubPBOrM8Hfi/o9ER84eksqzgInotg
/qtEsW6iW/KajbhR3rbS8a+oTlKHQ5wzIOQkIBilvK5Gz+zbSmH2CLF43bRONHVt
Sl7syFK3790VcX5uI0ejcegsSSVTTAugLK12qJQ/RmPPr85C10Tr0xf7YXg9Tybp
uB2Vmb40QWvGUQlN9DTtPt9wyMl70SMaQeIr622gaZP89QgAHgYuj3lKEtaTdMU5
c8sP2iAW+ljtyy/13PZDMpAYVrhNm8/2v1ApTotlLDaclOBN4+7oxvY+vj+etXdr
Q/DaD9G77bicMRtbC1nSvW2AyYouB3gwNCp1ZPRIURjHYXqf0+UP1+jfjUfn561y
lPkc6eKtqPN0dYlR38+hjUAmlle2v4ukv8uYuWGuOaEnaydy/hByD+PR9zBWt6au
gtt8bwDwrW7raWol7Bss3hRNOlOwxEjQBHtzCsnLLsGBYP1UYTm4i22DErr8bnXw
uXZidUocxhAzD431kokITvPZYPJXAgnIPCpfgHzmaL/FdyNAZ6TJJAdPSIMTuxi4
89u/op00PEEWmxLaWqk2gtGCQuxgNQzCeUA/7ha0zJYI7eDBBNRjs3mQEKfcm7rm
86cAoE3KftdJ1fg/s/9p8hrnBTheL9o759VA4iQeDIwNpyxBBKLcM0JRMGGvITgE
nXlKaL/Q3onQ4xE50ADKkWmAJ+cPk5gLBhBAbe/p6QBBw2VotGP8aZ2Rxh+OJRJs
yItcoph2fC6YqMZv5TMG42M6rCP7axYy9GTN8yM7eL0/xTEY5JHTQ+d21HbXPKnT
WJ4G4H4sg8qIKejerv/lI5Qtr9uPyJ9OlR0rj/5tWHpY69Bgj2oL/Kzk+Ef47cyU
tHGq8HN0yzDc32v7aIc1e+Ck5p460qNfMJtaEMwAI7NI3tQhJ1BTgu/Vd4Cs4NDU
vHlruPpFfu5OOu6V2nW/9HDgIgYR80HMR59eWaxhrU860ZnAgWGtPj4KlWk0BSs7
aYwVVot5UZcgviFikVEMOmD04uYymh5tNgJ4cjvZL43gMMreGbnIjrjJZF+M3rq2
HjOc+yXk3IW+wYLDQLU8Avd6hKDKOOo+JJkgYDbWjKGKTyQd0nfYvYpRelpoc39C
OVdRhdP926ZBQNtJtRzha4DJyRU2zxvIgW3rAAo69ZtH8gCzBE4Cl/+m2GbmFQ8F
o86uyFl5NRh+Urg0d9YA9fs6ASfjUvYSikxjknz4/O47FgQ9O8/fowDktpR6+D6H
J9iuu//iigwnoA/cclFIjhLRHvEZhhJQHepusIAhRtluyx8VyQLo3l0SGp8ruoPb
maud5BPlQCtj3TKwDVBMD5y0OzXoyR4FdUAaoBuEjgqaXwq5cz+ksa/i3B5c7l9a
eQ70NCzSCVyZr6APWAoH4TtPdF3q7KcrDwAfdwWW7SqTlxL8oUHYQq34BZn6HUW3
S4axnA/SNqzj8+y/ZH9bMmH9dXJguE5RPKsrgCccDgu5uJx9osVRC1+8qkK+MNNe
m8/7bkxQNruSTTwPvjFU7bYi0ywbVRAm1K9/aiEKMDOIp/dXuDp7ZoIyfuN7w2g3
OpGX5jfo4+vQcp/crQnXQqJFfvCHdjWUUyRiEusxP0WUUwCDW+MIcr9EbqhNjcGc
rXSY2r/uFAJ5rQVbA6INyUNOMFgqYiv5+2lRKdJC4G7K0mmJbnNUlGQEwyDlI7t7
9VxPVsq6UlKkTQi8V1Tkzf5y9Zfmr7MoGl14zh4cPuTefdbPt/IVCdlIGUA8h10u
C4iWDpE5AhkUuFfiYKH2/JD9HjV4YUI4JhI8ouKZBICPpWwEv2XhDgDSJbWUDIAc
Rmhk+q2Q3JziBZu/UUW7secgLXz209dFDZjq9ICQvMYv/gQEQBeKUdHaMOFRgfr2
gsKpN+tVs+8RLr0uA27WBFJ6+OZFhHAUr5q122TuG+qRl0GRf8rw8/vlPMrdFqV2
J6IxQH7HVm1SdG3+lDfMpQ3ylxCwkwT1Oeu6bYqYwgi6GX8W/AZzb07csXgzj56A
pTlgahyO+pM9dm+BRvHu3pOEXogNce9nu2NroXpq17/ciMo6PoDg/R/JDRRVRWvF
CP5d5ey/E1ra7+IjRlqwJNsPOrVy8R9s1q3cWf+XdjkiOdof6KSLZBLEZEErpIlW
65X3hxHRMhzJEmCfiBOnjJtcoibXjPDIEBvLUuvF3WFCOu6WiaFyv9Jd7ihl6j7Z
cg7JybAuT52zFp+HeteyTNuu63wwPXhd0iU1jSjfWYcRXX2lCwXL80hTqIRvbauJ
DbfvphyoINkm4x2b/TQj8W5iw1sSDF+nt3IHpxcWPGOLebpa7beXNNFvvMvyJ3g9
Z+uNmm1E0tCsEvCMupHPDjhFFXNrNoKio9hqEDCExvqaLiYLk2YkPa58uuA0Zptw
JTJhm0kBI3418FOBdftWYCBeOQyF++/WFat5vlNybxGPXxSv6tvuyZbYlZmLc04C
WYo+Xi3vH0nSylJZtViN1rZbNoAo9sDbml4GJ3FGNfMtVi6kF1PyBnmR6ZPXBfe+
5O4BVM2LM6l9xTd9ySBERBJ4dJYLsP/hyoDcnpjKWg8BmY6e/hg/sKnD5pIvSDSc
bXPjfXLnPRlS4Jzu9aQrpWirVNmbNGRGgoZe7pZU78c631DPe3JPJFpz1GGTu6ln
8mUUOeVIDeeY1+DRVfgznhtKvVRJEFnfVCXTZ6OrjeFJWtdrKK56l0cX100lWoHr
FkmvkwC+9ZntT9jZ9vZJ4+fbtyoklo08nxoH2xR4q1rDjYFiIz4KwSuZikr8NgEt
TtkbeZ4xKoxp98cNFP5HU6K7jbNo2mcdCr1tQdpxjVFK71kePYK6+Gbj0fs0xXOh
ZKxarlkhG2JCbJEBzM3PzK7TQ6N9/yXY6M/q0HXf0PsRdhq/4oO3EIESqm4oV14a
0tTPiFOg3X7eqYwqGiRX0PQftpVM/lvzRcvjxxW5NauJntjSJRRbd9Q5DyWiJZ60
SzC8s7LinfN5eKvgNa/5C6pT/3C1r8aSJciIwHu1v21N9tUYi+ytQuq7uLNHKBNf
To30LpP3ciJly8fFn8y0u/yygqNW8epw28lRNcnmQaIGEjD5shL+x7TSb1ohrRVr
ICvQyOhlioL/Najc8/h1ag==
`protect END_PROTECTED

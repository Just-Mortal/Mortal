`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFyz+sldqnSILIEUufbJSs3U3cMPt/T68B5FJsrkR/USCOaOuxFtbDrOB/II/LHN
OXG/NW92zhXypppPDlNsGn/m2I5YkjRk4Iq/CbSt5zSZqrdPzojJjRErbD0Jv68A
p+4ofTfNwONQD6QJ5XVUjkVI0D9PfggGK4umn+z7Ndkz+TXh+soF39ZIHmEr28IX
qhqGzlJJjxaOn8mBwqzYVeDPI5j8znpW9sSxjI7DDES3XU9ij45E9Sf1B4ihtxRg
7wcBofGOPTTcxH2GNob4jHqVfC19hs2d34gvAImDFU+mlnnbI1ylNPos/k1KuF6J
CZwlukWNYPp2azOWVf4yxFMK9cTh3apFbPHCmwDll/8TMkuolj6+ynNGzdrbgBN4
3OFiwWv2DGBo1sDQqesIE8K7lfyz25wc2joQnffR97A+44oerTNsupbSKb/OJyOC
xYYog3nvmI0kzkB50acPRCdzRovKavz6vzyIgosbEXzC1ZExeD6s2qculxRQLw0Y
ApCwTI3Q9s63oAwR2vLhTvh8MhAOcIS2ta3qKWWnh5e0EE5h7rIqRY1RpO9bFnuG
qhg3bR6LxGZCtzG65LabndE3uJ3Oy92tJjUXtLTYQeV2pqCjs52GOYTOC8c8zkaN
WOQcO5/MV+sIajxwwTfw1DI+BoIfaaKGr2/++821QyDSnb2j4s4Ivz/WdyfsAksc
q4do92Snpl3Zx1EIIRTIVKltwz44Cp/KDid8p4YyWeIyrG4NAICFRBXQRDB0NTuz
uGWAyjW9w/UUJkFbrN5GL6o7+gUP1SvNQ4zg7B2At7/3KlEyh3lPPnjWu+yTUEpS
+I0tHyn7RGvG169pIEGn7vH3YV74saQEEG+ZvUzqiJj/r6YXzBJAO+avh22d5RiZ
uDAbEp0tMEbSOZDmufD1Tdo02ANGu5Mt1aCmMZml4OWEW1o0mRoZq5OswTq2nST7
KAeOiaBepP9Z9O598zLjhJ7Cs/K5zv4uZlFr6ASG1XHSAX/9MCrmvy6ySp4faXqs
hWCz/2tG3eFEhbppy+FRNmtNP/xmGr2KBSkMuve+4eHMOfPVtaEKeh16MxMikPjf
CtHfZkf7DAgjBiKRaIocrX6GDsc3mm/19IcW+Bh/BqkqSb9GoM2gcgIh0YuIU0Y5
sjIYodW014BaBrdiZJFQC08UikCu7dRkUvBOR5l4aZAmxvGRFH+lHULbPGQt3RBA
V4iZqvk1JfOL2GfOlyMxSvw8K3ZBsJQ/ouRPhJ2rLYlznEmM9yKCjJp5eaemig/h
uvOK5OV3U8RlXXYPAHXmc+gqSDsmr9T4VLD1eLrFeAw7+Qyzg9QbhjCI3dsj41de
y+hcmTrzp/FiANjf1JZSujlABNYF2gyefO0eCj59hZVIGlON+3EZ09cTrn31ecU+
CTY+uKRDgTn6T7ZnpqiM2RlfFm/0zv3Bh7kgfsh5EI38p4lC9bTJB99UVtpxepvA
lsgfDwlg0aLnjjod3MfrtZOict5Vcih/uqZnq2cjtyAM86c/wOnLFkreAnZHMDK3
TcUpP6Q0WiYbi5Q/8N4+UX1R1zXc+zq/x8Y465JQfWSF0j07yD84UxNpG9tnVcek
AyOZpxGN01PbSrW1zVR/5Q==
`protect END_PROTECTED

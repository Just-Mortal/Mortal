`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4NjhvR+Qps1n45LFfIgnblZm30DP05I/nrb7kBOpOJSB8oB5FR+/CIWyJskURyO
IDc7PHNV90Zh6+E7gact01DArshKZTr7V8JK7WQ3v/gvJxZqBPuiedrpjH7iDV7t
8UT6YhfS8QFPTF0fNmaWDb4I1qrXo55eTOQzariUPefU6lTNxRy7Gt5yt9MEyuIl
yEu4wBSDPKUpvkP8HzIO1PLoKIYdTpikmkFRpQAfsKDWgNFX8Y0/uE+1evedG71R
OHl3bEeUDgVRcvb+BO43KZ3XGqQzURs6mtw88MlQopDMQZo20CkhW/5XITj77a+g
g3mhopr9aBHKf1EvJF+jBIvsSqxpHoWxnuvZVz/8F78IThosXR1EzivYnRmJuY/q
s0/WNmRyFlx9rQFqNrbLW4wHFMSB9cJoPb/kPyIl8zsx61DOb+zmuDXk6kM69BpF
bYBtzJ+pzwC0D0E2N7nD3xFdCmS3vHEsSMkRTXzihNeJZWNipKzqn1ZIrOtV0eYS
ukT6IMovbh28jhOO4c0L2VmfJW0TdPAM+Jmbhi3sN2AYm4GxmJT3axrl0dtOjRYi
bbTk1dGQOFM4FaDhxPeT+hXZzOe8NDEjquBwRqlbZ8vz2L9T0lkHSxtn3BTgkZyX
tbrwWYj1/Z3yL5rhnagYlJSZ8KFCWIw4mAWe/Lkb3kgsgPlimcVljM4S4us8eKxq
+uHwqpljFrnp4d46ev1MN2Dem1pF9lyR84DHt0ejqpNwo0bViBaZn+BhSftAnzrm
mgkYJYD3ac4HcIzkuUTFSFIpTFL7/seQ+ZzAIHxBHBh9UQ+clwC4uRtY0tnpxHT0
k0wdI7vNTu8l2ZFS4HbvY+jHdAwoSaRAfUkXJgH6B2J5f3ZYWvN1NmjS1u9N1+BS
wLeYS/ObHsI3RbIzRE2Mt4WpLHaOiuYOGOStxlQKQ/5+dcYfeBNA5DrwJmgGg4L6
xNfwsu7l//vvl1LjaPX2shleQ5NqKCPZtAIpv/S5zTBRah4fjhUslyAkhv2+AIvR
dosfQfqUyw7y9V4b86tMGirovxVs3O/kyLmS7r1UZoclKJzhMgqZQtQojg1MN8YA
Kx6CZ7g+S6xWHBiBXujrtPAHROARxk3uqzlLs2QPKQffEEVOyG0D5jmrnEPVbA/e
WLx01J6BzMAPHOHy0K1K8M+qNi3uIPjtFzsDOAowYakA6V3GcmKzVk4Ie6HT8PD1
DjNZi3MluRZ/pKvJLVQF7Lx9CITBo94OWqnA9W1NRgOSNqMEoiqD4IcOxgIQtPcc
UWHLmd6Tv/9tBSN9A2fM/f3OxeeSrfeAUTNQH2ZEeOCa5o/8lxxDw/0Wf/7+0oDH
1Xxyeej1RrUehs5GEx0ZQgcectfuS9nxkHn7GRcqmqRAS4w3PgRZVRDUu3WnyqTa
lIvdQkqJzZ8EFmTcmTbljrZzbXFUXAVW3g7sYab1h7FYesHQ8ng2n8YVvOd4x2PZ
cjFgdq+EBNN7m1gcx/mCiWcj2CpiDuNR4xyAsR45JWHY65+xD4ccXcBt4NJKBF72
EoqwtaBXtf0GVkUg3qKWaABVsigPycJYDv3UQDfdxTW9SpIcgVMpExJ4qBE8/eu0
KSiu+mQ98TQPDB8ytSxHyOj6IaORh8WeA+3Hjst1p5RfzVmUjOhmvtxL0w2EOSQQ
/QzgXjtOPSzr/ppH7lyL6ndyVYtjEWACNwtd07OO+EOQvNl2bPJPgKEzueQsZJqj
tVwposPYVA4vsj8OpxhpZ2MO3QI2YCSQkrZ2DR+XaN/dmU1/qfxo7CqZSkEFeIxL
Gv2BsQyNL3z6KmYNNIyxNxSVPP70BkrSWywJM9xIfBy+SyweMWyRJe80JBSWxHIU
DnsRzeRKDm1C5Q0reggOI6ymiotHJBEHAyO1vQPnxATKxNcBCKzlBX74b15PBSIp
/dsX7t9dv1aKiV9u2GcEXpJN+Dfhq2y8zIU8Q9hTgIBmkss4AqWUP3N3Fds+bXGe
c3n/nyluGf4PrI8/rWxJCe2+MPmMyOh71cDEx0otIKGRor5Jt80Di5BZyDbtuR2j
z/+Bi7xyLqwChzL972YDWsWXbRn0h8JV6AeVK5yh66N37uGPzd3usUhV+yNI5L1f
AH+kOYJfZf3asz905TjUWcRp6y2uk9XtJ7JwYJTko/X+3pwutTQoBwv6aCVqNVb6
T1aVJvOe5TTfoDXc4EiPvAYboAEmlX9mN7m4hY6XK6sy0YlPDXG/s/tvPdC6wFj2
GrY0pjv9ds3JmPTVyiZN3vc1zCNs3qUpN3V0xiKCMzEoeuRnjPnu4X9kdl7v25cM
PCpm1KZxoaBN0IO+A7lrBhgPdC2WxpqQbTKzZixtS4N6vTsuCh+HDdwRpHL6/7Q3
Fn5ESAnaP395cKUiTFLo7DZXu+695nZK4SWWe3Phi/RbXO74kj0KXzhT+xLTvEUW
q+NeUs1799ABPUlRzf8lW61DgSh//awjhJwm7jrpGPvJr6PwFp0lBUPXegRqwsWc
LT7YUQb5Kg/anAD8aLFplYGSIg3BfLyLVaUYF4d6fdzL6tPs1qSwb4fs1/jTctYo
eZSmi7GjyKrms1GP2Vqj7sWobtfWn+Xy3PzqF6Lec8StsbAkyTkQyQsUwqp1LI4T
hd5qxWl61JSQOjm8kouGpDpPoXDZwPDvqbaoZD3kIqJ2sxUJLLP22rRwprQKlzMC
MRgRYT9U+ifxEk323SDVe/wl4oD6Hhqb2MZUzBGRXUu/2DfuZQsVN8kTlLg8jZro
s5/V/brRB+Tz94fUEOTYu24rdFsMJ7oVCAMTydnEQBy+mE/2JJ5tYTL/XAYgmakG
TRvTe+Agdn4OGlsOm6egk4qVQN66voVWvuevRnjLS+6MVnQs4Mcy5MWlmWMrUKbg
Gxdv3obsNkOUg567jsrcflRu01yAaWRTz2fxYFIt3IvvNW522QEmzdfeVHGHhNXp
+IJaqNUjJJapgSHzRRGUEV+Fz3rmkOgy9sieG2XHn7EqTUa+m9C52bQ3yv16FXxo
wSTCmUqmeHGqBsVvwIK2FI9p8EkbPF37172xWKQdmSWaNYwzLGBPIeZ+ebgLmicN
9i1w4FNpFT+6tZt1eBRIAlnnPOOYK5DH7SWDksM0Wu1dkg1fY+t8/8KUokxB8z1T
PvyljO7LASzy/jVyNbGn34rZXz7oYC4zvWb2JldfFP0R3SUrzRivMTEN5GX50+lS
vF8jFEWVflusuonU+UBLf80cF6CimpaRfbdFNkhEPREKJTJiW+70ORUmqM02/Md0
oir9cv6IQdRTTKvjbskzu5mwiKEpDv+LOPt4nZAWM986DAde73ebYP07F4R7BK0L
fdL0KMmRY91GxXZQzdci3keYqJrdg92Js6c0ct4ZcQZEKVEcgwBbYtyd5BVmeKsu
p1pCPagDwpB5cEIr2vxz/AaMkFa6impO8wZnua9A6WReSB5nQ4UzkXF32aDy95XX
KD31d/bZV2FM9/n/azuwcFNRlAE6A03A9l3XbJd6Ts7ORiJNqzjbKm/VM9ZOMfmd
x8LdUJsdo8V/c/BDv5HpGWmjHgfL9QI8A+XZE/LPZjtiITPkYF04gNoeK9GqlV6U
ueXmGOLTrZlWkcaVDt9Rt8pMwkr9ZzRLOI+Nrh4VpMd0+eBXqGQSaJBLn/DqQcOv
SG+TOjD/vDo2CXjqb79EysOSz4EPvsgxHGmg7uw9lyh/Lj3HCLzzlx55/ocpAdUf
CEIeGpyUh9XWH+FiRH9whvQsodZVcyPYsC4TMyj2sL6vwRAscQM5rlf7Ja1m+0TY
Z7opbM5BNfc3702R0pRtteXPsG6y1qluqmKV0XD6CFmGCHZvzgasQa8yZ7ytZBcP
vK8KFchVA6FirwWgYCvz1I1LL9zeAFBCC/tLDrm0obVqcoOiyCQAGK0aBRzMLW+l
p6ca3/t8YkoBO1yeMsKwJW6Wcvl2GnIcHwHQuJ+ELXbdVn56GRptYF7Hw3/eT+R2
pYSFhL7CGfYpd7bAXMgaIDajeWWDFV2d909Hm/3o2a5OQxoF0TGDKdZnyfxqYnej
wF7Kzly4Vdamz7W/rjMLXeTe/OzGbxR1pdaONh3PhZ2B9BH23IByOquOMy5/gkW2
a9sL1entk89i1PA57onvY7SRxsrcy4/J5PDNgfa1yhAtpG1KeEmkkgYb4NTPhZy0
RS/GPGLw6vjzuVvXMQbG1xmsxUDcPytlSXoACg10wgiAonQdAyKultDiiBniSoCG
QU1OhreNna83JUWnPF9nrplzAmT5oEbLSywTZZ1/BRH4xeBOfqH84P4FZ+j6pWVw
oVUBVlBjpY5LQ/vIA0iRHgA6KXahrUQrjXQv+MjYDhDIWibV+HkzWAfuB01ijgLm
16KSrhTX0YhktOqujpr80scLyG3ngefLR5rD95BOygknGep0TC3UyViL/y1AINFN
7DEzMVsvdj5IWACwuVl9KWsZ5U0brv9VNPQ4+ijeYl1FAD3M96QQt4Dx4AeSNBZf
c6eJt8tZWWOWdm8wMcmKDpqv9dEGLyN8/Y5Jl3wMCddryUoeAtwYBfFmy5EG6EAU
7EAOb5MvXGKhaGoTIyV32+HKovGHBKwYm5gHWDL2kB8R7JxM9oAqUQfaHoddHRoM
YAiPSXm1JdUFaifJM3uSA3fgHWcvc1hIaDAlW818/Oh0I+p3zteSV2ZhYU4BQGCS
15iQz0sqi47Qhjoy/n1kntzosWSBDdhSL7B/Gkh/umlj8E40gFr/z91qnNSijZh0
fO1FFGpXTCdCBSuZx2JHWryWxhj29ZRXHY4t2nHleudIXD3RCvxaPBso3TLqlqfI
mBNz9XABhmZBOjCdPje3lJ/heiLbhByMj1C94deaoLIfrREZgYk64dOC+EzD/S11
I2jUuaphQB/lj24khXmHz30u2RCaASWi3PymoxTc0sJYrwNqNAnqXaV9KSYrvtYR
eALryI3qTuaDLmy/dr7BdqzNxE0477mZManm9BPNpOModSGFmdraxi1AqN2TKcEb
bs6QTMGndZpXFo33Kr1liiI9ikWhLR+qM0I8p+gomhEbNyd1D45naI+NI6zYN+ws
qctsEaLITeJkuJ+Y0B9ebgOlOeYwFJft0F2OSx/Jyusz6P5E1JbOv4Tm2CiveeoJ
sJmySwfb3g7/V9VuTx4y6mhjTLC/iL/a6bZegEt053JrQeK1gVbPBAecFGGysBQC
f4gVyfWuSjBdYlK45NR8AsviUC4Tep2YGC7C2IRxSLpUdd1WO1cj0J9KEbtcWyhG
9gp005XtJ+4E0IrB1WljoQNGHIm8PPDk57ismRtPzZ/J8olt6QV6I87zpncpVCK/
nuVikd64idcrYDLQGmG2zJSbbbbJh21JIFpHL5ZotCJKhlBkl5PQc5Yh9W1+7CjZ
1d6Bvs2CL2nStjCiaG0J23BsTxiUWZHr/4tGVEbJu5Oc+BpG5AniwaY1txCtTF/7
N6qYO/73u8ORjpl6D7xg5t2anmvHKBMbWN2p0Q4UYo4hu8sjrYA3uT9m5xEwFT/M
J9irFxwDRwqApa7Tzv7N8y93hdL6xaCwOn9hIMY270haeG+3M7s5OYGAYM+loShO
oxhx71L1+gFCC+2J/h8y0bDTDin8VGkIS3Mi2je1xONCXQM1va3bVs8QVXxITkNR
UO9P4EeACOffQEQhnCyV/rZDZwRuHK85GN/v0li5XU/cthA4qz2feskS4oLND2rQ
ay5+r3Y/pQuzOkmSTp6IH/dJa/HKI54DUV4GaZdReUE0wRCf1wWslP9qX3iGDxiF
dL20ND9qHlLutrwsvww+6hGtzIfbGdQN5Ur/Ap277ZI/1MuuXWPDI9kwD9ZhZkkc
OiFR/Y1SfdqWOCbNHhvcaxTK98HCgA5B5DTZ8ifCpztMWNIRy7mzfR7DHlxEoToj
6NR0Fm1+iLl4C+6mT5epqmZCRnLmJPaZY20ueL9WIw92kpsNAn6JeE8zoslmhOnL
WwXm6XV9v8rarudNPGFsOpdN3ff+dcUClXClM8yFJj0+wQQsJ3mBI90zx8/BJIla
ZeNNcCNN1d+5N29tsevD4u0SgTIGgjttrhFYbe1N51NXeMnPr3nE6N/moliKcYY6
1VlERszwyEQIQsIEtyh4jPG8eS9Syk868TfQ8p2TOEoTubDbIZfLhjJ++9I65LZd
E8kBBTRGCLLs6NPX7PnN/ULxIvPghQUp42AsAJ/zmp4dfadl9kAmd3fS8MkutyAk
pN29CZPZDh0pu7n8BZXF1Zs0hk1rHT4xzXtz+UZmYtrR7QrXGDssJm50ImnYe1zL
foME4FTRs5Dz0e9zHEWXanSsq10NtKcnHps14tm9rz8luXTEC/Ih4Flc3P3zD/za
Yduy+96+EpA/HJkUWeeIVyfTQ2QxE1espqhH5dm7MXJltT71sHFmTkBHge9L36F1
Bbm6odpLuFlNEDnP/jd2/AztebDpwg8S2AutgJvRJEBVPwHwPH0BH/PYghGj4VcR
CZezMfXq3u3eoPrXGV8TLq1jV1Txicw0MhrjXDyzJJH8G7DwpMmcnpNro7uX2Mp6
Qob2K7aV8BRtPoF8OtsMLo+Po2ossckuLSXGB2TEPrAFyy4bhXn81sSDti1mVdE/
E0S3ZupvlIYrDaru0jAo6a2oF0daRBktG1qHiMLIPEiyEZxA49HX7mZm3b+U740l
QEON1fSTPRzrMkHqnkvjKcjmANWCk1n3b2lbAzJMN4Ev7gnUoJbOQAz9iNuB+yXV
YnC8IExoKO2pgUCh8INMfvk8W3MO4fRRgHrKL8ctRInYJOU2kT/aJujavqPDzWbW
WCS4xc1xTueQYEctPU8KiWTh8u1GH8rOohX7pIjmLIFa9ly1xYC1wR+JKgg4rqz0
L0MQ55DLUhuKfe3D0SGkZ7cjNXq0f+WXsO6bzkl1Ujv+ApXVjyhTxN8JiowV6gJ5
OjWXloEov+BU3AKmdY14UrHu7kMTTj343n/JVuYgy1JHu4ywKLsLLBgF+Q+qgLsW
ruFkmlJBltf+Atl1G/Inu+XOJGL7n9mGamTpkFQHEIVg2Tat800rKN5jAsiRFMfs
LJulwxWH40uPNQZaTIJkrsy9/uquzrpqQkUj9P/Db87ZmjZOzfWQlxcdMRvrZUaf
Lt8ZPwk+buObRq3pFAvkmrAXilQG8km5LyRVAxuNTdyMt9XR5XtnGsfSXVPFuOhI
qvNTZpArDUKvKNVLLirMd0fkDYEo93RsxqpUuO7G4eDL7sIipl3nhZdy9Jg2q7kX
QDo/OHFV0DHK2rfIoRdtOf3kSduLbY+Zmq5+WywXPsm+M8xszhfBDQrRf36aH5cy
U1vC/eM/c0OQUSRULqZ1PfW9YW0cjbc4Y/mtdrgSJ81IZJKAvF7khzCb1VXUSNX5
9zJB1v97LbJfIA3Ew4rk/KtxuJD6CyjHaJeQeLggAyQ0VN1hZaOrRhoJGOmLvdz8
Mjg+Alu927vrr1o15Axr8sDH8Q5fK7yIOHlIJfLSIbtYo68bY4DhEgbz3+q3fzNE
cS2RLTCU97mrGm/CWyKpRGLVE1qCzKnmmjjzWPdeNCAX5OIhc2EpXWqBEoW1p7UO
2MhoOc09LDop1GIXvavHaTEqNiOMy9X7p5QryuOfbaq5TNcBOJYIpaQHZnYKaFnh
y5v5rzPwhaFjG85mYMvpy5sQdyGF1vpXyo+qRk5a1dswaFW+X8MCT97gMiznaYc1
K27SjTZsKI/9PODx1/jljYti9X+hB7Ly5AJI7KrzRKqqiNNADc70aoiFZytB/0cr
dxHtlPVgWWGQXbUIKccdYP05F8rug6maIWBznemeOyzmqQOVEqH1pZOGNdvHmbbH
dLbX1t6fIhyFQF56lVMb/CusC3WzFm5oNAjLWdbZEzq7S1UuigkSOc2CokIvb8Nu
pT11kUKW80rIF8kq/HXHN7I30LjIEqCuqdFTQStbq8tDLuM94q7ReeGmMgRskDoy
hM9fIUwViyxs7n0ZXoCPjD5rDU4vbMzSYVMJA/tKMm1Y8EhaCbam819tHZedPKz3
fVBaAdD4Qq5iBUJcrAiwfeA2raBlNkn7Q+OWUFr3bAtEu+d0kLopMeQc6BBybjFH
S/G8SAqnCIlqpvpCmhykPsJjLmBQo0aUSlzeOMtoemW7griEoIT9vgMKH0y2zK8k
ZiHrWVT3fT5pcY5jOC58Na14/4jgRU2Gqr7srGp480WpPpmAYqRTNpMHxiglTj6i
k1OSpPww/YDuTUWYCULnr9KT4fNVpzr3bB1zQBWrRiuKZkwRR6yQ6lPWqQMgdanJ
suc/cZi0KTtdSJDst3b4ZvnfwmkxHm+eN8SyzWnSmzQmGs0Zic+D5J5O95m/2qjZ
0lXqhGVydIf3y/iEA9zY+gBhEMLeBaezcwg/rUMIncO5BKMFVw1t65bZNJg9QD/d
G9Uqjmo8ImMqChlyKB+np6RLmt0gTBX9JuzpfdYlw8YBh7j2g1fv+VoWdFBi6kFl
dsik4SNrFx0bppKpQa0AiejO/aTr+SQn9mTspZechUdOakiPsVD9mAn3XoLfjHKj
jvEJ5TE3/MdqKYzutMYCIZaIVbpwwWgAdhH0n/LUGPEU6quFo94ElK6pZ2qTqHsh
1aW5pn5PpmSOf1lJDG0zsw9u6nzGzb9PpbygPGbdqMjIctmdgJGMsvCFAs+JSa+1
WZKeYtCSJCxxDzYLi+cFiP12gMMuOL+SAb+AEESNPHZiysJfAeiaUi7jzOZMw12O
BUDk6Muf8g3gCD90twAkD7zTUp+9356Nh2/9oTFY7tJpqsblHKaEIlpiCEMro1Fe
sUmfzdZwm28eVuFkxEwlWR/JRI+38FuNn13rwl65s3PUgvLPJhkyFfh3GkrJBoqX
kPG8DLadWH4ATPwDkQIw8yBmxazQ79qjklG7Nh0SVRs9/epDUT0/Iux3vNt5dekS
dyo0fkfIJ/Iy4sMR90nR+oZJiRRm9i4mwhLoduU+FA5Q+m+RoC8RExYvyPTwk2YA
CW6ZZzPidYVBQu0iAz9GGzXl1CdayKvjALhqrSEMjYdT68dLZu0Pme7TCEFN9oiC
9Exp20kBEl14qhtzO7rYsOIyR/EBqC/ZeW+OelTojtMExoQBQplCRbLjO361FfsW
x2gfQTJrem//RGWeVXzbvXheG5gTu5SN27wCvYlm1fHasWwoMsCuZv7dk+t3LkUG
1tMqzdu5H10t8gDr4sz1kdo4+glx5icUVTf0KUNg5HE0gIaE0GyGT0mhrKXqev0/
+Y3PKsmQ6P9F6TU8nlRYqD7+zBKnM+Lq24kM5YDZFsQVsoCI6OoAvVDd8ZveD2Br
cpqp5eVOdNm4CAPBOQTT7vhc/UkJhJHV4cabMOkJHHJLW8cOVmPw4DQOhJeIPLcJ
azn++UARUn4Ae3/qyi/iQj5Ubs5aa24UMiqXRvL1zxRm1SW+hv0ujMZP/47ObhTg
4B512dff3y6ecqt/3kDEbV8ZlPwxyaZ9EmT1b3NLI8suMKtkbn+RbltWbwL8U5hq
rJt/zdgE3HgxBARcCTb6n4Fur4p/gmKD1WOMuixtSoEmMFmchW1VfbKrtHSlGMJb
IJ+T9uUacuyojsW3k4P7mvn/oZbyF6B1El1lWc70A15hwl9+iT3vKVYvGZPkC6Fe
yMq2+J3ope2bYS5VnVUSSwe3EYRaf/xKpX1jChwFRuDoZKsaZcXm0D1ZAiDNWy6S
gHyD/K7HJ4u+uK+wwlhq3TRWgHxqIFihOyKXcC/sykn4BXqSQHOsYu3gira5ADYt
a8kavnRc+UZr2rPzVvkOVdai8ddUln7fYGGMzYFt0jWnnBGY+byZhU8wvsts3MV6
sk4AYhLUbG1tHoAUA8iF2+el0FwpBk/y1pFUv1TCwS96BF0xlLdYKM+ZPGeQgkTY
5lKgkylaNAA5SsvSWOS7wN/aJPPlEJGY5xmLCXFgEcMMMHr6zrrb0sTmLo/f6xOQ
eAowovF3Q4I//qMNWU+qZNea//Brq+MHc1FGMNT3Kcmo0BbklZjaFrAluGmc3oKt
S9ACJU1hfr/dp5yH3xWds7VIaX00YvblsCAmJPDgld3mO3JHXl6dk9jRFD1tj5nD
KQNFD/9HCZmUqaqtRsTsgCH5Zjp1ETaKyeJ3o8qMr9bfQRU4fzjnVoRpcNBOvvyy
z6TdzNRZvR0qt+EsDkI3ZevFgkWEB4kmrz0vle96BLmFbzI2JjiSFZeV+4jI2sy1
5+7jVqYCcdTPuJ1yuxAjY8xxTS1NR37vc6g6cv82QejpdiyxUYdoXoQFrd/oE13M
y2rq/AVaqeHq2802m+K3+G31A+7Nsvrc45grKImvHdJO8CYn5Dyvb/PhAFkIObSS
HjAXhTBuxdqmYeDt94HG6plSr1d/u7vU8qrm5RlMgwnGUHxdTeJ/hl6g4pqmh5cR
TAaU/0+bFrGb4JPCW25etuo6EzxQQttMFx+S0U/JeEsFB71W9XgKme+7KQTDzTsq
bknCmdQB1IDcGnJPyxoJ9HsgdnCtnnAPc15q5PvSsD76WI2TtuE7FvbmEV6cuX36
ZtdBSDTEf65z/GHZm1A+j/MSEGCM/SRFf6YZzHXOwcVpKsr2RPfuP9Z01/asVtRY
9S09DRmU4KbMJLfhYjNBe46zWsKtY287VgUKBAhFoViGSSN7CBMFu2ePZLisRGdZ
fSjGwQHzsgGPKBNWZvhYBi7DWVEjaTB1iMy8gX3iQXMEMZKkCaGQS+HNGOr4njEJ
leTXOX8EUL+TMp6d9Gq4S0+oxvLaE3gHGe7kdRKgBwJjzAvkOSv5cF2Hdw1s5w27
tymCcxeGS4IVTFIguhnP2UKZGhhDxiP8oAkJWYlqaUkwRGhtoerZ17TBhr/2nZOv
efdfqP0CHca8FTHvGHiAepMsRyisqRSy3k5Qe0bLrHjYtGVIMwivFSvv4MFJaK5J
3q2FxxhR1Ed+9vN72J8rhU6E15z93rEXLvjiqaa7uA7sFkAbHKROZtJ4Dpzpu8mc
u4588rENMcF5bUdTdrHVSycKwuXZrbOsDcsb/EYMTpZ3vUv/Pgj2cg3pmljzvT1j
4O328Ji4b1tSIyQIbiZVv1NZVtPCYxLx+W8SpetPnP30bhfwBI/Wf7p5hQVdYDUZ
EeVz0l96x1Fr0LO0wyVyZEcEofF9no2p39Ri1HLmNCQMddkGEyRCSDDoY8m3CQYc
LQzGGXCVrpjaMUgx1PcWnseHclEWLuFzNs4HknD+8PjFEt8jGjS6JCqf67sv8gzb
HA2Z5PuSlKKhMLDp4AgtLAj4JYbghKoAaP249adoxMeLHHPL4iIkhrG4Z8p2zH2P
RjMWyGihUvZJkPsx0h0CUU5kX3BKOqmSQ33KfW3cb+kyEul/EiYKVQb1ZRa1iqFj
50A+wiY+q6b3FkXxrrbgTJHQrvSlFnnkEuEysy3IHNKc6e8pQOdM7os8TCk2PPdy
aUpqIR4NIgOfjCJe/UsrY0PzTlpJjYPNMV03vap4Av0oCQ2CpaF3ArqYaRwpE8f/
jh2CknDYBtv/KYDBhx5ugjvBWMtEtUfsA5oOnf1naXNxRCikZZiegyM2MkbKpLqf
xC6Ypl8Ko/UB0e0wWNIMzMtgT4qyeS/soeS34KwJcoKoI0fbXZuv7beCW+rFA1xQ
+Rg4wVoohXyhT0pCXOvTuVfBGBBgIU/XcGd76d8xsNnVWHjwpHOduhl/qKDgBITF
lFE9mspdbG4xnusVWm6OnJ7cGkDdcQMTn4et7cYc2VjbTq+HM1d6G7YZAmi7pGir
sb615LwpXK0ylHSntfpS1UygMNoMzebLa0whZPTf0FuO2ukP7suzlWmETsQvvsNd
WbcCDi00t0Wg2dZaq9mxi3RXf48Qom/ezBUOuFRptubpKTmNx8V7rWsUA8UtZ3IN
3AHG4u4zp1XTRsJlF7KjqziCkvsR9nTw/kNnKSnrx7YPhB5euqhLIx/B+yNS6/Uf
xUIe8UqT/+460cYrGU66TV2bJnX7Sn7EmJifAt50cW1Uxw4rVAYhW5guZgfcoYWY
q4ZFfgIKmaIMO/234dAwy4/I3Swa86T52W9w6VInzYghveL3J9Vqd30bVUvsKQWD
sigIZ86kjRHy2xCnMuyYFBkGVQr+mmhgk2BBlipmUXuC4CqM3uNZV5w9hg/A5lAw
/GD+Gi36UAZT5HwT/IJCK/3XXsBhf2xceDMmWFk2LwMSqPA80x+pK3Kl/gFCNf3t
y96YcFx1Rh/C3WtaYz56tBfAnTfZPi5oU5YkvM2zbfmKZdkImK3VBjDP/9Z5V+6p
Ri0+Yjjgfw3AFGN+Qy7IzCNY+t53bwEqQOIS6F0rxkNCH8kpVe8MFDJK0u32mSQN
Xy/guc1/kmx+2cZhy7E2yYjyhmHU0kXg1IqwvpRI3BbSmQlJujNZOdogFZ1a+Nca
Kct9PQ6FNVDmOOGs4l9YMXr8Sg7O4rd6nJi4wSC62ur6doloTg/K4ORk4kSCSU/w
d5ieFBzuVNXZWcuz69lKc4ircuu1VqZYTnUuMzHvHWnoAtxOBpr8BSgjbv9lwQBB
Axe8O22xxbQF0HAB5y+2mzsbFCRIil35JHdOSaZ3exDS8f6jMlMp1jlDPLx8tJpi
KyPLJE8aqCkSUlR40BXsz6U5NiDpPA4H6/NNXHYt3Dzx3IG4i5W0Qz/ZnT/uMj56
xPUGygJtMel0iHxEY6FW6Vvomrw/N4iBHuCQ66Bv9AsG4pL/cRoyLELFY//spzXT
n7sRGTX9zm3/bUGykHVTzezh1h9TJKIrUTjy2hmHoJz/oAlfICZP688hM6z2x70s
H0v+ZpJFE2XqUsCbwQOm0jGODq2h/1vGoun4d53uVfIzZ76bQPiMYILb/HGuklAx
3mM+ed945ryww7/CQMTM8YUmb6Gi+eCRY83go76aM1+UiWod1aQSSAxt/F1jFKb3
ymFCDZgl4kIGLyecfw8ipdRqG1HHyMFhOki2D2KZ1qGCKe2uNPGort8d5OZDcm87
4NjCkqYIqe2TdXkrR8wnpX+GhTYx/6kgLReiz41wgitm6Vqq4wMJtWCz+HoOlk0Z
eSIkZAMZs0sjUuzTi3vAHj3RLUXNRSUkXCVn9LMdUddb26v/s95rCRwaFXaW5bfS
b9RaYFPL0FuIawTj8n5TTiinXp089aHUe0g20WhEM9ay/hzI6FebuZKug7d3l17Q
U52JGJM/kpRDdmd3Hks7sPwdh4BPj71UJ/JWpNPcvbziMh+IVRt5lQz62eMdTReL
i3GNk4UQ/F5QuzqVOM2AvroZRvdv/7cX8m/a2plxwgKoqAqxRgNFkYJH7ouuaVdY
imwez+unXfHaxMOGtbeGWjEUm04M1Nv69Q1+4P3DNfbls2fAMaojXXSPI027qSw6
`protect END_PROTECTED

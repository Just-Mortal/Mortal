`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BX9EM4ZVkKp3etZSfnzybcDLlGwe27Smi+2xYNEJrIZ1mY/rlVn6hWk57A49J70Q
zK2ENPnmlhPcywMcMhSFcAPBHqkyhy7diqxecK/d66YexcIGx9Cc5jGFY8gZF2N8
eZ7RV+xsfXln2deXPkHg9EhlnqPBDqYdaIgamlrUtBlXeSHoVDD6nPzrrQKxspbz
d+8yfqUzwMTO83ssikL/E5EgJPBJACEWi7pJwg+0NVOUs6zVcAofDwHEuWTA/uqC
2LcQytBPu5SAdqA42JTsfm3p2HBGyYnXalbrXEd/pdb2P3DgG9xy0n/Wq1CVrvd4
4aQzG3iISa/oI7L3MzZNWwCLEbdo0+P8VUF+H1wSiw8o/KeI2uCOGZfcBufCK9wq
1RnnUrShya37Gx0kfwGQw1ttrBgUwzqNFeEWQdudHOiV6fEJdJ5z2QSizj026iwA
jnVMn5lphTOkpOc2P/RQZwcda1EmjyOjOQMRcXCLAB+2WAOMOzC1/+Z+DwPIy9rY
clzmxgK4TSLq14nl9IgYbMUcsP2SNn0gtYO3Cn5odr6IqozbzQcSDqG6EW98ys7H
Z3hChKcBlFjVxE/2+b2ZfhU1XLeG1Ci7JHSq1SVWpZ1osDTW9vs/656U6znL4+d4
cbRgMKqDobkVI3IIFvklzLHMO5jwGrRiKR28kie5zzgy0vZxWrrHzuFZ0zumUWRD
TmhG5u+K/NKMpVNAPf7zqvJdDPBu/JYGrpQ6cuWzXY5SFFeUg42x70Lk+3YWFq5q
d/zxTXmF8Z2cxZWhImQj6wSMVg7GM3ZMbY/a8s41+klu4Rjcxo2SRl9kfhx+54zP
SrJFp4Gi/oWDxy9IA+gGM7DWjzHYm2jUJiaYnnsIStH677XeBC0FRaJVTrRqiCGR
i+33ZsT/aFtrerlq8FnEqCQu9ECydewhQbSExocObQa6mW1jD7pMO4A3Jjp4AIQl
Ok/nU/Yltrw5qTPDd3DT5wziVH1ZLStGgI/vRA4i45K1a4kC6L41Z6xFy0h7yOGL
6e1D7zV0t/4oi1y9rX2ZMPApEyXc2zJe9a6mic3xlfW63xX+LfeSsm+rSegJ7lm2
ZrF/rdpzdJh2pUsouKcUy2ZQsomtuVU46TY0HftwfN3br3RTdvwCPEOiEt7LL3/2
tZ/Hf3gEqyYGxfWcqZEFSNHejL5QCBbIUwQBs5iHj0Ly3si2ebTBirt3Taxo0hvj
ycPB6KVKeU545JeRAxfXHz6M8B6co0dYGOmExCOgScO1NmvZxpusDcWhdRnkwIGa
Tzi28bK1q9oLQzoyIVi47ChxeDGsggTjs3hD9me01p3OoOtr6ud6muY3yX4976dt
f4z7TShFdfCpbDFt46vajdI91mTUonH3PSeyzm2uCnKgMvQ/ubmNoL5CiJiP/hCF
hO+X7216XOpxU/uH4xX9y3t/A7BBOcOD8fryfzOkCqq9pU39wGN/XXCfgpw2Y3YE
tAfslxrTLs9hf0sBH6zgTw4dliIX8wFlb+BTWuBOlTIatQ6wIahaGkzDBbKDwLi9
teCLrt98PVbiaCy0NW4+LID8itimoicIA+pdSzXa8o7RxZY3qThmiLcf10oCYiHR
/vX0EsNcwOxmIywqzNqsnVReXnBsGIwjraH6/tOkkArbT2aFVFDi69uq5AXvYCXG
ZPgJ2RhFqkLnEV4UdlgP6ThrsYs521Sqvgmo0bIdSYSdUh1YEDyua/J7atkq+Rz+
WZs7cyAAFg2dE3ibAEnlZjd+gzQX0GoZRKq3qvsW46qgOJE3Ki2C/Fz8OU0h3yE4
kfp6QkBn2tLSQvpV+Z0XQ/bWudR0P2CmxYrlJBh3sTh9oD4InAVLAsaDAXqiaaft
puEH6wNqC3d6fS/ITwZ7NDBdJCr7886Mafb6Zl2El06R+nZ9XTwZXy8h0cSzTxIm
eezuPCvH08YpDa3ynvQc5J7Ml5el03Ry8ft2GLg7PcoHhLEUEZ+thkP3HYrvf9sq
y1g0H8K1tZ3IKnWiklnb8NCmOPnj1DH8NeYpylofJxpT5Vh3UfgMI7gQB7ZAxYSG
5HZXODBNBPixAasTBH7CMuKAOxk6yx70f+xR/QnvRRzJSGgEOfihRMnIIjskWarG
FKTkkjKWLyxjgfIpbEezYYDmCsB53vdHLPT/uVO0gjHFAxRmVBUoVYDl7ECReU6r
kkRK1oO7fiAckElm8IhMjMUD39dLtMplogM7JfrD/DVfqXI1s7msJbC+eo8QvUwT
T2XdqpOjEd0BXzK8wSfRv1mvixpNPdAbpL1WT6jlckO5yhuHxpIwkkyLanB7LB+i
KIxF/rRGnCfUngVxwHDW4E9u5aH1SB9g6CmaggIFpbXDRir0tndT8hgE7FWIOt22
rZ2QTV5W7hmgPhkLZZua2WgcLZK5fCiR6Zya1jmYuCzijZFsZdLuw+6UtPmZF9RV
1kh6EJiFeYj/sPX9LMXDXcH/KQ+fDk/7M/5CTCl9pt/LBl6UjSAE7zBm0W4BseI7
b17Jqxjtw9MqvfMXypgRrGnx9YXzFWuOOFN98DAe85+iQy4pSuCerp85eJQkOLvM
g0NPf2dDWBFBbz75Q+6/dD+xonk8WLG6vDruXsLppv7kdTm1oTeA+9fm4PBT84cc
9pAc0P8wFqTxNHTzS5dNJWAxiaUdXclxuU1nT7mLxx9XnJB9OMnzbtjUJyxWxU7A
s/Q0ELJ0kWDgvL4Zrk5ywCTxijvIe2H2/iXTePjj+KdWpeg5gTBMD9XTicTbJp47
qNrtLTUQhtmEDl5ztOTjUjMyOM4PCVYuXTxF94I/0Vf7ZU18hCqsLHamlBwjlf1E
4ajfbFYwUfAXUBtkhb91/h+6I56PpRwzn73+tIm+dcbNrPThjK4poXJwKMQesz6a
wSHHpKzKt/Mrx8OvHERql3xcd2mO8swrDGX+be7qImhysgQhKNIho+OU8KxZyVV4
BDsVFUKo9lcRoRG1RMQFWjhdat8lFi0rrF3ICZZl779dvWY8BVbJeElheNdLISrR
d4E/ybLeUHHAw4sCsHUMG9/sxtbsc78qItjSlEbzat9UzA72iuL7QLul1DoCiabm
pBjBwqepi0/2KXsAi1EyQU6FonI62Km8SZDqCthcSAdc4w2dvKYGUJqT/I2pZ+f+
VkkccEv0zzFY7f3G9Wn3BVnwnCoplEFzKIRFR5wB4kqqVPk3bLQvz5gUym97oWnN
MtUv3BjKGU+F+7lyhlE5oGGhW0PD3W06ypCUtek8W1zK9n4PuDaCW6qShYWjjccx
o/KHYRf5AwsQvhdkD+2PJYvj8Djg7/OvjCBGH7Vstd+wx7jvEm8HXHnu3KgbalkJ
L6UWSc/FeVEDUDcc5eeCCZhXcSI3zjZ2cE1ELugS1LYiaSmpNg59ZCzQ2tMBgTvD
tYFhgjfYE2jTGJC4nK3izinHHuCKXKgP6YC/niq7+qCgX1WiD1tXwNqn1bL1qlIe
XaGAkSNbTSr1IT7/1LckCHnSUkU1lNRo0h0kSsDXzTtU1XIPKKDWFb1dusIgZpfU
Mzhccx3lOFkmjscFvySR+fo5WhzSMlJlhD28KCs0TnB7JFTl8QHva+5oFc826l6k
KWqaKysne9JqYVNhQJPlaiarEXORxgXbdJE8Skzl5D+M7957xz4BZ+OBqvQAcGDH
HSDGDy3ddhxrhwOb8ffRDhYUVNlBonwZ8W2hot3/pcWRnoU+WFSkCa0zzgTLKmkB
p+20WfTszCOlbWS9jhMvr2c+jNZRwnRw/GzXYeu/yRNPPhSzSaovvx9gp+KPn8vX
quATKNoSqYXu7/KQyzEDUjr8K6/7AXg+Pro+8ssDeNHeYI/Uwjcd3SXUsIlDYbk+
2/doW9T9MatwPgfSfm3Msk1IWANt2ktsvLHP0TFpNl45bMUdJlKCfo49N9hSzpTq
7hSC6/6dkMLARGDw1JzOVdi82qdhIO8xKZquK9GE4T7eUDlR4+pWaOyv9f0FquCK
L1hkWVndzVDSzx2Lq9dvTVS8ryrvKtypjr/G+oqwbJuaeFHQ1GOL1qAiatna5K8r
wt1dv/hs2cFJj5Z4FEfuktneh9ho4VBP64voKTop9MllAobzULMZQxjyG+uYWZTb
Kvj59LhM7F/joNfUDFfxTkAii5Id4uTzMyAWGlGWrbWwOuIT0YY/OxoEQVXK3KKy
pixWtykB3BM1PpCybv+u86S8TAd6j70fyWjBy7aakgYArjkMe0jcInIAVJzvu6Wg
qmZ/pRIaQelDuv+o+Qu4vL9CIFiM1tpMSsoS46B3IRfrfsHFOJvd92QqNSEPr6EN
iC1bEChAJLj6eyEx61gqeHTtcKw0f3U98moW+1Zul+q6YTIURP+mxfjc8cojvIyE
wi5Bk4G77oFJHgmUEXkNtIM/SHQhqtITXq4ZdReFw11odhgSiM8XDHX8+RKB8SPL
WrpMV4sXOdkeLzo3JrxhBygksN7Kmzb3knO6mfEyZufbN1vJyFEljpe6nXK8itFo
lWacbHxGN2dfSsJ8JcmoygHRKjsYsHUqYqVWlEX6MH6VmLp9j3EhZHqxrl2lPpD+
GNpLxkEvgwe4iN8lC8sZYXnPUC1y5xlv1aE/nhKgFas6Om0WD3oPigTKvrX7M5j/
GuVflbtqcBWpOArDHNgz1VlU6vyfsmWS4b31fPmdA2tWi42L86aBZZV9XmIPEaJ4
zfpIlwx7XCBe6FABg8M/lj8d9Y1k1uj8UTr8LsShm/GvzsLGq3jfzJRXJi1U1UdZ
WsQ5/EWc25Ju8E9t4PnynOglyeE2m2dMfaL0kF5SaVWcbYGxwOK/+rdMFVWwnh25
onN0OAHoY8VWNp3bXeTkEtoLxc+dUB7ldThngn+ROgLDI98gxR8ZpwE2fshQXxJp
eALElSe1bwjvBcD+mYLyME4a1TMaMsA9uyWe+HeW8icOo2ED7km4OeIl/pat9FsV
rBA/xaLeyrdt3P9dXCqpK9FP8zStbEuZUkRAYDZ4Qir0+wUCZV+wn+krZYAV8uD0
GjMltK4aBjESZKnusrk/deidogUlrr7Th0KAIZsu8gMBHAW/cCdoVJqmdWeN9YKc
n8hlxrBACs4KE3EUSp6WaWr35kRJA0vPbfNcW6n1YNZL0anKho6c1xoH7DQVaZ67
nl/OZa6jYS9mNkT3TBkRWovoCDbkPm0JMzCQKcCA46Z/2wxrYrc9/dyvyTawr+AA
U3hqOVmgTDzWuyqcj9+8Yi97bXCqcqAgupnV70aqxYwyVgZkn4IXRwD4zf0N9IeL
8KuLPLPWc5ET6yQ78Al9h9w7m9SFX8t72QJsDGBe/JKe572TlILoVIzjpZCKj1rc
gZMN0auIdfonGpefAWDLz+ShzsrezrobjDqmEF6Rh9i7CU86mSdQXGQjjQ8GT2CK
cJiLri4Px9J0EiyfNIktES93KEdLAb1QEoP4ZFD0mwAEmZHblORBVR/Un+uM5eaA
FMa1PFDnKQgL4iSJ1Kc6FP259TP/kkbGmFne6vm9M+nkjk0w6azSBHeei9CD9XZK
EW7ETi975kwkAzTSWSItpWIEXAhvtK7gpf2v0omXLVqzFPrKDBPWb+BYG0FvKooA
kdY9mBCIDuUSYl0LyaAfRyczhHvfRUWUq7uRaOesmGAgXQgme4+bYl3z7P/ihgSg
MWYlSuzfcIaos4wk+JVUSm/MkDfq7r1Zjl3EynImqRPeprkHcziH7lt5/2LwJr0l
qJw1lHgFLnfyYpBSCjgp6//XWo+iIEuvVEuTrgnWztS/WFENSS7vD3b4TR/U0xXV
5ESoiinTD0kLEjhToegmymGiCbB7pLLm14MNh/vpcYd3ugAuW0mRx5DaVb6B/Vmd
3uas3OG3JqFu0GTwWsVx2KqnUR6hf2hVI5ayT/KMbHOEjRAEQysBtzJYYLx+C/GI
cwTGtwteTAm4P2yW10bLVDHx4f03+Rz1Dulr0Dw3yVAaQkO4zjsfISAaS8wOlRhy
bxIt+w3UhxoT2Eb8C45j7r82QNA0dS7MU7SP0LFeKxD1ZIks16vzQcOjyOlDfXoP
qQl9NiwX95zQsao+KH6WYziDqujcUu7xDNXFPVBTVDBxNTYJ3fkO6HwpsHG7qQvp
F5WqyOpqF8d0WbcJCSd0Sq/6I/2cqEhTRba7iyTFiRdqHzCooxT8Lke+ZhcrndrH
KCOiL6JP8DRWPRirVfWGaAzgur3yvEMjKTy4+hDeL1hKdQHfc4ryR/6z83YguIYm
5lqAFXiBygUs3YEddJe5R7/KeJcFWy4wnUYQqEWHVm3d55ikBrrXsPbzqTqjvlQj
wkHIdsfum98LkKGpHfelfJ1rVJPB8gCl3VSOnQLUiXgkaXn+4Xe4RwL2Qf3Vu7lU
Fu9rCgnmPz9OsoCabl6YoyTvPHLx/IxONvPJx80A+knkZIiFfQd5biT8OkxHPFt6
MHnmm0ux/srkQ/YbTCM4XShzaAyR42eSIbkFEFi4KQLJBg1rD5E1wrMfkukv/IxF
sdqhGQdLEUMtyFBqsFfyQkQsnxFzR1XJKQYruqWdFwd8rXfe1/YOZI1Vfm++kClJ
b0BnjTPRjK0SAndTQG1KfVIbBZaNqNqM78QS5gNjmi+ON2ypY1va6RfeWrMgQGAG
uAp3EQ09s2PxAHBBPWQF33p6voTK2ZQPS64mIX+mkrO7kNj4fBzBVVW2imBr2Q3J
k9JV6kGyWbchudcCJmzge1MPTlmn6BBRBDNed3MxBrM1UObGpPXV4eg/nM6KAg1Y
Jk5Aw6z6aUtCnZp1Kl7J+Lhg3wPO9Mr6cXUJtAyb7ABUG3blRseJ+YCVDy2KmEKH
i2KS3AguNMAm9x6ivmHrWreQHrWvS92iBDj5hq3XLTv6kmiBHqNqPfAyEPqS5LT2
E4A0avdB3g08OVVQZOVfjiQv4XjLYtjLgk8/1Fu9znr0sj1xnzWjF05BHICUl3t2
N3qi4W1EIuaGLfh0vmtHLOfVXTMPNe0CHWu7aRlOehli4xS4Zp5cm+zD+lVd/lnz
XJ9UOQGpJF5ExurMxFkOAlq9WR8YhV2psyTJWgbcxcTagxdFWO1l/wzFuHqCOEdP
/uayM+pysL/2r0Zkd6cwla7audEYREno37mApJEVki6GS65gvRFb8Q5duM/Gvry6
ixzc2uiZfVcIPc95lvWkgIxkKKWlh2+ULGBybLbtpb3cQWPam8/kt/lo6iiD56Mk
Bh7uRYDbtowrVVcB+E7TkkoP9nUw5n8yvwFaVm6RxClV8axKoFnBkWNjj0E0mXPq
HVu57ukwEjNEUbrKg5h06oKErS71pKppjuN/uqPb58memX/rgkRPzdctTmOt8M3W
YuGDVvl3n4GzQQ62emARxbtMWt6gW3fGZKkOyOqNAjPRrL6tWT6Hs1ys4UTkroim
kfm1fIGxGc4aOlNEMozH5AdlrLlCW9/G6wPcuKTtRADcZaxzNwXaZHAQ8aY0NAUh
CLNgViHyd85eTEKcBRPl3xwBVL+IYfnARY0p74RxNvecrZYH0dT9GRYsgwaJ3xo6
VmqmuaIFHWI7hJ85hP7oHrnH2dW8pucQmWYjuQ7EoepwJ/L3MCgyvbw17xPww2Jc
ScoK1n+NCwI82mhVzoLWTUBB26PsKQF5CiJm1EQkq3iQMKTahsTK4t4bieTpKtJk
7NvqzrLbE2VSN6DM9Fn1TzABZGtGP3CrHNlSSIlM1dpBLflU6C8cV5+71nWBIcDa
SHUGZjHUE2rOBx5Dcp8v+/9MKbtjYTL2Aju7yugfSazotuC/ZcGZBrZm1r/ER8Mu
sBsmJe9gg+60CUY10YtfpGdVfEOotpwNdopVhOuzLXYIY6Nb3isN1qPJRTj3kOVT
nloIMtKfQXFU+0ve8bZFhOJH7sA9n/AbAEdRM1TshcaurVz2nku4kXqK/CDyFpKX
8amdzd8itARV+vFY3pfy70l0fn9ZZRbrCoCXOOt1nrlbrZUaorhtm+fPKz1GmnUS
u6DIr+j68uqOwxIGfDkpajShIQxeMmFyq704EUDMvE+QmLHWm9bRBcrSwj2Lwg9R
DbpULdEIn9fhtfC+JSEUQ46VHkFje+JAOtlSq5aTrNAGSH2TvppyqTZI0JShy9zU
be1ZBqujfDW+nxh/X3m/cKwMs+IgCYC7DTcdUAEpJIlKSngDR0qsDQDfwjgMl8ZQ
L29bty9rIannaVK9NF84pPzjSf6RpsbWkb/MqNqrxRMc/zieLAEIYK0IjMBtqP1i
w+zim6HmT+KeKW3KIW/GnUQCNLa0nJv0K/7ClrfIMdrPPti050IGywdAUOkJIVSv
Y8g2yFjkgQk4jvJ841AlSjyjiyolk6q1zFDzWQMrKDHn1okAQgPboLUzuMWyVyCS
hx2L9BrLgAi6lUu+Xr99nvhzgVKtO6lAzZjU9wx7+rvpKUAQLv/oTv+QvywOOzay
/D1YQE4GMrIlLM85E1A8rBqmbjcIgSEXJggHjbnJ6orgDrIZntUZziU7rD59nkAb
uvgOnrTc8NBQg1T+eGkgXz/9WDOkwVF1lOSKEd9MW7uiYaaNsVXZqz7VztmFNCVk
nGQTbCIt9x1ko2yrbD/Gg4YWBevCjq7jMrC/iSOh20bRKbgN4f2j31lbBzraAIFC
qamtjmztZwJGP+k3xXrYE26AODfV0L48RvNznzzyxJBIwUgwU4xdhSQ0ftYonvHX
7xp4HiQVVjz+nGLb3wfY/NNAxcAuzS8/+Fa6aqKyj+irvWjLKNLfJ9FzA2C0u5SG
BUA+D8Vs9HiyDYExAtsm6BUZFyFUX4ZgKZxXnv0PM623fkxV4smTbH6EJRNEzAof
8S9smmz/tTjAFXDhCmdMGnKAjU0mULwMAt6Mo1QQ3RS/56/GJHObLGkVN5a7Aa+f
ngfA/hbm2XrEaUDMzAv2jJAJo3oyV4DwmyyeAHhHQbbZszvFGzw4lG12KZCRRgtf
0NiU2QIb9O9BmlX318kjkifnwnD3qLfc30G488pheufpjXeYXv2sQAkrYhxdAtaI
s55LAa7BDky2pJXHXHeZiHgtpZxLV3J5SgAbzanDRDd6pozGaUmSN5E08ykNZFmO
Z5KWRxRjx/7m5r+rqUjPvcB6Zga7rHRlcez8v5maBu7QRN/sOEEF/e9QBnwouRiR
GJfzFjAamMCeznWyvZJX8hNdUVDjnbpfcjlba9s5gzMZBzf/hOHd+JLQ9JmtPBNS
8Lbxrh4jYpjeMM/X1kBsK0iX/Jo4gVf5phnF+Y3WoFDory34uL8UAt8r9Ul7WlFp
XgoRiFyxKUsic6MAqT9wymrYzUyrKH1QrnUYJrp6RR/QkVYQRPtNrmkD5HIB1czv
+dGWs4Plzt9TMBdQ60Q1u5RYJtdbvieLD8xi8C4DHKSbfgfVyMAuEc5uCqsTNuEH
p4AGHS0h0EPPGBBlJUZfiDpXCFfFqS/Xq36L5J/WFE3lJGGp3KP0bzv6bmwI5DvX
gAKwWHBg1fuIfDj/gBMCnKXQONI/Y9bPq1VuxaDkYLWgUHQviwc0NZ3HDJujZzBq
Mk7KYq089MRhuoUXbozhE9lxdmb5yxehPW0rtFoujOrh9sUitMqs1846h1bJfcdu
lSxrxQQolURWqEc+E5AgK4hdUJTUQmEAqZMv8tSg14eeCbvEOijgxs4yzPLhQ6YX
iUQgzTmrSNkxKgvGgxTaku1bR2/rf95NX5dXr9A7+tamqHMqgkg5GPJX42VMtndp
jkTZiqwgI8dLMXPoCcLYoN98Ivl/dseuFuhQWLK7gAHJvYxE9NqgvcPQXUW/CCHN
5RRwgB+wGeJfGiAvaz0VHKmixhwKoyHw0S70cEsB44+oVaZUlmBAd8rtENEufCbV
f2fEruzlc5d1/qEt/veOZXg1UPZSHCs/8k2QK/aXJA+QGup4FW37JqfjyMT69qxb
vYZFT1mc/cWiWmqWIVbnZB81aPqobEIkTWCcXnjIfet27RUeo7I9Sc+ChvZ96VKg
SqmF4h5crV0Yc1dXR6r8KsnbyMMD+DX87XIbWpM9g0emv/TDlyFQRvdM8xyZw5uA
POQoUwbqWKb7GqoFCYB7PfH8bd51dB/+cW/zhpIwvtqXaSxe29WWFLraR9dCsssD
3LCr5JMelETn8jAinYEp2gHh9Io4a0j04RcnVyKDVD29bT2Sb9YU4Yh8RjEzxIG4
0pzP1+7xJNNinXaIzor17Hx0Q87MZkGthZu5muYAulh3hQiewIzFiWif+jfVjeyS
SbLrJxvNfLcyL0ladfZoaYpyQlwif9t8+HZn8fFMuIx1De/iGk1ttsVKgiXqAGuh
NYGS6AQHGYcu+JdDQO/gHddOB47rlQSbxD22GBHtnigC9ulb/h3oFlYr0a2P+5y/
GMNhlbNt7fzdbMQSxUPhSsverMCoDduKP/CMlYp+iVuhCxhZwJtimdyNkiF9+WbY
1P+UyCXFR9uGSea/R0A4kw42B06SV+nsF/0glB6g5i48U6HcbKl0POFR0SXjNwMB
UvQEkmSYBfatXj9EMPJAl0xAykv/VmYTfu6dbSl8c8MJ/yNLyrZ5t5zmOW521mqc
IJAhyWlzWSJ6kwwoIg0wanIed40VG9LR6BC7KzVOkSMHPDMBeDFCm/lpMaedJbAH
vkfoxGAxJbHua4RoXUaVlScDJvsMGg4f8jVvJYZWOq+A70bXWvdorl7483/89lFH
9UILQ9Cu6UTEx4fUQOtgKL3tuQj9ac1S872420q3Au7Z3Hon/jIloGDRLf9ACznj
D/n/dfK9wtJCYNZlcjp/uByd/7daPzD5I1KUdaVQMVuGsmi7Kll1/mPrZfOmP8gI
rNXAYAJm8HNigjUyzdkOPYuuG7CHOIbe/X29+EkC0zrZ8NjkMmHeoUCIrXvLm9/n
17dEuw4FJ4mTcRn9kRgbGS0CtpWQNBvpJ8eyeJd1FaqqgzjzNXb384XByAdxprrU
ZRj+hDL8rGBE9eZ2l7WOoJYTsIdcCjQP8I6vYiWbaRVLjh5E/cjJhq7fe9P7fRSI
RfAX70CwEBPIZ5PP2kar6iBaZnFOi65u6yeF8mIDJ+3x/dwOay7jKKAsTkPEr9jB
zn0mKeNozAbpC6U7oCpX9v5NA/URByZxQTKdg35o8fenxoQIxutUASl3KGe/yQLb
6v2HWmhr2tMYdydSyGhkIJ3cmikG9XdgjTWkhtNX574NHBnv7b2PiEwIxMQlTPWO
76d6INcx7u1PjEngbs6Vk3n0FUQDnNHBcaue/BtslSTVtIaPX5rjCcFCBZ+cnNME
3OaQizbfilB+G5AThxyTvjIgCCgJsg94J73V5w4uMAoFHpaykF5zzW+1sPV56YM8
J8NVYI0vekVT0Ezq5o/mIdmA9G1n+b8I1NLInVBut68NrxNESl3bTHcJx0YWbvnV
4Z92SV8divrppsnHnNAhBvw1Cix7x3rBqzsEX+uiYfLXldCE+d8ROLETeuxpkao7
iDNihl3mBkiofarESIkHXAqR2RiXUpgqbZiAbpIG+xBTI75if5iTz5tq+8+raOe3
nOECzeVFJUZa0Xcnq7PY8JRjkpeOgm7VPXaOdc3qxaulzfiYifb2wxMjAnc0SKgF
yOaPcNhHtcuLRukTkYYuw7Z1g6fxQlN+jHof0RqYHd54CN0VtfR49jy8wRtbByuL
zx+QfbkUJpBYPPDjTn2Nu1fLeIAB+2H+B42QwRLP8Hg9W1BMLeyTHAR62x7Kzc9O
AxQD7NLUuG8sq16NBZ/QrElNTH1266FPEk4fBW3XLd/yT55mmF23vdCCGIYytpR9
6bViM100NlRT4Y3IQt3iub2zYoi3WoiKRBBV/KN0Ac4hePbERcXoW74JPPKAOK3n
YP+syXUiSvuiK8TtzuAFNtc6hL7AogPI3UOMw76fDCDkYsqafng0+Jfl/pNDL5Z5
vOLAdTv4q1++G7Zi2uZce8S4nGQifwhuSRAFzU5qhNykR99sd8SODCv0mpOzNO1t
YDzsyjDmvwrE1cnt3tIZ24Sb2LuSQeIoMDBm2xCUYTVh742jREPKQfjiY1lPE+Yo
ydQvxQZCB45O6EvBtq2usJ4Q4FvsZ2uCcHVerCOaFJ8QsSOsloq5qph29/QMHNGy
MLRCiIHwerxr5fcarq1laDYM4KZKvX3DtWcf3jGORGK0zaAtbR4Iwo5NmzXkySFf
innuqY38AMZTN12lgE2Mup8Zvf7XKojn53qaRwpGtFDdaBke8YT5GTyRBwJtD/sZ
/sPd5VvL3MUhDJCoF6z1CRSXjMUSnlqZTHpwbFviCK+nBAKXNfHoHD5pDc0niTPK
MPDBMTaDCEVw2Bk622Bh3kyAM8PaA2AyWLfDALzzXNZeyaei43LmaoKXRWVyscoz
hSzMOorPTpGE8kFeUHdUOQpOAjbRgFWCP/GqWu/4tkHAjtGu5yCLK8saDpe/xh0w
QVBlNllE5r5L1ep2tO5XM2eB1AtJMZrUFhdTHSiih8o/9SS878jElI+hMIvJ9tzs
CFNPYZFaWqc8mEKLEolanIsaA5+Da6LSFjltQdsAYfvt3H+UmtLOe9k4VGojx2y8
U98lHkV1xuFKbXeme3almMqYnJc7FRDF1b93CdUqEKMw0Ci+TPMMiQEX/ZVOrFx6
uB9ntSvbYl8ij4t+EqsrcaUCa5GP1gSuZaDtjrBUda0ubx/3LYQbgwbfFzUyF7BU
XdphNII4UxGuc6XmEjgC9JB3jDCPA8Q0yANCVvNEGlJKnNPkYgT9z+H4ZWvqrKNc
lrFZR4gFyKEFBpntRj2jRRXw5Tp4Ut2z7wa2JrE1t1V6WmmhkWuU+iXSX6MjMvuP
/MjQqUn/m/yHcR4hjQIRnB79PumXLpIjouDKxDPWgKoKQkA3WOgPdZ2oCYkXnpcm
PpsUoZdiTJnuGYxWLum5L7JJlrCOouEEOwy3JG8w43CIhupNXWcQ3EjoGJsRz08S
IoySizqce7qUWW46KeXqP1OWLru7A0bZYfX/z5zNOUN+W9RwU1ceglJeNvAUD7Gb
qtJNwrXLxUt0UUJ2mtcAIQGG7RBh4vwP3VNiq6vvDquLjhMfhQmLrDDcmMudEdQd
m6g+d4zOvvvrTT6p42RsGVxU7HVoPDYg7H0PZw1wF1mVWzwwVyFxxL0S2oBbewul
65BoSp7Pir5UJFod2ANmxIlAiVmnZ3x1DapvwbX5YPjPGi5EEkRhTzMBp1i0BGkm
erPeXhx5Tr43brfJHt+wKgT5sYMwvGESl8bvXK+FulMCFQe54IlhY7aiEEbta6Lp
kJz+huqslEZNlURVR5DBFwwk+aeILJycCAHRkD68+pRbEIY4f7L6C06GfN+I8i50
mmbG+0kQlTGTUYJElxcK104T2hzyYoPNvF4E5LogGgdyHYvOpLMfUcPpjlLgVDCa
t69ronhZDoucfvei5Ygody6elhP4pvZxY6TLg4eTlaubYWK6oyeZpH2JnM7w2HyD
sDVV3tTjQW9d3K7UL2BY30qoP8cwS3mGv32PMDysEpOA2yOMsVfwhmv77mkBP1ci
DsF5EhwePweivEp3p8W+fKsYk6KwkCvFCrLcPMBvvjIjplXuPTcEVP2tcvLEZb2A
jJtbLtX2asjYp/mVPKzs8nqCIn4dA4tjJxLdOkT6j+yZBX2MFMB3wVcwYdSHXhC/
enl5JxnfC00TrZMgHJTyHhyV+/2KigCzrmjfY1At0FnU/G47owhNmfPkrfYvWQMT
VprWbPclX9M9o8TJMSBw1j+BKtxD+pejW4CndThqa1oglDKHx7nnTC8Z9VfBU3ob
IOdD9ZKVspG/n9l+gZVGkoBWYZEWfbZQ+NzowIkIpruJLZMYXdzUejFoo4A6Bbhr
PwGpeh3tnQaICFr6EdER6+d21msDDux4+YuSdJ7hm45/DuTRHfclk1rasMT/257l
1cmz7HrjARNZ/SVGnUGPeEM7NLNNUqfXCSPvFy+zZ/tHNVY0/mFdeUKSphkqmZRP
1jW6JVRxR5NPOY0DwK7/QVQk2e4e5iiD/tSApWb7nE20r8GpdIZEPxtkeIl9wJ3s
FxXysAwYff/W9j8wX8lhFWwcu86Q5rfHLp/PP8lhJt9fSdKWQJf8b0tyZA8w9Hlk
WOt1GQ2eFexX2R4im8DaTeFiJxwjYnC+mfR/cgM/05ESlpEjrpiGAlqTgIQtBU7k
48b6QrZ5aM4Ch7jhNWtxXogJZ4Qdt6sFnq59JY122DqqUNMYtwoIZqI53Btv0EkI
mtMg5mQtHETrkjT6ZnMDYKHobqFDeiBW5FI7/itY6uPcoFosw+nRmpAuhCkTg3n3
dYvBBU2X+P/XNmvuO7xXNbSX73aqvY62SDQSBb1lcISnaIc4EF22Wc70ZsjI7IRR
LQuqqkL9ryZw0oVwZ2iILgl/u4STSqsLc9733LOQoKpDlWXpNyb/gUCRaXFbpc3h
0CygjB1/US+ToHwTFQj2tHVDC0B1enZKjWJwtuszUoh7iXWs/8BHZWqGgnS8cMpi
ado3GJi0+hPehbPy2zWTcVl/mD9EgH7Ie1wvAhgPxs72JbB5ge3W/jW7oGb7W1gz
WK3V8PtB9dvgPVhtF2b63pZOw5IpydO4N3yPt32YemIqcV1G6RLJ9J3BCiWamJPp
w58qEtFB+gggTmz0MuOiGQ+JQXxw1PjrPlGgt0KLAXmQr1mnT/0q8jy3yj2qSNPP
xsw55L7qayv/s2HRkrEqvb0r3Gbga8IRIZY/Ja/BE7/7ImnUnaLQURPm7uUjyIZZ
YTZfogToVctblbql/5y3a7fCc6dS9LG2XwwC/vQUP6d7F4o3JJdYdjAlrFAmrm+m
DXw2JZZ9e2z4D9g4AuC6yoSRsj1zve/wdyWSlhnwWyNA+sIQjwfb2sRlH67PNf4w
gpaRSix8kinfTlR8hIYQoZhwK9dZkGY+pdKovaLfArTjvOxbUyO8f7thj3nKMh+o
FlMlvpTLHRLie4uwKx6lx3eVSJub6xod3ibGEraULYBnhJ+ov+iCgwFH5Q4j96+1
vfUy3+TI40XnCXBnRQ9PlNh/nMwm/jZWYSwxYT1QUP6yJvr+vRjGQGOTs3qSa3ds
SfttcGsSjyy3u677cDOcP4rNpiEBY3xc5SzF3gm21HQGRPHQ+O6s36LsqmPrqqd+
wXHXvC7+P8loPm+chXvvKXFzi2jIzHfbM8R1teHKHC7SqK/eKsiy3+PoXewJ9rWl
yte+r9lX9ZZS3hpW6vuLdIIhSExJydCeUqiunTxC30Qrpd56jb34IzCshyF+x3r0
VYujKrLhfBkJQ8KbVAgOJxPL1el0AsDNXM71Jd90qtl1r+WVB4DLog4OwL0YYTuZ
J9UMuILxDIlVDTnmYOhhLufPAySNCQdGrPFlRgAmg8AMTgP7x3nDRUlYxWYMM9lT
2IgTNupjAd4H45eC0GP6s5HaQNbKL61o10uXaUCliAeZmDE7ZH2Q12ad9vKRd2qD
l+4jJ2b/yus+7QauiI5lmEwA7TKNktQHpVWrBShJ9AHrINNrKhrrhZcNkV/GtgC4
k2JbynYRlcqMm4HNjx5/5SUULYBZiwqx9bA4E5Ud0uHqosvu/k9H3cs4R2gYt68X
Jx5diWQxdto6NsM2Irxx37Pba+O5J/lqBKAPIdo5rFsIqT01GpQY5izFayouh4RI
fgempMEv8vP1n/oR4cMn3yReOINA2KVgWWRX3PUPU3/SPwy1xlSC43HGoi2Hp6GZ
drjrC6Pgi27T8sZKQLSReEFS7+YnCeVTB9dElpoWHp1bGyIbpLqPG34iwJyQvdvk
Npmgdc9gIkI99PCSyVNkHxpRggH1hm+UemBfYMh+Ddbw7VP/oBKov5IyInihsyUe
KIodU+Fz4ymR2ZZtsFWvmnteklTBympfUilAfl42OC6Qy+6yhWarl13nPawmQJU/
chavtGcgJEU3DEApka2GD5FKRk8vyDLsRRSWbvLN8tNPhUwL9TNDwu8H9LBsFmDg
Prz0IHqpr5foJaO3xhz2okQJGIuKUAyzLXnp/u82dFnVPJvjXq7/04i9HSW9Ss7/
JLkUr9FPl2VRnXwDESJ4Ts6u+stopcVWViFG+WLaNZRlrJN/sH9qeUmOv7K3YWBc
e3qXgN8DkI5V4PTHKFJWb/MdA/N88PfWI/7fl0DDfVg5hBh7u4oArlI2BmvHIT7m
wtWeh7F0ZCr7YJ2WNYRqTuje/vEIdWS98IVDNqQ4X/BCI/QKVYzhOlteRt1EI2Sp
IX296IfFLJQF4rxmpydgUCu9VoB7Fwrac+2RAPxHkUjmR51YZdYOTZokGPjRoFQV
f7xmq2V3IhCyUt0VmLM55THbp+pDCQldGnKMnz9MQKBw4blzBFwV9guHM+aIlYO2
auuDcCh7ThrQhI/LKRdDBGzEJwOGtRIN7YHkP36d2uGSsU/RAPI6dKwaqJZMhOaL
54/+2brXpR5F4SgXZytV5+dEpFaM3CQGNLISwZXqezkR36FffQmO3c4VvCZkq5qK
uTt69cC9tRHextnHwNlYticszSvfFv5uFxvYRfictEIGnMrbj3QzHn4Hf2ga6TlC
DL/HlOEnofMO9q/UYzCHqfLGbXDx5z0sDsyLUJVQHWR6gjolnBBtXjt1L2GKgnlh
89n7WQ/DMTlCWe/5/9nP38OhgZQtbAzOeu6KwkD98VHBeDE58ZpEHXpbWuPrxYRa
qQQdvq8R+7A8afB2GdXXd/DHAGEUnMCMBykJzr5dU5dVdGstXLAzBfaOyzqOUTaw
mreUT0zEqSjRDFGpT0yQpQN4ZuKXa3f0FMY8tUoTENopQ/i7EbnAsnwwizQklezH
SkQyxC2vas+GX6+2b69Yyoq7Yr0J1C06O5SZc1RQmnNviyAapqZGXlT0TYQVeLO3
rEfBmh8K572ap8gPVexSjCcIbntrKdjTFyGVHWlx6pwSymH6ILvHoVyghX7za6fc
oKtvwZa01UgDbH1Zp9J4C7Dq8FtAPVlsOqNJ/PbcsjagWCL+iDyyTM8p4n0tKvoI
gHUvUXidu8wto66U46rEa0wnR8NSscU5u279K3SnV+OM84Cdom4UrJBtMEP0oHxP
xEqrBRhd4cUznF8UXNw+iXTEWvOnpmSuS1qjCH6lombTp2IvGciuMCNl+zfvEug1
sjBIEG/BsqpliDOUowTal4jmZNt03/Ykx6in6ub696BLfLNwkUiSLD5SoGHpW9F8
uKEMHtyKfHn+8M0G5zVrOHTnUeV4FGqRgiImAG/3BjH9R4jwMAYvwsCaG/YAag6i
nuLNiX/hDtNT+FLukV4GX3WqinRuPosnXtjst8sAwiocW5MqQw99S4J2p/xsI4xk
EZmldolo4XK9P4qtIN7FJekR8PAWX3KWmc+VtbTbU3JrVA9HLOiwXlff4h+8uSJJ
hfcazwAwQFvZVf3AuVbXcJHkjUz4H/l8qIwRXj5jYix8osHET+t2i8DNl0Il3Rqi
q6QsVaC0dB/Zs6w/rAI1yJwc+dkGv/L5kZUXndU6MvCDJNHbYNQKaB8BHLK0G94y
6T8G8CjDr4/0UH7RQxKHxxjq6hc479y9W9TvV1+ZwbrKfXduNn8pC4HAOdECrfy2
R/wOXI2n4dS+CKaAY7L10IB+niW8o0cAJbC6MCfozG9mqBbO5pUxg3PonOtvp6cS
tLP5rXTWOZ4w4OsfUhwu2TnuqhJvLC5cgOISLL+G58+MTOvP+nqiM+4TxoRhrF/o
cxsQPbCReA3ZhTrSGLbxSIwBkFcgY3P8w/L1jOS4hd0ZiUaRbQWcJZRiKeMEHWG5
hcYPLgtEFwRW9Mi38XF5JL6/aTv2dby2KY0gGMtyF/fAthMMz7ozgC5aksDDY9YA
q2yLmAFAY4Yai8w5wOqaWcyNi8SXESYq/2vXuMEwpydU5Zw2vyrR07hm4LGxrHGU
qZUud1ehsGg1byqd9cYa4e4xhZodFyCeG3AmnjsVDufh6kVfsXscForh6jgTVrSY
yZYqbuf8Lxj5R2UALI3pe1H/seTeccQpjm7ymvGpwi39lB7bkFOrIsMm4ocZXKDo
acrBZmBODicrw6S/I7doDLX9QOXqy/hvKjv3orfSAJQ6tZCdSLU32QJU6zll+snk
QTdnOTEKDksX+k+Ai0Ptlk9z9CGUbB2u7GP4FR/PjxHYEuAZmAEtp8IzAnfhfQOB
HRhnlqqMl9YQi4KPkxiIv4m75aEzvVm50Mlquifhfma+2mlkNojgf/n45loOO+iL
s8P4eVgNx5DHzY8Hop4iiLegAqRFvuE02HJN2AnKFEcgmxTKCJ8TgKoLKIxAdRPG
Zq5ugyr1Hes3sl4/ZY3XLYmYa5XmfvOLutKXQ5YbJEM+0bm337bgSkOyozThC831
QCtRLK6g3iEtMT56bwoBUsha/kUou3dKeHVnBwZfSmJG2JyDTMsKPuJXzRM1HM4m
5dUbtZrBXMueH0jMmDJeQscazxePNmvqoyA1UgaEDnlysJvL3Z6MI41tn8qKb4Co
RhEwTuvf/VgiXIiXvlRCDEYoh1iSOjVF66qtfrvRgsxeVTPbvIppSQ69PKoQzRMy
JPI89YbKOzk/jO77oRBlTvjl0okU/r7gIRzI07SgbyKjYvlEg5ozxTr62kE1uduu
4X8ihepcsx/9VdvPbIlwFZLVnwHOORE7HXem93b6m2T301zVNqQ6oE5z+UixHX+Q
zrLn3uSYULZPsvDDU2OVlQ2xyx5FARuWS2mNFG1pjQRfDDeML/GFC+kcfPtAt0b1
nryaz6A5DbITeShnyVPjUo4nnb6lY18/EiFhYO/nwwwOdEhofwD4vOjcE1kmaKCn
ZqksnY+BSew3c2u/L+KFPxYucWIeZWReVvctkj+GdHOtKY8jsrAxyUUKzI7atYZf
V9sltkZ1pofyBIiwOiIGyzj+xI8DLIAG+ug0Mw3Dq0SpYDy1tGqF2hhazEL0v/s+
i2jC3V6kw9aNW/yP914RFaGsInux+OsI26UDZHNFl8cE21YTEsTBMhDDbMVJfJkm
JowVwcDzoyHgE0bUXqgiElxU1E+UKoa83DwrkOCbkqGq5MFY/mObpgKLZNPpuDOZ
z8S5prwArJbLhf1i9pLHWOjD0G8tqntqEqqdVfbgjUrkIfzlpFhHbw6goGmRaG/Z
a/dHQmM/F6+rUCtyVNgH7ofrP3+4M9hK6L360AsSF8PjfGEG0MSHZr/oqxT+wLd+
Emz7ezB4o7non5EaN5ZuhbgMqcfHDGr/VPE340s+Jq/S7BekrgkSO2uzY3U8dsUW
HHqwqEB3005NIOcMRCpNIfpk4IxgUnOGUiKXyax2AFRgJduGVQSGVwGZLDt2LzfN
gsGryHZu/6KQXV4RbLqj9dD9LsftP5VfuVPBRTRPBCAwaCRNOYGI7eRCpV9qio+X
CaVw+Mrhpq3VsWU7zf4RInKxAPG+kasAvJrUprqMwpgkvuv4Qm7c0+e9UOn7oY48
yBsw0WnAA4Xl1OhPj1cOlPzokYmHpmz8plPTuvhZMdXBvacQJViHHSATLQFIDMA+
zKJqua/TVAZdXtf3V4k4JcaNEj5ksLNvKrVrK2TNEpGlgYMNYfmbSaoTWaCEgcQG
3LXDQ+4/wa3LOcDjXiwQhW8yVEmcDDHl4Mb3HAEZ/BzySwisgh1vm9OanLKRkqOp
0wrJJjjsbnkvuI8Vs9q+mKWlfqVtaz2l0WTJF6gh+KsX/YlfUrNJPM2qumQId+se
Samai897ifbxrz9+T2rz1dam8KEFEegpxs/7y5tg8W6f4f9XgeFxkyWXUGG+1LHZ
l/tXbm5m618zEGHY/GsfbFpZ7hs3k/PJRJ3Df3fa6blYLG22Jw8JYFQe1rdnoWUs
tcfmDonIsfzlPnvW10nFWrGilLIbgQiVTVAYIcgR99pfB2Hh4VH2RMIcK9OgqTv0
k2QeUiivIb7SjajrT+14uY9Ac6tkPz5GbgEQn0YOKSB5j6AZIL9NjoTUrT9B9Agc
Ts13SdAW11tzP5/e7T3LmfzYXxZ1hrTQFJnMmGB5mv/+1NEK4J/H9nUEn/ko2ag6
kffRxZ40hmh/A99RVdH8VLg03HzA1d6TNYfuLKd03AE8pz2aCKd35qgKa+/RJUFX
dN3e0C7JbYCdXNjUud+lma/zG3iJDRzVFHyI8hhdsuNlC0D72I2q+UNL3WFPXgdL
Zn/G7W7dD2jCUyMmoiElmpyZJyy/hctXcEI+O5i7y98p0LeY00OH0vCsq6e5scfu
0pMiX10yZpKG4nP0GEaYytvu+0KDwOiCQkbrHQ+C3j1F9Lp6i/TVDa0Dc4uKuFF7
SBzTz1Y6WCp4gleDQRMFRrb5x/45XWdUnlCGtMJyPaua+ahv6f8H3ZFMk8CUMgna
44mr4qK0kINgKyOUCt+Kau+iXxnaVlepv+hVmHvaJ3VAljnIvseddwBm0iGqOcR+
7c4YAXjteUsSVRK27XtTlqiOtjc0rMv+NaUMJnmGxdUrGAv/dfSdY9Jl5a/Mon/u
gHJMCju0PZwFRSFXTuk/XuTiINiTYiCpg6caIaGuLH0hHhcUwkAisXkbyZGUm2P7
ZruGxvlPuQPbOSaHh2JNh0T+DcqwTgMfllJWvDfVkRY1qvNN+Gz+/ak/f7lGwpuZ
aOoVp18+Qand0q1IQ7F11fGMr4vlnj5qk3NP3ZuqOIt1PUBHYVhvdWDDKKKtl73A
byf4Hqi1aBCEECQEfnkGub6S9kRtI6XDiAkLIESC0RtHWrm5YTaBn6N667ToPoSI
0kBiboT5NQGMRqGSgT0ifPhxuzXhLW1cNQ5oYKZxeHlYbfL4+UmQacF8O3JvR5X0
mgOGsQck7HBQucnlBeh6wz7gwPIFqeWhkMyViOLAaXmnlmrS23xxK+JgxYo+/ndl
ItkWO/tS/KcUIo5uDuB94PzLnSzk/2MZLbT+secm8zxY/P19JgwuYhsgsvr/4B4O
uuOA/Wb6PMh0YuEucgk9aVVne0nvEW5UubNgUZQrRjbltkxwWum/yKVcXH/qs6sR
52BRc9yWRqc1bRgB5D7vjw5lRkm7oc9TajmwaC8IE7O+2tjUoauzRNrOyCNsJt3Q
7/45yZfhFY9R/HUneHtjVTeqO4XgfMRQ/5E5+2QaXgEe9Nj3H8zcKVEwMYqePZSG
KMYFIcNy89QpE820j08G7qSBxkdMOsrpo+7Crn1M0UxzGC4xhBpFqXym4txHHPin
+OANATv+mosvrcvMskJkHJyBuztJEfeWJBdXsJR4Qi/Me+KnuMx4afeRKDUTksGI
C6n8tpXCeVh6Eh4U0oplRNhj4uBlhfYcScka8cC3B1hneUW/Yf/dKDbj6SZcl1Mt
L/V0YBUgOW00YVwPssDyEoM9YrriBhXJd3Ju9xSiBNv2Zfiec2H+oxDgTMq5UNX0
EEhW0SvNWNzjn+lKwdwAz1Owf2i5nO49yIGF+G20x3OYvz/v3FGmdSLQruhn7t48
gACfqWtkUSdEegouo03/p9ry9PGfEV9fSICockmuZwvHXLjeLO8GQ8zfV387jozU
OxdrrdjIKQQs7Uj++Zc5oNBR9G5fqSTOKcM7Q+K+ml6I3Gr1JZrUk6YF3U5OJ9zy
L12R67r8ZBhtQ5rWTiEKw0jdrNPVNBFKFUVcIsxsw0WJBM/cVEFDrs4dnWlN1Unm
+hn9ETW6/TtLblf6X5Qn6mD8UlZTqmjApIJCz8KtH7457kHi5BF41uHoM1faIQMA
xJcQ+KmluVPUXHAjcRVgEgg3bdPEf36fMmtPYBqusuyw+Nafj0rDubIIbnB+wPG1
PUp33Qjukwrkc4UY7WOKe8vtXdd2GGGCPyd3zqXNi1LbGz25viReaNKiDUOuvgRb
UxHKMnAy95vbkAaAEk00umCDOQx+06lz20fi8g60JbhyvsvGI3bZ2htcZgxNMXRF
BcablEP8KXE5f+LUi4BTjuU/RvTb+MqLLDwNCc2/UnYkpujXqNgyAWLxj2ew0K3y
TWUiOdZ3VtTOImpnATAm4gvKmw9+Orkkw1elo9txXPOgIgemWkVvEdG2I1ZysUue
3VY0mCil3N2fOA3cPsKNkP7EixAH88dbJ7KMzNCjCBFZWOBywMM15+l0UWbT7vvR
47v4MwobWPornyq1iZxUq+op1ClxUsys8vK95pHZKP89Kb6uVWkFZVkD72qAp90U
SLZxwSfdptuUYf+YNFJXK3inhCciFxASSf5cIIGFmJRJEpfutl/4n0hrBvay0b/2
8qcTqEui1KAkaPdsaUj8z0nWGQ/Ewhfv1QTh1V6ew2T6yRRlCQelmfer2QZZQvNY
tY3nGFPHYkYpJx0qV2OISEQvqDRho74Oyd1jMnGJDNI6HSyrshYfs10Skq6o/tGU
7nhj65eAYD4347y40su35UaZ7CQt3z41whSUAWaJ+tsBZ7wklTSRan6zP4UYcK6b
pFCZW2WAcl7zTW1BQDm+oefPigut8S0ce9eojkk8gokLLDg9iwCr/G4p9WPunwAm
jWXN3WyWeh30gm0hmUGljMJGXqrYzJsRtr3zYWBrxYJ+iD8OYX8Hk20P+RYtJU9N
jJpeeKTAwJ6bMEiML7VSupz/1rnT6LQGOgeL9BOaKBctoc1NRayBMwDbvSpDJOgq
NlWHzkEYKXFjgN6KOshCw68aFMsKVT/97MsAoy9XdUO58dlxVnnFUOVcxgCwlebQ
hhcBl/hc/W56782+rlM2HA9O7ffMS3STMV+7PgN6l6RIV1WArJWs3LkQiSJG2qnq
u6uYv5fNzauflGajxX/tBKZH86USnJiBBKMgAkT5Eel7RLSSLdx3Xh4XxqtrEMp/
gC6G8/LlTkbGtStwX1SCIur2hxawQULabLRlIMc+sQMJUtTxm2F7bCZtwKFQEL4j
HAJ61WufmLcFdWaWIdMMyJ+XlSia3AYEydfpBz8iJZQW1px/ppq1gKM4NVhGd0vg
zpcGVh+yYRafWfw2z4Uvm8W49Dl+JgTvRbvPQjsj+uQ0bxLNlwmDIHSkmct/jhVH
dCupQT6gYg45kVWwahQhNe+AnS4P4ZY4sInbEi4i+CpiNo2N1mZ/478YZK9aATme
CmQ7UacBIFOFvOze6PgAq9K8CkwLpBM4MVjcIqcAA0jKMHIWcbNYYajoUrjsoUEe
ZJW11TdC25dwFaQLWlyW3qVbllRuJHKy0PCI2lZ4WDHmbsCNmz73YzWUtSiqdNfr
whRCQgS2cNpJ2DP9ej3LnRaSwDTWH+sR6g/7FiGyooyhzNPvDoe3eBZisVgplzEb
0DR4sqAZn64RGpxkC50IE8Ge910++HkAjayCccfdOA31VhKEcMm1i2G8PpbWAfqN
pMgf51iuryZSuD/MhLhIYF1Ar0X10+sQPrYCa/j4cANBgMtSe3OHiM7A9gr/T608
BphDfLtSmJWk6+N3TTIWBaGOFA61i5wEHvlhN6idhObc02m+Y4iRFRntRiWFXgey
x44fFtgrgdcXaXOotVGzrZk249jyOy3J50MpeuHpDSFeOKtXm1PL4in9HEjk1CBz
67vdJgCnKkv2fQNI54lK2UnhQjZHBZg0Jd406++QtxNncUhWepnEqZhMBe29ni1r
IN/jgX/N9/38idm2BsvhTND60m9K2ZrdCotmneAYQfD0BMko2zMwIjO4YXlTJhOd
02A6573PVBMuc1mBHBoDfOItZTvWcD1HdUI8quPICZ5xK6PUWJkan4lV1BqSjymp
V0W3FUQHoVLcoTrU9quHE1nFNEr/gn/kLIxSflWmIiqZAxnHZWbPJLVwV1k8tAtr
JRIOpOJU1ZSOr4pUkupoERZD5yTtpDHW256qDaoQdP60N8cuXmK/qRJYwGVTCHZ6
jCSlrUaumetxuPga26WXFM6JttsxZrjkF7HiXmlVWpDy0vRHa2rLt138dEIqIx9C
cPMjvECXRC8DBPy0GODrw+ZLZonVlCQQPkC8wTadK7reHref/wIX906b66/ZDz06
V1QJ/Xl5e4dJf5esktFaMJEKmjX1EUEL3A5Yy8xBwt7Kyae8m1hcV/qogEuIG4jm
dbySZkD2gTZI65eOZN8K90XySO42qLGcMaUfP7MQEA1yYWUmDHXa67NrkcLS2Dyj
xDDpuPmub6u8myUaY9cR69P/i2ETskV92HXUFxzX21E2DOz8fkqFr6nJrkeJ8oJ+
nRxa2OfWa0WlOJ50oHn/OvD0ia9kBuv3u0VUEjZOw5xyKMiSh1Ivdrw991UysKvU
riD9ZYgaH3+9sbOz4d8zd3M/RRCdiYXrQNpfMg2McaWE8bT0SHzJzIfd9DNF6wik
L6rWi+XduxUTP1ZjlvL64zOUv8JVpRTqrvQ0dl4N+4Z27wUvESW2jRxBkOy2AT9m
MAfuqNutvxGkGFQq9Rbfm+mmV7PwtrbE77FI9MU+VuoEbTzoiPdudgVYexecrnrB
xWgVIbogGp2gunBY6goRgXiJ5LSV9a1QOpg2DVdZ5/j5+BO86/b8kCsedhmC8TgB
zabbcbrIZMewRb1Lv3edD9L9qRAGxRWM3k0KQYJpTG6ehePgjUpjb8qmYg4C5l+q
eGPpxAgbyzYod9SCMkmopN6oFih2PNpcKwoXC+AArKZpr67SAKYLvzaO0RzNliW3
hq9FDwir9nRJT2QTHQEm/lMJ/aCJesJN7SoRle5FLwy25odBcdDphqyhdoXH72zX
hOm4G/ntUldegoxfk4Q0dnQN0yaH67odNFb+FVTcF7dJezzCLYTNT+KrtUwyS+/Q
RN1PDOlH4c2fiOnN1g9AnFbMMWWfF9Od9iNQcAHhCnEE2tZLguJDuWxq3p6pouwg
B8V13+pZUibgrw2cSOAr2AHQC+6x3m8j1Kc2PRTO+4JmdzgjJ2E5z6OWZoH69SxC
5VJ+S2R3EuMZ5vZjp/QXxDRIS8wTlM4Uyb3MiEVc9Ju804WGDmC8j8wcICyjLqnp
k3bmvmr9oilcG2N6vTMBbjMYgzCI4w803SCKIDpswL/qe7p4EePKZ7Bdqd4+9WwR
haICgHnilJNB8aSLnV3Ekj3eKHVGaP9jeuYl4AqJzE3tkLiDngqN64nRxALM0byM
ub8p/K701fkYR9fTHYnbPqG7c05TbB9q+5GpijOQqt4SGCtAQ7+UM0eWFpS+SwCO
rs+EXEXoidG73CUKlZq/z+d7AzxwftLl47++UQQdWerNs4EYG8AEwv01AHBL0e8o
PKha7+eBaXnpxzipC4MPMhm7QcvBAaUFVwPVEtJGymG//4ec1UF43pI1/VpsgJJf
gRU/wALhwaoEzH+w8/FpgHvQ8Oxf67VvNMSHVYEjSkv1R/ftaUTQq7OkDLpyg7Rn
//cwMN+1W6Z48vvAyS+s2ZKJI0LDl6gsEGVEv+E6jKH86tGGQJ7ZHEnr9KSYWnJj
nu3nBmP9MvuROwnkMPAjsJJ1KobWmHp69YAIzhojjHBdhscs/mZEAL3iToTkyV+H
JOk0GgABWzKNxNgGc/wOl0/qLntYg8CPKbJ59ebqiKOOyg166u1p1iuEkc5QgVDZ
g+LeDqUfvC0/trqAvdnmv0DRLBqxjXrpXauQ4SEVPjS+oUdYrhSG+eEAIIw8kVW2
4eF2i0wTksd4c3CIfovMydi0RGk6/mzfY6eR2ee+kecns4TRCNnhWlV6bcSs/At4
18wR1Jmb3VCS4ct0MBXkIQ/5vlF4H00mPX/J5xMWcoVmGfGVjpIkqZzVguskaXkC
MDV7dlBY844HEF+abHQeWEjexFv93HD7eeSzHwRRwaYI6+Fj4P+TOQAZ/GaFGkY2
bVjEpKdHsVkQg6jI2OOwMgOYtM2CQA3CtLD0UZh89cgFM0tfY7W7cKuhrkFarouB
mrHzYl+EqTV1hpp4nOvEvsEGM55Y6+cl2bNM3v3gcGvflWOvQYAZcc7wRzpLyq8S
kJ/Zpksj4wtxuYtgYw2OTQ9pJJSGrbfgMLUmEbh+yuFnsbHudArqDelHaoaJonyR
zhJiWc22YkpS8v28ceVpH/KCbbMmAeo3qREFEpMpMNsH72kgM/jKEVRH6agdzXAt
I5rMnkY+hbfZ1Wbd371CHyylP4e0I4CEPVdwp6uVQoGtQ1ph+Y/JxIN3fZrSynnE
yJhDG3Cup+UbRCChTmIaU0A+n1mgRzaATs8jGA9Ory4GD3eHYle13CAK3Ophe/A2
A3RE9l4APH1sn0ncxpjIxtE4Rc+QYcSXgkblr7dDYmR3Ewvjioc0vkXp3fa6iAMF
E7fC73zvwqey3BpW9FhJ/n1c0z5fousr9L7F7dfSch8Uia6G2vo0/xUa90cT1/L3
oX+rslUFgVSxONzNysSL7P8V7SomyRTr0gkzx4uZ1FV0JbfKgpreVewn4enVGEw/
jpEoamZCJdqQm3CZJPifIy0J44O7kHFfuS41jQVkWRM4cifh6+kaA8wwGZL6yWhk
g2RPq+w/4aAbRtyYQjX2EUGVuoLVdfa5LJp3J2LAiDnL33GWgUmNv3l8IKHq10Nz
eiA4P73A/ty41oPhquL/uSHCywhd4j/y1h0+IWy0CP38pMDfyIOGrFmIcI2OPtoP
P3hmYZLFbp0xiQQzY/nuWtWpfHhGs4cRO/uVMawoyf55ljuZe0EWYrk++PVOlYak
Wsg8MkhtAIeu2Xl9ld2bSom3XoZ6wVW7h+V9IZ8WQgtR1RjOpjO2yvxDiaKm95Pe
SXVDJi8QS4J+klfF8RhzErum244MUk/7v8ZdJrbKnN7cO9ZIXQi/9aeyMbO1iA/b
UBWaXG9s8VZOffM/nZmw2g3ICm/OndbNH8XMtq91gwZQKJB/D/dOM4XA8bpC2n7d
w5SB7tV7pa92AO7SohJavFMTEPcgO9hYxYvDEPK5CqAtFAYNPNmkDZTu4GLJkYXa
ONQecMoHWZbn1GyOMcm/SBihTDRW2omjER0DuPbzbVY934V9D8uUCfLuWidJlrx9
wKP2TEG1gJiV7lGOW9R3KD4DbAhR6Mp8QYKhDEW2PW7RSNk4h0msxWS6p9dYOhw9
yV/YKsDtPP6gJYxcNGXW+6SdOFmfORqg/QFHIHze/amHzFAPunM+rXmnH9RvhXxb
tBgGW+ogN3ahvQsbewLIi7CVGIZOLA1ApxEI/6GX9AJ13sIo+T8rWlTBzA8Yawbi
+CUyS2FzJr81gIdyKwXOH1apeQyDl1qzhdAG2kPu6FfArcfEdnyKY98YaHwJH/Xj
sYPSu60KYV9izi80/t9Up2xHqK23DHmavLjVjLBfjG91lvS/hbEU7RmNMn2Ue6jJ
lbeCN98SsgP6hLpupkCCUEHXElsVwv3Fw8ChrK77Osg3gcGkv/Bur7jd79dFBpQr
V7Dl7sDRbr2/spJ+g+ZzYS15mQdXnhRnksNi8AOxJa/uwe95w8WxYSajsT2aDhQ5
2yG615aQebG8FnTd/BDS52dskpk6Z8JIOvQl/whDM7URxNLgCX8fp8tbLYJMvQ5C
1fjRThRyOXJ3zcANuqyW/q/vLubRQyUXuwphcMMLVIZ3LSLmwXv29kYLFReS52f+
BU7DEUyl9GN6ctkQrVcAfdHUeg3YTJGYHGtUNY2LCwTnlWF0T9FswpnEVV9GKXx0
GUWW91m2I809/sUHrEbHXplmEha3SjcZaarMHEJlvY6Lt3hAOGVI9s1pYvuCa2sV
Ubj25oO/kZZXhhE60ed+h4DGhaSsFBfhxn7n+noN0EI+uxq88Jrvn7mb7DhfMtT4
SlS4aSX6FCRxEYrO+80kcg3uVVzU9Gx//cZF/GYd48LwGHqJ/+XXrxJ8JEHXZsRM
YmjjRAGOkjM+NR400IHmiaYDNNt0kaexI3sPOCMoM7o16PKAxoUEtgaipM3/0vKH
DQY6885YR2BpMJpepKg3w4mny5A0RRBXzFVYPB7jIg5PKBQBVVJpjjnzpQUxtEXi
s/Xz0U9Md5g5FBSdpiuXm/M8XuCpA2i4xu3FGTXOxpCKXhsi09GzIb196qrtmc5d
fcZXmjYP/ZiD8N7yd4/4Ren32QvfvkukY5XQXgwhLC87AN/5vViiNezXpeojhIBx
La7KCQi792Y6va1yyay6QhGYSupWSf31OIc/YmUYKgi4RXsF0rAmKRszhVAx1Uoq
ihDLlh+vi6twIh+TO/1Q79F+zB/OxX5ob7PbP4TeO/LnWdbx4TyLeMm2RYnx9XPM
Z46yQ2HozOyu7jp6H2P0lPW0evMb6g17x2StQOhLOzO56XiqArC703/WjoiDD52x
KB6QuSmouAB+fzP5GlrdddZhMLjtfNlDPuIAhsb6q+mjkKq6PDYfuLfYIr1npZ0h
zRRGLK7WnIisdnN/gtZBTn0dgo9Sm1TbURRCNlvSWlqiyxh0aGWh6yWWHim0yrvq
vFYDq8q3euJDraA3wsQgNnkik1Rp+q0wAg5+66JwM5xfDRHcjGKILcvNWMO2PBv9
4+hzujGstCcLRhkadv0Ief3/3DkZ6ijrBNtMYRKuTPDI9XGIMOelyryoh1vLK2DL
4SLKKHCWasn+3GbrAWgHp6p+EaCgFk7ujDstDl0RFUaUWHaEdwCN5DAKotw0sMQg
CBgjk2j4iCFByfE4Qtd58wDZeCOCziBX5h1qnKUFf7703hOvSFJV1F5oLoLJLeHk
Tzm4qfNht9HYs84f0iHC+4mSnKv3g8raLURdi0ucyI+nFFM7l6SULWNYf53Bs1Ow
hWLkmxi6pHFLm4SsWkkPw0PLHlzSqTZuN7QeeS28m3cWZ1leOjXtjqwz37gRh9+U
jLAjoF+eks+PWI2XS93iRXhykS8J/VF0b50BQXJRBV87hFsjw6hW1W7KX+qj0uAK
SVgjzDC5+Qpk29rkPnBswrULYh210TsYCADD+7Bqe8Bu0dmBH6DMNtRtI+w2322j
k6AuXGwumdziCouHgTgCRyHr9DdoWvTK2BJQ6MVCYbmmTzkvCAirozZdwBINFPr/
zdRuB8F7ho0o4PYlASlGSdN2bkR6Wu6yirfRXvvN1fnU7p2YfayWd6wBpHEI1aPz
K2tdsSxP1sW/u5UMm64BpdHG0DXhX8fPs1DGpPYK0wjciuXvTdhifym0iOyjho9+
+NUwRYDSON438akrNs2UHBgSn/k31ovo3Dg4bTOmoDjtFhusr8GKpTDGL/kLjFGt
c1Ozd92v+5RM5QwwRaoSLcrmQL5GkUfnQeos+cIRWUiBi8n1Dkz3wBMVOgF4QcYX
VS7jM7dn0gHQJZgMt9hfOiB7ZN8YtQ4F49owkso2AHG7Lk7wvw7VOgN9ytIoavbV
TdF7hPORALaJ/BrPbUepydj+bt9fiscexeC/muXdJbfm2Spo9cAdpvsrjNyF2j8a
lxcvVbsv7KC+6seHpWNT6XEdihANBkfIrehSer/y0wBEPAP1V+QxvS9etB/IEM2L
ZNodlM7sjUpcjUiC95a+JryCawOn3FTHLZmaPBW9kzKcA1whJzCU4em294R5V5Ye
/u2qy4AlKvIkh1hfYuEWPoNQz3dWdinHJhqxAZ+3vC4tazXMY4CStGHu4YRtmCu9
nXEv0Xb9NT8caqSKgw8qRiR4z/OYICZAWCXbMJy5H/M2uIrbIioaqrgTdcIycnMr
v1y4vDBHm7S+ZP/WQY3qo5lTEuu3iF2HVLLOQubNRxCWilkmakXsU8KE86y72bU0
03HYsm/BBawIlMHfzmqohpHd6Ymg5V1S+BWvG8QjWJKMZhNEA60y0pQ1/Wyxa7fT
T8QRBbjn416WwHzdBW3n8aFijWtbyspOrg+1luMNkw8gQXTQ0ePLEB04PNUG7ega
eIdOmydg81FKEx+UUol8R48qMEKTo63Rl7olpRrg6MmQe5hzxIBBoJsNCXSmh8tO
FMdlAQ1ByOKvIbo42Vio62M6NFWjvzp4oJtSW5Mc4HD+w0jzCTcB4tGpCJ6DsDJq
zTDMsXdPvKUCMGMCT9t+KYyf0YVo3yeE+d7C37ZsGXV/ZOrZrqJuaPEYz4gNtKHh
BSpw2i/ua7BGDRvn3fTDqGZSZcr1KhQPxDdj/IlAC8cHgkaUrV24v28el4uEkwSM
J7L79dPDUgVCqic/yaE0Px90w6Yf7Svwlhdyqi2WzTgiZ6oq49bw9epxh6mr0JSB
0oYGQFW3AfnhCBH45RcyY03OlqAURywO+Phkx/ZQR1Jg+7y9oDbqZJdn3r/iEjy+
FeLNGMeY+e8YGolgFzMIZJZT05WvNVrd0WQrFgAnCYLo5OA/1FbDMBmCukRITxQQ
mE7GklM2V2QPNhT2hNYqdKjwpdubyB4KfX6F+KpK99bfLfpHFRb42hVIOXHBy+Ou
EOVmqhZGfmCAiDOichscRQp5NnbLo5kKt/u+heP/yt0hNS4T2uzBo8tHJ1XH+fFD
oskItagOeDO57bzKvZOMRmkduNNwZw7U+qVUFoUKmqoK62nn+kcuonXfZAZ+mULR
5X2iS8Erld6AU7f6Ydrlsefwa/xTUyJle+wJYdWOWd5U4KzTXqRW7EkIE72SS1qU
DOJLOZfpiitB9D4iTwHvtV0S+fDOze/orIOpoLBx9tkk3LW6x5x/zAbpfhsrYpMQ
bJsUBfOxmPS1hbc+bqFfwdAZ9vjO1R1Enx++ChnE4V5rCVFr9UIYMubRZvwNxNEp
dRwjoRIHtH2cjefoMQH+LO1OIuMTUv7eij8Ao8eehQgx6lDPeA3NIZoAt029sDzG
+dlfpAiiGbDQPl5Xr8qsZPskwKbuPrCA91+S1BRrbbuUq6F/sLfNAUw7DXYgKIyz
WGMcmxrP6MJifstM1yvbqfZ60V5fQDlUW/bWidMmSbWQ2EB1UC7IU/4kmLs/rdV9
j7XjvoDMRs/jP5E4p2CDWo14MQIW/mxXzEnApwo3z2ImuZJCF3dFgIm7qUpC8QMs
HRB/ZH+G+9LY+K//VOnmoltai+ooKiNNUP7+CIxi67VlH+GiKsUCHriREYHLXsGA
r/VGOdaAymwDrKPRsjYYkJGBbnLjj5lH7muM4Zv27jf/nt6IJflxBmVkf1gT5Dk2
Fmgb9AGBvVA8c9c6lipHrdDGOXbIbHzu+sqOYr5RVjTzcmBWxS6PTHAkjt4maZIB
veurmKIRLAllBi8HUzc/fxMjnCwv/irOtyykuGGnwrTliZbIMu4kdfMemhdg309Q
ZuPc0HvFKKF/ZiuTFM9I0FuyVRQM1t0lCXTicXgaWMPsNY5XVb5IMmWrb7aQqAUG
0n015Vj2RJOllF3J+dtusK17d3WiPsn64YwXaX2V5dI/VwH52lshPl8Mz6WWpv4I
bXPPCvKcxUhZDvNgeKpnraXetXcpTkk2EIX2a7bS+7YyTcOmV8qTR0iH1Lgz4Yma
gRx4GTnSmBCgmGpZ/iiBfJxApcFOk0mfnmfH3LNCws5ZpUnAYnsDhrpv0xppHRCn
Zjha9Uj2pw8lOi0Ev5kEOxRScPwVYR3lqKoLdibDN0ha+2KkoC0k2/Bh0YJw5TpZ
Gv56vRZR82GFcl0hSmkqDxx7ZTmrJb0HRihWpnwk98PHXG0CCEYraUm3Ke2m22Ca
2DnfySdYoUtYM+D8UpekzRkeFWKb1l5NBUpkBn/jwDKPwDizIE05RmRjyOhIQH41
RRBx22o98ItMtUH+vkQHHvbBt8LCRoSfV/FatWrm/3TeJwlqcRBMMJLyGb0Iq4oR
BlJE1SSm+BmdzBkgWNxhJ7EIsclFMBgEPiUburyUBPO2mN6r7MHLPe5rHax+uL4O
HxSuJeY8ygeI2oi26hOoVWV0yUrB+8hTwgcucTWZ8YOqgXlkxrSYR2GPF8Y/jgxb
XHIZzImRacmBHmBQPG65lnXgOzvrrI+woQx2PJg5tkcvXGNKUOcPnVLZogWbuMtB
E/8N2nSqR3mJLULA+pEawwzREj/EaLtSXbh3yOpLs7ukFrH+lQGrKnzCUBSJMOuF
DunWVhOcVzyXz+h725bZQ4sI4vZR0ja9JXZZJNvvNr26RAHqKsv+8azeE+wOpzkG
qZoTmgeXhuVs/14y3HNu+wL6/0ns6rdCH4KHJVRu8upuOxon9lhAtPpOOPeFCxUz
z04nJj6E/0SmfUNJe+0za08SN92kPES5sIlWe9MhssvMr6+K45xeHg2NLde/4pSI
W6t3jzX17jGbSB0hxMpo18nzqo88ovWR/3zZRxhHxnaUkwdIaBB06VA45y/jRhYY
Pmyo8iRMQuZhehHtgln2bmAFBiybWUaK0p1Yxhlp4Yv5rs7gy++YYEwL2PobtV5R
qBKygaYwqs8uip3BmOq3lkqjPpumJcBqpFiT13UqraH2PXkFvzmxO9XNOyI9qCRd
/CLiEKK6WZUj1MNY+GJx3OTkTb5VyO1DZT15ORh/BpMa5wpp7dgwYj3NOoIwyZZW
LtHLEddJDgiOLjMdOWpxePK/2mPnwH+MnDajpg78mw2rUd2Bmlz3sOGtkgs7RVc9
QMWWAmx1/azwqd6ZrMwKqxmkrbgbpRn5uW8LikdE/y7kH09hvn+ZkyfA+wov6YB6
FU1wsZototw39A00A9o1H4dbqGyJIWi7fnIoKjZmk2yDTSKOPeq/nMakVuLCWV2S
srHHTqcJ1P0WXRoCkcGF01gRwc//aEDOfVKtX3msl6bTMG43oqlO9//YUT/7NBem
4TDG+PBc7ctlooKGZ9INFfFZh1pZC9obhTMEJ1ZrzbdFwqKX58km97uRKYV0pfZr
AtUDuRPW07Sym3vVdgjD+uTPUvjRsRIH5XVpRBsRVtlIH/XMxtyMxN0LzuFb+v/K
S24qytb8HoNPhiMbpKQ0nbcCwiSj7IwhsYjVXkvoktpGR/4AQFH/jnu0ZQabgO7Q
sm3fe237CLFYrRie4AkDeav3n7C79ZfK6IVl4bi0RT1Apjoyo0SpCjGUn/bZ3bqY
wEINBCCLrQa7iK8IRqqCozsrOnCukpMwWuA6Io5Jbfu0/QHscNfKJTW6rJtU1kZA
yhJ+bHRTNWc2aEvgdF9fxj8JVhkQ2B7CVxBAJPcDDYPRkTz0tFRWknMncIU/Kg5D
q5fx7VSSBNlOBgrs6kIgC19IWFhmMJ/dBMMVQaF162CELfmrrQ949+/IxTDf9QuV
36qmLduGy2xAE+hnmYxULaJ/1W/G4DZ1i6ahtDQRtj2Zzofm6FNoZq2k0D2teYyu
1yousaSLH4tt3xNxu/G3F4noaDFwwfTm/u5iHd1h47e4nSmJfl3j81ITBNHSw3lq
pksSjpkPHwyiHyin1lzZYuO5lWwoLi5FFqd4Pw1nCmKMVoACsIVt9AYupLw/jMZT
A9YiXr0YW16serXLfW6Z1+oTFIcB4wB2hMOLD49Yxnm3wQLIC1G/aqF4/7FwLw9+
09Whh0kpDT6qylNsqtRZGacVX7MCv6T7BZcbQv0Utlyy2yix4zkaJNUxinGkq+Ef
CF0vA23HYrJyKtP/WwMZ1Tw4wybBqjIiyhMftIytPZ0CXVCYUoIQStfpokV1aUG8
X9vHxDsNCGxGTVKS27o9LTYpehCC4ofG9ZXBXD+BLkUaC+M70WkkBItyLUxE91yz
2Cx87BFe1zN8OHk8LPqQVz9oJDabblf56hSWmDodjYI+hcSlPsBRIY+WEjkwAtob
THETPgiNGe6dU4tt+meecx7Cf4FyrgdZbEO0r3VQndO/pZS9BAY05hQr81OpCQWa
fniy5QsPkF5PiShcvPEQMGpPu19kLE1VQ3NCHBZA+IdrQEBqZPQXVc3nr1ab7HZ6
XN4qB4ATb7iOb3EbW2/LB8UjMuzjhCqOiUOGJFicl3edg066YCjz2vV9skwb587E
bUvNhSPTlK9BJNriFbWZ4eF6xiJXQ8sZkjqN4jqveJ2NdBEiU3RNNLe20yKc5c8w
sJOApd1caFrhq/IQDvMY8d84/6nyGhAStX1LIbxS0q4agsVa1LZsKqIso7bCrsFs
MminN6H395ECf89MrV7vDgnbRxbyi7T2dyEBvVnHukIVVgES3HWuniFGgCCB37mV
s48NPiXYbpoh12e8+su8NaIUMnbKNrvYBjR/d/j+cbOZYkn8e4RAnN6w8TVLJACP
a4sDSnZJfIQa8jnwIRU+tJno35TgFGQ58HLQnTEQoEbGwH5VTSSl31VTS2/PfXx2
OEbrUk4VBf9/YTevmXC8A1ZVOhrfm1L7aQ5yrLwU7ciKSMWKF4vNJBLLUro/o8W+
qPxQ8uwsceN3D4abbtkgMU1BuDh35gKkkUS0zAD1SLF8cPSfFVPUcn9WquFgpyh3
qq/hMxRLoxwJKfh1Gr27SjO3fjR+mmIaId5y+sZosYI9hUV0jqmmoEUGbrOkVj6R
bd5aQzBwwPdSR4SxoQQaJK+0huhyNUOkRv/BmPBdfzbJWSvMCjpwfjf1PBLWILPL
CjL4C0PV65iK8d8r0G+GFhRWz4aX9ivf+EDPgD0372dQFdG3qxUj7/NFZpouNBBj
jv5w/a+01Dai0du3gAFmJetwG71n3g2Lp41RdJ2y/OYYciAvdLBeliiiFBS58Ilj
NJ8C9gYTHf+fgsNzneEpgOk3mOG9F/iH2GX3OfnLSa858/7mLZRE1EzVCNHWuxnw
krCibivdnReIxGwDOaw/Oue9Qd0Fhw/Ev2ddauRss7Bw0Sy5/hqPacISGoETzOe3
y6e7nZ5XmFxY9vLR03Rni/v33yFHhZSbz8aawXVfAU1gfsaMMKy7d8mAi1qxA4tJ
+zA5oICS/cowAS5UXbqtfOFodJUWnbfjutrIX+0MhvSQoayBNIEy0KGV2vtKSOqq
VSugXn8ACn8CXVHHEe+LqNqa8djrNkumUN4jqEIieFsvhRd9QuRqo5rYU5gLL9KX
cePQmeVY84bztdc2hffc+JL11GmznSK6xTugTkZEWjVJ/1wgb+llUfLIau1xJ63e
z6CPQLI3exk5LaeLyN2q8/ysaglb7vD7IHZFSfsEikBVsa6adEBLCIg32CnVXrAp
81DjiZbrOG53VzLQ3S1iiI4E2LLNrA1Q6HASz9MIWl/89X236QHd5BZUgS03j9vZ
BR4cJfMlSlAnbaOF5O1AgnL9L01hAHIegxMpBEE/Rc6cFm7jPZJiuptKKuFj2B9m
7rN7YqUkEojN+ck7mPICb/LJ+MDenyfplQq81G2zrrWTgAAfvMnh4liVp+gGJlYj
DFY0Xwe1tmidaJ0SN66m988cnyLGgaZNSG33sJ6nU+ZxS4+QcmWI34eLrSwhmq7i
KJFACTmrJXSYt+f/AxLRhikYuhXxF4IcGTjialab27qplXK/d4Vhu1RP4GRuyWUp
j0YeTHdvSf5nXAFa/wvH//t2nqFk4xDqXGhU4YPyU4yTpM3Nu+6ZzXRUymMbphDQ
m94Op/xdkwFEUSH1fiEmBIEIwH96Blu7BLIG9mIS0Z5qk5VpjV6CDfmAaKX5bZ0/
GYGQq/aNOSn7Bv/DuoENHnj5V/B8lUvxiyaPrjs/alM+GIhH4nf8Q4VZtDe8lMT9
yDEcUi4BD4DFODM3xoXPzhzpa1PNw5oOUQIibKH39feSsjI5wwyvw4ypFMJGtc3s
8yMFVmLH+fsC9g/aCYPV0QYigTTvKSfWFQpAr17WJjCZEvySa2eITq+vUwrErJ5+
D5S+Kj41jaUOlmpHfpKz9Dq6okRqXBj4lkpR6EyrYqP/OZfkNL9hyY2EG56t6Pv6
j19X7HD5tvo7VfaNb+8ECeDhoiYMQJUTTDDrtzAJXRF59Vaszj/OSzaCMmQfrtIo
+ahltHzvffLoqxJBcnQ/vxQD3w+XNwBycte4JWC47NSeGWUewwdwQudk+68F20MO
sx6dKkU45PNqigxKqe5zt6v5987D1IGAScJ454wiTcuMTtmweuMykt6AOewZAIne
/EfX1dN/Rcf7qHMaq2pJVWlHqL9f8a/EVVbVAePzWhIP9JZ0nrjAmWvUyY4kXSQS
wS2OgJ5A3yEDYhw/32QaWO9cQxMlICu55bXxyhwrcSJjhqPn0XbOdqf7/xaL9iHk
nkPBhT07slQo7T2ZoXS80/sJwytNTxspcKoVbM3Ki06USFUai/PH0ME8ME4jnoaz
ss10XsBTG2AaS0JiCpNSFqL+X9POAZHbQdLP058e6/9XnT289nAE2xNhxcXR9hB2
DRX3djPvA8cd1hMar9iUWulHVnZhmT/BWQ+7doIrElEKwpAYi1tnweYCXEtHf4Lq
PzjicrLQh30gpav1Pd2XLabHZW2cpYjKIcJHMvzO9wuUd36+5/6TkBiLYnnssLGF
0KgRfcemcBF22dZ281tiisgl+544ZYQ9mgllJsSef7lau4XN9m/8ry8B3ckaFYNy
DBEwRq2KU0sZ7DQeTPb/XiH5vh6npYSxRW4phFQfw5b1gE94V3C6Q39ShtUFqME6
nbcSHhPNk+RyoOp5+ewiMZ0UXQmiC+WFoDGzlDrYkfZl1UmLFJKAcOQDTC4jwnVj
RWjcB+7MwnXYYtHpknU3gkIrUHNXEbKybL7qDQiH5+fY9dwiaHN9Y2hJY1JyeOZo
VDwlPC4AaG/yWpu4ytlLsEPP/EBW4fS1Lemj6667MQnkDj0Yn66CEE6WjcD+oTv+
64fmqNbzY6OqGoWKha3V0xAH1sYyqE6Mcsm/klsGDv5LyZAD7voLiFeeMskvkTCE
AuH3shraEx68DAwQ1nzsMbKjZYkLdvwoMiNWkCZbo1MFK5BcdnCB1Tx1Ml6l8arn
4f+eZOzO1j/hMt3X3Zj0lyx1cBht71nC8UrCPP4aYajJ3Z/LvbGBmXjmpvCeoegr
Lx2Yo3dGypdjybGBi2/6rHeyDPjFPN4JXwFXrMtJeN6Y/cntYQOQK4+dP4zMIlAQ
KrQ7HW/j0eVrNVk2DsKTKA4pdy5Po1H6Q+kN2Ug1LYhVcVN8CUlmF2T5ZeEX4ZYQ
I9FFPsi27vQR9PXHYbAyytz0mh6KRA0JYqmLY1wSrPUxlOeLEjaAQeUTjljh5faA
In0JwkYhoHSneir6wBD0QaqGxBoOqWyWjsym70FgWYvuckeIcd0CgX3Z0BnldsZZ
uo/np/X0jdzlBF2RU9LS1bnUSjbXOeZfkflqQRRC2N9JVwrquHJcC4G9qnExrr+M
KWb572EESILOfbyqnnslq12wciSm2NBlIAO9zY4vhPFCLTqW3Dh8/jemA16bN03V
WJV6khcbWIMgoh9UgM56b/jfz7j6ZHJv41nSqfmVNsnV8eeBF5fRxSxd8J95Qwa0
9mFvTd0A+WTGpUG0LpSJru5+Bdq0rSgpsyNUz8e54SFI28zuJguEif36td3njuiL
n3UacL5+nQraIgaeYE1T6/kI5xWTMUpu+SR3ZB6AXW0ZTP8xRnkUUmNtK/WqqceH
cHQsZU+mfiCfBg3hDUno/s5UksVCe4gk5TSHRqkbv5NW03p+d5X/0ZwBBxTfnf1/
gesGEUuu3v4EkmId+/5utgVd6mpJOa6nEvIKO06jqa03j48ADGqrr010Fqm2GfDv
4bvCrW3jOr3BU+Zr3QlHWeWQwEEo/QPzlt8fbLtP1QG5zeUh5ODv5BbMqIhNTq3S
6tNVc3jfBRMaYnF4WcUT3RhVplLFCIMQt7NSQKt7Mkn3rd9WYCiPUDkporEIEErz
GqQBIWF0awArSD+Ds2MpBudgzjbgG8W6ftEK2xjfwNAmPaFm7lWz4d7FbJMvIb85
l7GuEeXNFY3WwmKlio2f2GbooMy95IJO7cW0rOijJhSbggLyjbYydC4pwWKT9UrQ
VeFGCHs7EWq8VADpSYgS457fKYcw4p2z/fxazNC8LRf2foVF9Xhzn44uIZDdj9E9
vwSGu/0H3zB0rR+gqXvrzXyQyFtfK/eh0R8mGnJnWj6R1L+x0q2hlS7KiOnE4xcf
6khGawwiRHg0ArCDn7mntbVYEzaWvnt1pX0KXSCzfJv4PdsEP7KwLufebx8oRYGJ
cGnUdfzmDu4ccc7g7V9BHuN8SU5UJnCItZOGmnDdf/2nta6bGphozdkIL1Bb0A81
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZX1ccnVWL+M8kH4XHuDNQ892GVI7Lht42kRJIO8Dwz0rKkRqsy/yadU+PnDoZxW
Rr0m/bgaNWqFxC9IrTNrqgeXhUQrmwm+Y2QjjqP6NiaW+7+GmtSaiE+mXgSuyxnz
1MvecqP6DH+Et2tYIAwUxp9yJpexzgU3GLF1Ok7NwrD4/z2ULdtfXRkEacCThnR2
FoFKdbcDDYp9fvWApAOvl52TPrY04t86I9JgCKjVt2ibCFy00XujYZ9fJxvv3Ifu
C9SujtTEwss0+l0Mqn9dRLV9mDcil63LAD0wxjDVqJ39KcLf91idLdAyLd6Oiah6
GR/sSyrgos3RCbTYaucM/ilcE1E21+klMLC2ya08AIQTW2eWJ6SelTpCugcUKuXb
hQiscW5ZIix1L9aUVyKijG7HuIUAbwT1z/zkS2ubMtFuBzv5jF5JT1k+f0QVwmOC
77WiOEMed/a+zkxPCXnBOEwQ7fzTl3KiPf02aZTNfot4tGVxukudaHFExaug/5cI
L1r98K+Z+/MY0hoYjVV75A==
`protect END_PROTECTED

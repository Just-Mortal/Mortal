`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QU5ejx33Y8rEOBnvet5pQrXDmB4gxBFCM3OE6jx1IAecyqEMwPpvDY6jKgLkEjYa
1XDXY7y02RnFHSlMG4OapLbvBkMC9fps5HrdCEyZp0+xH3TwPcnoDAO5fPmK0VQr
kYDmP++w+Ed9dHIs0sOGvj+DIy67gmsGeozEQURC0zErwzNZ/t+YUMWvqnk+8vL+
Kp5LKydlTcXLYr0WxvOEGbR0wlrV7yLJ7YCVr+J1eVsMPXnkYJRJPta/ifLSBOBS
FSBA6gb79tUsZyuFBos8herClpSeRoQQyaU7I9P4Kh2OX3TuPI37t+zzHiWbbuxH
9ixYlHEVxjEPb7Hz+4ej+SwtvnYF0Sxsx5+U3tKNWz5jW6zkke212/XR0C1MeV79
7+EPUp0CHLaprNyYqvScIQGjyHOe5JcPbkKEQJQu5rU2IOUL5vtU4VaaBro6rNAU
ceZ8W2N1uOfHHr1RgB0NKnwg/De8ya/Gun7fWmGRFTVdFoC+Lxuyh4HnCNdoYRLC
AHsDL9YVLePPYLSkzhm4d9fGoRiNUs+IrGwK1OAxd3eiF+WalnO13P4QK7Xn7sF1
nZgFzIvQkwNspWIVz0xfwHmatGKRqrCdAMAtf31mW0bTpSmCTGXvbiiVKbd+Fg2D
jien6MrSHQtNlqevVboEp/93fV73LgM46pgghetVBiPamZMIpziKXBqoH4B/9YVk
qgFsE8v4JOeWlK00j54Fae3Lwus2GHj63jt8AjCr4qyYlon0sTrerqkcWbdAuwN6
AjtX8p7sRWVy6wDqUbIfJVOBJ9DH2LyVt9dsO1VFlaafUlcpetJOxy86I5lzinUv
M49OEPhzuPgTR0YcIGejDKdBK4QiaHULAseWXrTKWk3dmpCakBbJgOpp5HtHQkFX
O1A+9EOBdrsVjZl7KffVJWqfjQyESDfa4kej4ybHo/MW44uf6F4qEghJvGHhmyCz
PzoxXp5lGWraFwU7/o0aReb4LjJXRL7kfBoG6kY54Jyoj8ruftlFltrCW1THW1aR
pN8EVfaq+jkJDZL0SWzDp5fdifch/E67eD+CzLhZPVzsZlbDx6lftFtA7I3l4N3a
3WeNgJbz0y7gkAD7DZR1iyc3yB+FPjM2sDempsi3sbcfnRl//QSufWm5EzE4DOiY
PPCDbsvqdDRT0N7o/UkZmkMn0iBSM3I1hKkaexE2AC2FbKCltqywpwwwfVObGyTE
bS/i/XFI1q3FcAoaKXeBNxFDjAddf7uhB638j0PHbL9XX8KUZ+TGsB75TLx68rVn
ce2RDk8FkZX1U8YhHdxIjdRGsTX5xjkdWRoul0uhIlT9b6/5qzEoigmH6IiBbFHy
1n8vBcpPT+MNxg9DYxMU6yNvBgplMxrJi/3XgEl4FC0BNJ9VwCTfnaEKtFG4Av60
Drj+VT/dbXU3PHV6vucLas4xW6S7OLv5zXy5qkuk/eFFJuM+Sy1Q8OVccTXrE2Zt
hD9iP2qefpXEqKoN0/YDjWjhj5FGPhRjb0OQeJWuUlbH7OAa3g55a6bfdcggvUHM
aJo64iVTk/SsOWgxc+K17U8uwSTgf2es1Ns+r5fZrpW1p5mh92xdtG/WPqVLv3ky
0cpnyC0d8UH4QvSYJo0WFYEaMkUWGHvzgV2E84HTo/dwnmxK7ARjmqtJ3Ov1VYlb
Vt/Wq54+LGi37vczT0YKfIDHqKmEebAme+UbpOr3w0o2YRWHKNONan2TdG0m+uio
+a1OVEIuV+JPfFmAZqlUfJGlhMUzocogPADduiYE1II1zli/W7P5yofQsPmiRilN
WV04SRg1bGzcC68pUfvSMtfYlPtMVH6Szat0pUWUe+igP7Uj43uMbNnw8P92Qvl7
eIclbd75ugttNIkMIa6N4mJxvRqvR+f/yXFgb/2GB0Lon392Xtm4NYdVqTt2G/BO
dqnELBvwFKgb/y7W+ncBSSIBFbwU/j/YKhB5RX7b1qiUghKBCq8TtsSjbB4CoQFr
m+D9I6P+TP3H4rtupyCKWtSV5aCfsB2u/1ovhHvgDJOguby7UNmrCJGSiOXnSzti
VjFzaH92+v7KhdLxcjl7X0TYnEfK+ciajQ/6yf61129bFtuLVg76eXkMhefblzb8
mAW0TNcJsnEWJnE+amO9o3JpKRnWbcpJAMXzdw/GOJE/ZT23rA0w6f/YHsAEQsV/
TBv7Haxrm+mkZo6c54QQrW8qcQwx+t9Dsfx1N5QFImE8GdT7il2YTIcWs64htaVb
UoEUE1/ALopZvqmGiCHakPN1tV/C+2vlaPGcmTRnTw6b3PgjFHtHiy+9MFgrKxtI
xUMTG1zntZrDLkFbv2HxsO4ckh9YFx9CtgwP3cax7MogmK+cFSc4H7yCBl1i6W1c
xzPKIFa2nVQ7cSp0jnHBjOQfxIEg9zRPcwyhzTvnyRvnr/feK916fUiJcXtf78SV
N3NfUC1Tj0kpXiNxoWw4iDgcBXGHweL3j3V+r/co3fgPiaL7dvBE2czxb9s5BVnh
f+EITWqK6MF+4oCgQZDPZapdX0Igt7gsS5nwQ51WuKAe/Y0ZBKb09nxKNY1evs74
bXjNUUImZ/8M0tYbHWRzRCFnlk6OPpaMLY6N+809MMHM3UnbHiE+ASfawQ60CqET
HkkWdo3inycPfKFxdYSSHNcjvCrMb6HB0+4bYik7E//EDWV4k8h47IQy8CKGbxno
wmbTdZj+oa4+Tcl3bZTxmfeZus2HlOS1+OvjvHr2DNNvMYHNMv5dVApvkPaolIww
10Xs8wimI3C1baUf15MK/DE6fHcOpceXJPafvLQ+00XXMv9OBgZR8pp66JqxDF3O
52ySVYiY4xAqBCjiPe7LHYPez2GhXXVs+v+DMbyWXNlL9xhqciWbTceDJjf7DEjY
y4ADALYmpNRAnIDUhmU747n8VkPdYvrM5qoiwjpSZkGEK0T5zlxHSZbqVKVUHHw7
t60OfJJ/6muzB/7P9bFf5+LgfUNgb+aK3MMQX96/F8eL7iUrMdMve2byL99911pP
BTmY6gqBsdKMy4sg5d0bmSSNhfLf1SQf7yRImstAOWvywpl2z0k/Bq8HhQLL5cPg
KmH7UC2H7/EGVMZfzEVStBLixv9O+blg0cO5dF9KmvBGN0y7RqAJj1m0+gxoZE4C
1NFzmFirF6rV+IQJAeMeM+jVaFbs5jG9AAbJFoPTzadOhE1ZBNBol8c9KUep/9we
Li55DiRLGTtjIIMUWrb62QW+a5ikB8PHihnmEtsToPbellWlU94RHjsSKAcKP4a9
E7QE3EBTKIOxIXqHGwh93KWa1/tgHL0J/hhZkN4IsOkBkjxki8lATSRJbur9nkqd
bdqboFgt4Y0RjcTYaExhHT5HfkVDGSZ4ofSMkvqlHKvQI+2as0V9Uw0ROvNQ0nlM
plgMPArTMwTMNiJn48BckWWSbSRjuZJZrtJuXMWuGV85qBpBI/MlU6hJmGcerh6O
7eQ22OJRi8lB0+F9a+S0prGuNDG58VAx1ikWFh73sF9//JQivfwtroYvLpSkYpNZ
qlVQIaaj8akvHGb41ga9wamV0DKPB/uOZPCC4aFlRpGI6dAEga4xkJqp81NH8j6+
SAD9QDiDqMlXqtCrGKZnL7wZzDDI5n9seEdmrH9Ol1Lh7s3DRHzWxdpoijbE0oiE
OURPSALdqR7Zjxz2Gb1ZKwZAY90owZ4IQTcAaa7scKx72/G/yeO4Wza0oMW7L2J3
c/V1BDHlXEdy1vGLW4d3nZfa+wbLbsthKj4GeJ9lskVLvFyAD1acLyPORfKoEFfu
jnNRlG0QaQgXKVVcs0iixnNk8UyvlKabHzUrAsYeM2KlxBWEpbvIJu4UIJC6bwgN
sJgOuDAl/L4q3m1IBPiv5nV6uk9clc/NxQVlqOjmzfNLtVAquERIVpzSVqLHfaXG
wYgmlVX9llkGPZIhUSpvb3peKfbyaTpNbgc744L0RRIO51kium5bRd84cUEGcd4F
EuuCLvlc1dpYhrQfY4NAA9VlbGUAJJju8QMlMt3wBxtYtyulacjUs9weo7ZGQhXt
6khyQzFeChBIGlx9mbbGktb4TWTTivTSmAgzIcuNa/9k8cO2H7gaDi/nW+OqrPYK
rS1nEcoJqusYa+WFG6IOaxEnyKyO2CJeKqzLf/2N2OaXW1JPO582XPtbNXNPFvKm
/KV49fo9Mm+hCZTdh6G7vT9aPOoA+rbBl6gThWNbBiIcj58zLtaAjHRkXWMHUlfV
d9J3Ql2Adc/U3K2KX98S7DZ0RQLZnPzCGbgd9zfDhH4F0Lo4s27ClVz0asialKlp
Mi9HCPldDdo7A08IF2d+rtuqQ3I3leEifKAXT5TpaY7UVDyMl4+9fjlWeQe0Jiye
qZdB9Gn0krCRWmDXiRQbO5gteGoyhvN14vVIhJsijUp3ihfF6hny56DAx8KNRJ2N
gD/TqtuHiBhxLOFnv8VCJW4pOgftfVjlUUSb9bpElby+rzD4j0oU65fyXqCNriK9
A1r1e3xpfM1GE2Gi+r2YKCBUXTtoZP55/O2aogX4ZB1R8ZfCWS1yBBWfn/YATA15
oDzdlYKKHWeL+c5HRngFtmNCqmQbJz1Fvj+NCYglBmNOP+BGOyL4z9bO8He8YkNp
xND9vt+Pyezno9/ip4p5Juj/Tlor8Gmp74HUSD8l7Sod9v/eRe+krzLLHHPr+Q9A
VcPgZgjzhJwBl2ZK76eQPVM5jZdMpnPQjPWqFijbnSbY6avPif5PmXuFui4EnIOf
+XXmngeTC3nxVfc99ve3aAQJo9YTzIZgOCiUfbYeeVpGqzHLE6DpoCLgrVCWi1uS
KwCJ8VC8FGPT67YrTYI9kO69grbuyS7wBks2q9T6A8Jjzh7wwQdQNu6rTawFOfIX
vHq7xv/zwqyZBFClIUCCwKPgSPUjqTJJavgb/IwWwSyFS5WpD4UvUFH8xUek7Pat
PSU/aEVeAIQqoGqJCWtceY9xhNWOLbsCS+Out9Raxb0aTwteDC9BPnmh/MH2b1VT
UQAdYpy0WurRkNfgagvBS097ZrAIVsELZexLYeDwwy7zgStBepNqRGQxuHCkVa2U
Zb1dJdXInOV80QXpabu1dX71rsQWo17yBlJyHbOxKT2ARAHem50gzjLHURyDvTOc
qWIXuf7W0d0fn8CmAJO0F+3FguX78sVnWI6HGhWpIGW1Rl86zDuGwdg4/ZsLL+It
xOxCeRcqfX+15MBBLQIiHfeDr+vcFCumKa0mq5OI7p5ioa30rISsRVFW2XXLMi6e
7m/+Uk0Aq2NvAX3gcVMpDWdUsznLYvWv/7Xqq4jpisPzFpuO945spqltjj5V9JOK
hvEeqmFou2PVRzSf1A/gbI8LFuO0Co3xejUQVOLG4bwGT4WJ/P6ZWion92bnSkQ/
vrJp5BkdQidfnOupBTrF+gezCvYFY/rcO2rAcozzubrClj5bjCLVmh8sKNk4bM1V
gE+15Z8w5hQxGBZixbentRta3Xi/bmLpFf+s7JpcfR75vdagRUqyNk9jGww0iKcr
T7eM5FU+NLfrmeu8/UY7O8yBjwENLJDjocUew94AmMw07J9AgFZEf6RgqGVuWuuw
HJ6auNzC9KcqSrI5zaKf+9MEpFNCdakIGbQmJwP65/yLP/oYIi2lge9AEl0gWvsw
dKSVhoVaFCY2gTOqiUNqmzf4V1uk4p2IDdDCCtw9wDAnsIU63EueC9XIHkJjX7iM
+haQ1whnKcNFLLxjMSpOvC1RRNTAz3L6KrJaeJgosmKiL+MJgxWMXNvxmap7+HAE
rjwM8JQrLk87dWgH+emWXn/9k4Y8wZUIbkCcpY99y69I3OBJGzZk3iKAf1saJktr
Q3+06Gz5795GHr+onM+Zeh63R6izF1tonhpS8arBoFq35UfaRh8IJTYdcLj6iE8K
WJK4ZqMJ5s50WC/EznbBrnmNyqygqe6x0xC3NAaAicgMLwL5a6TAnsJBmALwKHbS
+DyB6ZB+n3K87M1G88LW7k19C1cINix/mJhzPZLL+rjOOWFqpBkmjY2F2VVXme2s
Q96wcpDYI0LQ/l+1jcbNGT7tJ5VebQRgsGNCFEqvNPrqlLQGi0V3BNFCrqqRuRGc
s67gsK8xI8WUAMDP7HxjHZSjZluyRiuxI2fhvWHW8ziB6xPPVAsKQyqGCcnt8oPL
RnArZfOX4w4fVQKFZd8MtpqRNKxpY9gtO1xYwjebO9HeOALwZjyE0Lpe2ZcDk2Wt
ys2DtEMG8DFiFjw4tsDMJv8tqpaKZAxekWcvBDLwp8zP7XNUeGTVeabwtrjN3W7P
QdJbYrKzHzZ/YOHPxvBcevUUDWokoBxjl40UCbSVsELbtDQgNRhw0LKrG+Ni12W+
Hl+IlQ4PbT+rS6Poh/s3cH/YGx/JOOhkcn/ETToAWw6JshP21lFRy6dZE7JZ0OIH
uldczeCIDZaCZFhjWbdaeMH8t5GvC39smmN7sk2nKdjCgpLzAlOf20AIjx3FLLWm
sMOQP1woWKTTt3yZ2x8YJYKO1goivgYVHNu5dlKi6IfUBRx21WQq0bs8bybJ0Xxk
THNBuYoioIjDaIv4T+uVZb+Q0nbQ47be7G1hqfjXYrQiuFJG37MBqb24RLgHfZVW
fI+AEiRu7vE3RDRo3ygT+Yw8lDpQ5cMrI8yklWcxJkTlaJ3Mh00IC0tf7vpHEVuQ
3gno0/xnnfgHwdoJ7WAcgMQTQEWrOWjNLU1VeHNSKL5tTyQPK+TfVhFqhSTZ15g2
yg8wg5v/7tODXyavUNg6Dujh2ytXi1gRCQSlYnwBkWmeUDfy9VklrY35481G9ZxS
TcKHGV5Er/kTVrxDi2qm0wRJmTD9U7Hdr7Bkn6HdtVi/cIckN3XV8BAkyIZJSQFp
0MSz0A7YDmKz2cxx8wBuFOLLpC3L82SmEuZeWscSWhxwztBnfhkdy+27IOOmSPGS
a6TmI9ewc7kZW+lqUeZroJI2MYQag50607vhG3uEee/Chd6HVY34ow4j/inovE6X
9MolHpnm34Q5hV200rlDxsnzmIS1IVcWzox364KiQjh9y1j6c3TfqWHJp56GVUDe
VK4knO4jp3X23Z664iNQ1gk1Fqws9YkBQg3qNyWXjYqqLifjph4p0nRm7FBBTEch
Gam/QdTplrBmDZxSygM2jwaP62YVP4dGXGDX4lIzwQuo/YYVs5ZscaMOfH4EwO9C
qXVFhgGwQJDtx/oRABWGv1UScVPGg36D4QB58bH0IZpCRu7rjSa6SGzLLsU36TSB
gp0XyCx3pmd39quDwyQqNGGDsP9mf0B7lR7BZuELBCUh6BhfjNrhjYA9gWqqcfnn
mVG48I9rEoboeL7hO/SbfctQA9Vfl4gnhaOtFnmFa8be508RPE4UMB2XbKpFu5PQ
9IKmqgbVFOv16JguzbpuR07wjPwnJFVTQKGFPqvmwB8oGLXIWeTPfw2ho0fGAptk
EHANfIzBkv95CYIbMDZ0T7gElE4NJ2P5E8KdtLyQ+L8eTVGbxxQC3aszc79Gp9iE
CYOEYYdZ/nCO+GEofK/AMrfjVnUEncmvDZOu6+JTbOhpnN4zPWVwveAg+wbHTavN
H/3SZkG7aLrfCaci3wBNPCPoEf0vowV1X7K/ML2gnzT/PiO4h7HL3wTAu+ue9Thg
k0ODnf1XTB9jjxxGlHSn+CgYHbOwhjSEQT/0evrkW2HGypBOzT7zev6sxtxnI/nb
ZYCC9QpFZGVNXSvZQpxp4B+eJZhuzxIpP8CeDq8jo2HJRGzor0tHWLqIuKsEGiFa
fTICNpWnYD5n+2ELOJ+66OjMhw/gjx4sZLEQru/NTA9diVKOvERIEQfvvNO3VkyD
WJApJvTGukrZC4JLSwGqMEfPffjN2h7iYfrMgDCq6UQb8kKaTGaOS1s97PlgKXB0
DZAiTuZefltjweysvtFKuHzf+CjoSXf1e3xQfNtOGR4TQ+dHsVqqxUQ63ES27PZd
MlyI8Z1cDAnRn+AsuZbYcD8qmaf+J9GJShuvcmH+eqzBLY1XANOZgectcdQoK9Lw
Zyqg9+S/X42qEx8+GtjvWAUkEG1B4iVAiskdJ8NYoqO9pGX6fGiO31JNsD1WS8sF
smW7mWM1heI6tXKeSwqJIbMOtgc/F0E2t9IW6O1EU/qsCvdtY48wluTTTo07i3Ax
zGw6fkWEkvUo3f+yalL35ruu76X68drg4iguVKbAJZVSutuqU1x5PQUi9ZcdzHJj
hNb/juZGSsYcsIFfebrNrboNjcb4c2Q+sbvcZ3imY050lThJJopbKMKemyo9IkuG
X+jitEJrTVModeg9EAK4Y5Yx2mZ5ylRQqswxZPUeQLFsR56UiFkKAvfkSTGbnaPm
pn5AMBpGNPpJyWz5HXiE31xQeJcFQ9TEoKFwzVCLfkeFcmLf5MQF78JunIgScBNt
xCmk1Cdll+8Xg+cY1LccyIjmrH4Pxdou/oDjEaogO0hsqjhlCgkk+MLoVWe5VaJk
URRkHt4Sa5mSzivsDLW8uFX5K5TninjtRx6tP4CRMh32e7YHhuxY3r58FgUpU/33
SsyJEcGkvOCaAWQHMZgxdOh/nNmsmAx6h6wxjgYC71bjBcTZZiGFL4RoqH5SSOQ9
hwH6h/v8KzC4T2kBEjMVEjrvchWALNFgxAWYpls53bicBTf0B9VrrDHgFLvCcQaE
RbpCuTUAsd0H8YmFFxzBLSGhJmRilJGR+Tz1NTfaDvOL55b1o2Stu89GhW+H8F2/
iF+cJCF6OVsCsljLac9QvabIbHAUTF+mr5tzEmjEtF8GCHxxwoohUvFWB9kU63cj
y3KrUGiDHVaql9qmYpJ1D6dlnb7GHLuqjRfcXD7O4hhwIQ18jl0TBe+kTIr+uQ3a
ijyigwGXmpxX9VL81znnhOHypIIUEkRrKINW1zhLC2FRG3ZzJciQpYYkDnKMn+0U
hGy1imZgS7aTn5WP1d87FHlrb7vVPmmsk+nkzhyfXn61F7WVNMJpDW+/lfG/psKR
pVFQ3kNHAS9ii3LfLyBrUNAa/u7j0fWy4oX/7pZ+jIL1KnbF7zaysmV8oeTM1tGG
k31eDY6uGtJTjNN6WRAFUCf3YQs76noaSrbTa4N3zpnj2LKS+m8UfTAxflxXx6A8
MIT/P9jANJZl3evr65guPMDTDgdZ+wf966yJWawZGHTtsYqn7WM0X8fkTrbqhWUT
yjPmQWxxJitkijRpDpznGvX8bVn20WucNspiuz5SqjVexRcSgfjYftz8bcNUzZts
CwiMr/tcxv2cXeBJUnTw3UyPD1SC8S/fGVQfGqvtQYe+wYBIkXP7S8cbAC1y9urh
+py6cNacExf6BvF3lN61xsfvPV+jOisIdQ3jmU3+J49Vw00wOeNmg1ylJc5xTq6v
8+pAGeQBQCuf9ZmVPyACx4zmNjUoAvHrkYGSNEq2PinXFXHfcteLNknGSnsgCHT8
+6It3O6OVsXwgmPDmEfkRSNvtPBLr2hNZo+ox3FRlsDWee27qPNCTiU95zhZTT4o
mA8ngv3Zia+uUYge6BOYX2yv2TLCNPDZ6dWQRo+I0APJHY1UtCVFYo1sQ4E/GWsb
+VdaVgPVm1Jrv2DiUXUQPJDIIWeMrtiaaKImqNJMux2jh1ySPnecj8b7T6TLUCVg
MER9qRP3CmyCDaCGNXPjYcip6yOWd/f9PWbwb1tU66rl5uWa83LiTAiwIHzllDm1
4skgVqbYAjzPDuOSOz0iX7fUyEniHj6ax4NH9xxO0f8YdoRYMtJKVasacYLT6PDD
dSsUeuzfCT6YrTDeiqQ2vDI2zJ2XCxqyT9tDkGkGlyWc/hsnRrI3JxL9IpmbRgSS
VRS9j68yQtch2lLNW4c7yjPWxO8gR1Ymmq6btHRhs/Nq7NKkjx0rn1tbkLOI09jq
dCnUr6XrQ9FjFgrXLBr0vOYfe6/cN7zn0e8koeG8VOrSTkwt1OG5AEJjFJCIAyWg
KrSeosjX3KiGqT1Kto+9f++cM1wKiIMq4mM7lzKCQ8PRI8P1jrXK+3qMveVB+isT
/TNnVujOfvhaUJi1bl4sDA1/Erz9agPUM45aRmUxUHVZ4rBXjX99amLBtDjMrM3H
ZrqZEjF1CW/QI08PzYVo5v9V5lNmj7QHL6KD0npD0ymsGJt9ttmEh+m3J8S3zQXq
TJgtjIOQEEWr7oGQj1Tbldurtnp+eYn7F3jSkrzF2xMujPUsreN+/UwJWERTx5Ne
qzxImmV7HjlOav6nkq12KQmObOI33oBUL/usAbg66C1BQo0huMGmAAUz6kkSGI3Z
B5R3DvYjmWmqVDaMnXIwXMQVyHlv2RBKr4rtuCODFThYiL+Pw0/VZon1SyOOCASt
pQVkiZ/P5ks+sZoGgQFrli/EX1yjUdkZsXQU4bKau3pQedFwKf41Yw6M9fDAkGrV
leb2QrVZDDCGULRQlOmI2i0y7Z4GA+GDvB0Gf0/q3hHAZqhLhK/NcrRgkkll3xl5
WUpFrmEel5/MqyjHpDkq1sYkSpzRza3jaqjXBCMYydLxSJadaFhjOUNjClokU6lU
td8MP45ni22n7/Q/yJsncNBOkz5+wo9dVauQhKs/FDdiO/pmmKbogcGBWYNlFZ0f
6+xknQz15oFiKzCpvSFujjVqLB496PwEOF9nxi8QRnwmDYCXIH/HNr0lslI2Sw55
440sEI3Cs+FEcVQY27kwHUe77ZzoIetFJp+9pZCoVfvSCLe6qXnwRiUCvYNmMLFi
QN0sLVIhEjWhglQO5ejL1+KyhNcKjlM+EZwpU4ghRhaCGXCXARieX+t4CHLdP6Ob
hP1nTHSLtf3lDPb2OXMDe1jU/47NcrA6+doEkh91F0mi1qHYkKqFvQbSjBvB2p+d
xuqn01Z4aPvNKhlDxEJtD8i9HLCuTguEhDV0bY9U4xWS55VVJ3o+/AwUgSoa9Jyg
Moufi4dUsMScSviZuF0y4aUnDBi5lDilZ/vg4mZbOY97/m8jpr5n/xyDkxQuqnUT
1SvqhOOAW+yJj2208Q7/XVc+4FsJkvYS3ZXWBtcSak50ljdxzYxDTa4K0l7vgPO4
9t1eRIfpVqwEEg/5BN0bGWYzh5CFV1sO/rw2219373k+lGFJ7MULRr5/b15MfX5v
0aRxwG8IBDa4IVfw4x7rPYDGs0RVyBQO1+QeftAvy482XkQDbTa6kpkaa6E33JFY
71rYETvyvSqxh/ju7ABHH/ksOx9DarYWFS3MDw6Y556ABbHgOKA30AAEL+jI6ZMO
2TmwkNBzVC0+/rR+KozuIwuoz+b6h6vYX7fqrtJtDsA177yQP0S5sGkh+p0dp4TQ
4/IrGvtudmqT1Bkch+TbWEa1BveBPHa+jZ840mLXTD4tO2O5+O/CAVjwwGOygVMq
0I0O0f0otZ44rESFENY767WpDEfVCSF3P7RjEiE2hVeOf4WRRcQdHMwIY5OTwO4i
XJGxgiz6QYrAybCy7X33JE30c+RqnmfbQc048tCQOgkncZQLWscKEmSk+x3s2hwO
dGind4dtIePyZU5zleemElXwq8+Mwz1rUgSp7u+lV6kVYTyAe9fSmX8LLlk//Dvf
3jvXXDxffagCKosw5jVfGxXynEauqM/PRIUFxhW1RM5L2v8nso0sQpkLEw/3lPRF
5PkXXOMjZTA5w/v/5vTGj326Uej3K1JDeRhYzYO10didl9JqkfgbWlf6MzQocyjq
LZfGSxOqKcmy0nu7cz6YcNXD47vTGwLOW0jSd7aEs54Y5+Gj4xMrq6jzyLUdcH0u
nL+ycFZdsptJ2S2LrmpDDST3aO38VSa8a3yaejlQ8fuqEnSieuP1N8KU93DjXcD+
wSA/kCqDesEzxALaidSp8Ab2lKM1D+5sM77OXm/YWD1kyYvdtL3YyQOY77mGmuAq
3JxaDrdNL/sX/b4qhHiqKWL9CoPJ6j6pPKoCE8zv48ITZcW21YPi42Q4i2FHomit
Lxzf95qM0Px/bv9Acm30giL9bKK6n2vKnfuXLwHrHLB3c0oSOrYEYOCaTi72vNAR
odONRKWFNCpvUOc+eTS7hsokxB6Acu04PU6m6Z+QeUke1tf3s7CZHTpi68Kx+uGA
QNjrSNz+MpqjImoUOSwjLm1hF6bZYW9fd4xehvXXOswHsEIXPg7FVauHOaytb4SW
WHBrsOU9erzXdz00GqXDx17ON1hZSK0uIEc+TYLETH+A4OSo89KgpZrKh2OtjMxo
xQiwMwtDn5SQPOQGpv56nCDAPd7n8PTIVzDYsi85VXl0+0tPFn1p0OtKe6+gIm4T
U/Nq5stR5t7UME/esdjWCfKzzgtlmYatu+ZL0786JFCuuCoLninTOGfft6q1EBSH
VGcguQkvJGITObTvvKbPgHU2Dfh914aT/tCUj8uxPE45c1HNE+zV1drB2wTCyhYu
Ex8Kn7nXOdPKc09mAtB/QinXSbHsmp076liHEnsqLQhK+e1p0QI4Q813YPqrPkdh
vCHDQWNxI7Bk6vJjsfBdjofs+5s+xSokPGn2ZF6FmClT8Nf4xrbHgpgjOaJhYE60
lXdmMZNASzK1Bn5j1vaBdD3lwsZCV9RniCXckwEwSGm5PjN80sKMjyd8jQKjJomy
i4S5YAoSKpL4LhPHmWnRyTCvyqqBQqlTtdJx6knrecQdoOk2Y8BkDAABIOSYbwvM
+7qz6aBynTH+vlddxxHK97tKmaw+9RFz2kXevEGPVO1r8Dml7hW2HLVokn4CMm78
JlngR4tQwgi+9woLh6ZXyiD4xe1bZdQGlINgz04SIIGG9tn3/5SCt1L5aqTOy9VV
ehAhe5d0Huxzdtx5qhJ3EHeJo9POjWLWLUuak8IoTJ/vVll1lihu5kfckMPR9o3a
k4KdRpRQqNIOecRoekZ7pMXyQa1uM4q2/sIm9jSAFkRsp8uhxPc0P0dE1LMGNJvr
9Jt8qahVO71frk0qKCKNRstWczQXrT3HND7pBkXKqJifp9GGHYtJcCmOXup7lL4w
V9s0VCExt8nJudpcV6zAY8qv7e9FYwfIKlfgRcBX5hV2GhwH8M2JfKZAfgy0HyMu
V/X/p73Q10BIbEYYfUb2PmtWs4ABfpwKnaMYdrDz/O9iFYF1U+t55QlKdvej6VFG
vKGKEXLJc2lV8WRaMF+AaDun++bcKUh5PuBHynM4AZnTdvRXlpgcv9vnUJ6xb6Z8
ny/D3xVYspIWzOK/PoibbtUFPcL43Z7fLD2RR4VHnSa5qK1GvNJUlaJI3SGrviZG
nS3zuz3rNHAR9uOT1GWYXv3ch9JeLvPcLLwLcGcBfmvfxneO+1Cnw+2l+ehhDe3X
QNjfmuPgdT6DZA7cfSQSPv1FD1ywTEkb2/7OhxLoCFKq4X0xAqloAnR9xK98SqVx
ljsu4kwluhpI7HNPqRJcon9QJCi2DAIUjbMntfW04Ac/xZiMoHw/qHyp8F/TB2Hp
BMqGaIm4aOeys4w7Xz8VVb3AAvFJs+v70E/4sLBAcq2hEBbUTyIrR4u3F80byPXV
4sA+/90MBHuPnYMnPT8AB7JP4HdYx53TGP6cAzyOWrDPC1vWrzKfQaHvjMpAn40r
7KpC2ToHFlyOASeM3dd6YvL17Ta/9POmvq9WZJ+Qx9nsVK8ev0js5h1CpPlMaIVm
7ctDyumwHgkf0LYRRTjHg5k6PUnXmiNN5KCf1AjMy1C8HadIg9IvtNgJQV6VFY30
o9siHu/N3MqvrNkSFgP0FewHzYhZ6wSDoxqDOTspuwuKHKeUmjpfsWUYRunsDuTo
L+f30tPtoOJfrIAfVmw7ORGIl3w3mV5Wi/jGPTJ4Rlac/KozLBa2Anz8JmzB5Y1b
HnzsrnrB3EeqcdTxHL+uloN/c2mWDvX0day3HUEV8Bc6g/1eH7aXvfoPzZ0+9Yyc
Mglha8il+NK6BoAq0xpSdlSQ6Hra92XkhMT6NVdYn/AvUxk7fAvaJscn1MOINJT1
cgyzpH8tc7wCRiZxOlpiroOLqHTIPwUqIEdEG7gCKjBRjvLP7amEJBPOSjg1Ky8w
VFO4OAAx1mueEE6zG+KVb/ItASyxhXtNUeiYKZnZK5b9Kdw6tPPXUtjw+1AZHQ6j
5ynSydHPvBwF8dOJ+E89PiTWABfn/BmbMOLXetb5wvEOkSiwDIa6k166aj7Bci6u
JX8L3+XWa9KAvDAO2d10TQmDiiThspPjcxyfLSmpmG1M8zsoM/3Vk/259YFBKtJa
WBL61XG4x3YYLSQBOKg3gUB9+lpUPpcPYYun5NQdBpz3Otjm8lyG98DZJiY4OY1e
YVcuoc7C6QIJ+FJZhLAJchOJ0slvXRpWyNWSbllkGOqEW33qK2I35fbXfHhRy7w3
JJ4uVLD9aWWBq9aoF4qKTOgnLFIxhV25y4wN3O167y9U7OhDOw7pMAiL7Htfyr/y
u8cyTphGMMs6bhptiPF9col0qEhCV4rSX7NSAEQCaKCpnbDcs4xDv9TyfufMZLaC
LfGVxVwpcwNqYlofYcTj5jBhtB2fFb80/rrDiWu5l6wkDH6++k1Ogq4ZncogSjOf
DUtJUjR2t8JctgYbtfIkzc2C0gobFVgTbiWZeCk2T/uR5drxd+mQn7hlzBJMh8ho
xVibRRcKC2F9Xu0Eb6l5imcQECRpPJDuEAVfHjitZdshHL5DuFAchcfZtPXiiE5s
3Ls5PIzj70MlaPTV5sFU/UppKqjLdlk+IYg2jOnWEX5MqSXt/Jz083LT8PvYGCoj
2isMXKYNqyWcNqZRM/88HnDdcmRzg9ZaoUrHws4eM8a7sFr5lNmQRsmrcesNbzZx
vTxtKdWFSfUncYKtuTlDuuF58/8HTdddVjJfhKTtYxJ7V/th7wSvVYlmIo0+VOza
ugtDVCnNw1cmOq5yF91ZQqjtxmwmsNJb9I1LU9Gv7P/t+GwcTajdcly69W1XmuOa
OephErzMYZritaROAFHeH6b4JfeNXhgHMLZXe+XQD28ktUyL7+g4hOxJ0r80NxTX
/Vyk5/CbMCQJVLVS++dQFf8yiR6wXsN2izHgRwc9HnW4rK9aPa6hQRYojF2JDXfE
FMugQUf9yGfKUVpIbUlHAJ9kHWWB3FvZu0kZY8SEAjY4ierq3alnF4PCzn/iSg+T
2A8HPURD9EVdEQRfhTYCdg59LxOot6vxkXqOsLBQPYeDrKsM2Mw2wxFxhKE3XtDU
hpYTkgF+TYBN+Q8fc0Lvgcm07u/Kyf+OIxZdZKdS9i1108jxN2ItFJ5RB049Dalb
9LPOSEsoIlHiArmqxVV3OiW7HBzwFB498xKPIEqhS+wHIr4ernH6HuugIrGYFm5F
loPmeUFl5MrdbnxM5Q/kS1KveYEkbJmG1u7p40ZNNfPYwUkbqwayZQFSapeZOFyE
Sc7RWnnIwzywrbuyIAwb4trDcKl7S2qgiXA4ZTr4++xXjq+Nm1eSfkSnPUndSjoi
IBs/PDagRk2rKeHJyQGUwwL0QCmC+yWcEQSb5xrkFR0pVUwXxZDIbaTn0MxJ+bh2
WajcWFdmkyi9djA8L6BX729ifHOTIHxsyxisKvG2mMakQZSGjVr7LngorMwiuTiS
c67/dlAepgtQoKXtTIyb+VcCg5rzv1bwsUcDEGSZX6xuXsISEojLvr5QQ1ufH+4a
r+zGG40OTLmCo2+QBZizr0wY5yF6xmfLBDUJp1Ob31Ck6cRsO3EcdKdjlJ+ZxfZb
VCGtVBKKZDst7En4VHXiu1rwNrFEf9TLBKsc3EpfHbuH/FVqAfI359EISNhGohl1
ierQeLaXS9ktPiHnXeMGT2zablxS5oBlNDILhDy08l0L3KfuxkyeW/e6XtUzowor
GN0YLHS6cop4xDI+3gGnu8Ce2XVKxR0wKP/N3FgIPAFhWYT8CQkTXtnpuax3RVqM
YKcwV707FufhlKcTShTnimyBsvCd+fwhdnu6X0rNaSfcH9LjLV9jxA/074f54Jfb
fn7insb7wyzpiANKTxwCJDpn5kZiJPqDLVUGRvyo/ve9W0Snf3qSF2orMuYa6NUm
009/ApfX7a0HbE00fTnfdIKqpoX9SIwK0H3ocQu6SSECmFZ7fqJ3PHRbMn5vUZzY
az2wkr/Wdr2Mv40y0kvnbOqt2vAxzNDQ2TGp2bLg+kCg5V2SwZ2hwFCm6anZV3uM
4YI1wmPHrNc+lJP4S2P4Kw4qosnbUvRk4bSQddGf/Q9VcUTdERTGyoghk1qi1+xG
SsUiTKc6+Vpz+WVxZuf+f2zr515cgBlomafkzszEKHNxDitWOyD+anop7VyU0B1b
XsyL85sEqH1v6IlJvg5E8SykwFK2r8nQj68DeILQWd1N12U5ssXfrpdwMUO3PCpy
FOR+9doryBqb+soycjP3eG/UdXFAUeMhi1yhbkqD/txk0javkFUOXp1tZJjiyE5x
pu4JeKXs3hyY+c7cjjNXOIM5a2bVfBqbz3fVW7kBbgEsic/v9+OaXa0B+ce6soAa
CNcPXt4KL7asy5tA3Seqh5cjDNjvJA5fzr7/UvSgi4bLQeSdVVwYuFjFaeQi5kpo
XjwXGTQ84mYAU8mbP+glJB0Ga1FVnqBBb5SllCOS5CmPRUjQXmvh00C88tG08zfY
kxbylbiRX+mjCmndZ0QxNQXklgRy0DKBO+Z0yBr62i2YMk65asMz26WurP18xzQc
L8i6KnzaGbEEJF6Z4l0Z+UvRKq9aYFGPJ9sUYHoBYhdc5GcmDssV8xOnwF04LGpN
KFlQ3BJ0BOLwk9YD+2LSCI5l1f30XTXNP3etktEeomaStWK6Id2yWK8M0UKm8xx+
q7PkUvfvyysr+VHKvcd+xuc6j3Fesd8qjoze9tUfi/BwFotKxfQcDf2Jbww0B9En
n/JL6IrgLQ8u82WhPRwHVHUyqGERcXGRcqm4V2sswPj0MiBVl9bRBBr/XkUcebx1
tFvUYer5Vp6Gza4Jjn0f3SRwV3nn1XUMn1akG0k0UFAF6adPw5tXTiNDDWFqHv3R
APPqFoqqANulIVGqRxb12LXyJnqUQ+dFfrfvuT5qBynTK+kGp0kJJaJcZPv8Z/JU
dL7RV99uXfOHky2O19yD1CPk59DcRlVCQ8pPDXL0ez8XCjv22LcyZCBvKmFhXXvb
sEqLEbwwNX8jc45aT3KnAkQmW/qxZo1v4hDsWJaodMl3SFYIho31rg3pM/rMEBSN
Pk5jRrp8HSRWiQA0JuaOc09VDMz2HzvosCA6D/P2qQ+vkvoAb5iEYOmWlBEtvhmz
Qrao1xyfl3FAPNrn1GZBrp6w7z9ttZ8mhjXgIp5NHpdVqptJN0c9Ts8ytfUOhDv4
Sv2zYEQRQOWeNGqPABEg/y+RYRskwScrDEN+w+jYeapaGRw/4Ewwszzrj9gnT2a7
HTlmP/QlhZcuXmkev2r6GXkIf0H3odPKkLmk07+0C3so1mNnrJl9Ejz2qXSAZc2C
tYGJCpGaj0+ewn4RdFYTgRFed1y7PGJV4tqbfopAfytwRoPJZoRO4+lfK8MI1Lt/
bKkkAo96HR0s+vzC6YrwEZnH4k8yGfybJOeTRkCuVxbbxJJ0LpxPg3u+LTkKS7+n
FY4NcBHZ0ncgoDowsc8QtDatg4Jc8OmClY05dnEd/Ln2gBhWM6oViSXksi9kuXFa
U6wvVu87CA/5drYD3JOJebApw4g9Xsc5+KqhwN/iSy34LUq6KrsMv5qiSpiNFiKM
RGt8uwhIovuAkLwj1QvPjIyIx24LBerLFI1NUYo2IW9JQhW9MMhEd1NL160jKnH+
StnUfj+mXnDADDQ3QpTPCmXrCON6J8SK0q6wLIIiyp8v+wtcU5w4RDiU04zrk5LA
NT4BgFr40SCHkJ31GQ9AA1yp+sWGtR5dwVZKdM2G9AMaBl5cLbNbs95EFRW577zF
JJhCcU4BP/JOb5AlPTdf9Pfc13mnNoj6zU8rUNPJRNdXvKav2Kn4sueWu/VBbv6m
M7r2+ptjqJLaeiJeGjMhgPo/FwVYod9UCc3ybnReboATqDzJiyJYKwFAD7A7jE4W
BkGXM9VOHOxnSjwrsiRwJC2BqVejpJjr8V0wermEE2KzTaIuy4EJficu4qp20A3a
PVLysx4PVR+kT1HqLfAwZn1+YYXC8Hh3t/kEaoJjXX1DR6D2/RvtiUOB7Q1UWP/O
rrb/sXs6jaW8+fKKpgXcmXs7yHmZbLvab9g/NRens3cGoMpaqvG7/e6pQStlMPPm
blffgAQ2CVT3Du+6sFts2Tce82iBB5HT/8E8dOF6pRLxIYbX8W94bb+FyAsFGWMX
AS5ws4Kcr7lp8tHg3o4NzgvsRJ26vsX4QuNejcCvsiMwYR6f+wnWVQKvarmtxiF3
5YQdZM8Q6GYWRDJ9yKKAS+27Q5MYWgV79gnQojOKUJdkh0g9oMKVcRnMVHVMiXWU
fuWYI+IpAknVzdjJathGhe7srMbVQv58GnCQsdpCBOYoauFW3eL7xnaY8cVkM+x4
oqafubWlfT0sQt7yuEa+vFXpSGJT7y0mSfyD0I6F3kHdf6kuN8cdjRhRBkM3q2j9
GIcaCebJwKpyU+RXzawLNJQydOYQ5faj5KlvSg4X1TUXEJutcC6CRwgis4u4u0WO
bynxBMhDOwPqo4x4zrN16dolHXsKNyOBbIYq6CsmM/bDBiwOr70BSZA6MjgSKizm
zknYCPVLLm9AgDexLN+I27y1KYPtDWfgc9vjvUP1U1jsIGdvvbGoPeQTuTiBrOra
D49niDFncjF3ntkLIfwknQhfKr/0z3cxrsPma1/mwH7bdDQc/u3G52ae9p4XjEyL
wn9TmhjQBT3Ng9kPMlLVD6skbhJaXNChmVSzwhH+kvtWvXYU6nJOlp6J9T3D+N6K
cO3dxAWopaFJZWqpph2Ezij6kH8kDigixEus9ApqmSmZKgVyRp5evDGY2smzp3zt
wJp069VaPOI4KhdkuHE8LSr7ug3btS+PSNzbGlVa+ufzLnMpYIUDlV59JQiEGJHU
SmMz2k9Z5jBuKKnfVIHkBjmVKRzpMQj6Ygf+gGwFBCCNxUpcnPzOUcFV/bXU/4gt
4rfH2TwTQ06zRBpj5Sp8G4EBZJzGIRJQaShCwykts+jFWRi2KkAn+G2Zfb74gV2a
yXAFKYgygbGp/46sK0xFLmKfP5StXhue4K28K3qF5YFlE2FeaOg7cnRhXPfNcc8u
UkhZBvod9kwPQvHoUp6mZsO7PkYFFDV5oE8PQ3nf5QaJp7QugJyNbFHy72F/70Xh
0VJDy5G0YtCHoMse/+WWKYr/oTYF8d4RSS259GZy6NIS20MvUsqGaCuS52C1Eaj4
2GJIVEo005Hc+I/5MDPczFExBM9sQa8o7JgEtSgE0WZ2/DHHFntgqCL/maMQlxnq
w3EwnqijJ2i5xNUi/FP3d0E44W7NZpQF9bb55YxOoz1UdKMdj+mNSvnPwQB0Cc85
pzzSMGGQaik+2IFvWCee3qBk3Gp+70s2QoW/sjGjscveljz8Bzk2oyNEl86C6BvC
i+Cpqh/ud02dnzU760KJT43QxHhp2Cv/wCotvkIcloh+KXtDXaWPQDlx2wW/GSHB
JOaISvTb8V4b13CKft6+da/Pyl4+18dLzjN2tmkh0rCVVeh+XmKlXYfmrYj76kN4
UuE0Yp2NMcoVkoZteo2aYEOd7mvBbJ5rfxFtdCBb0og62R13zU8NVDWLEk84LrsA
ZyM1r/9StjUQ8MlDkJhkg4waRtvacBeVVp6Jvw0YPtAtrriQJ7Y55vbD1NMumCon
cH1ie6DeRmy64T8Ll6ss+sV/bt8DvJlsXyfdglFRDUzSK5GdOu8IaKKjm7+g02sn
tQIctsidpw79zdEZFYTML6A6zzDO4DlsJJectc/p0S/UJC+cmNxsjS9WX4vIpYKR
QHBSTjNnOL+allPl30IUczw859uN+RTJVZzPPRpHQcB0X+k21KrWpw8GgcnjlSRO
IjC53PO9VJgi+ggTIwbP2nK83HpJ6qaPkx5pq7aMGLS5xcYrnyBKg4Xg4WYK8ElZ
2RFTNbGjRT8t66EAaiuIvJBAAG/c7+GHK159p59Ql6Rx56goaEbuN1H1qlv3B2mF
jcvxcXTT/7TNF5OJ+EOqO/xrM9CaS7AMvne1afYAd+MUrZ7umgOJhdWhNp+l+X2T
ZvK5YIYRrNjk1Sg7MJMBfEQR/RSEHGt3lzPDofR5Ms2sNyh6fX91Xt2BNhPO7gve
LqJxYweBbz+SxBAY1YgsCeV3qOXa1HIaRYLciI3VXf/3tCAyx2x+7e+6jrwp8FjF
vZnpSb5q3xzLa06FE4ZKPH2M9mvk0L4GRyNDeb/c9xN10mkDjAvHAjXT43ER7TfL
ieKW3Ovtbvy038AYOmkvTS4AmMNFWn8agsvjLrOjMjmVkgI2LYN8yQKYqQvihSDA
WGYHKTz2HKkTwZVSZ8AsE5FEjDOiCrVyIMBf9oc/1red6+RarpDQQbBuSmuajpej
XNLYGgQ2r0W0gWP7qFu9HTo9GyY4utNPOx0fr5+wyfKBfcATq4qAJD7bM9JXMr04
DvDtTHvQJ9eCy0OVNwaNkWpouydDLojHoT0BVnd+MmJKFyP9MumWoxcqzeqon9Rl
IHHgm1wFu6yIu2SNIy9z6KjTZp/1lpdLC7N2dvWe5oPIXlSTb5UhMYdF6XAmiCIk
IHHFL8qwgqUdezV6FJFMacFM/nWVYpd5x3kx0+RxAmoJXJHxE86q02b+eqcJ+Smd
Dt3jCepd/Yithn5KJJ1//Nm5l+FLFivCL8JuXRw50gBKIcrSovK5JKX69Wxa5vGU
w5wvj31cA/l9NJTjNvEakRmKboq3Prxr59LMkYxouW4loWGvi3J+XLIq6ail8n4/
tJB2GJKU7+actAxc3HZWNlFNSrj2dEhFads+N8FOsxdk3cdPs23P0gItpMSAclgs
yt/hAATeYWSoJX98K45jTrlBaD+NWt1g7e8dIVyp7KIqM+HffqEmIp1Fuo+gP4Xu
mRQCR2dO8ax/MquXpS6SJlbVgLiD1qgp3IQtxyB+5+3Ph3pU19JPsOw8VO3Jcf+o
Q1F0c6xyc14YSJQkHuVHJGzQvcq/KB7CLqCWxEzkeX0YM7icYEbFyHqlE/RKzFYT
3Y8+KRa04ypymTD7zhlh/+u7h8xfqHiFq+Dew3dd5inBkv3ufSWqTL9qSOMn5OZE
7fyeth8sCIGDPdErPrpVCJXOje7z/QsObjWTqWtPaYtu5vrdyjrw6WEeDClONy0d
ZZbqUP0Qy9FW3ThUxG85WVvHA6sqXvzIG8q9hJ0q6A2HNUEx3UUwAp1Wt2oQacIE
KcDXtwp0IP2W33iMAm4i3wvapA75tP1dxJ0hF+4AXHlysrvOyd5kRHrIacVBDlsb
MDOSY8tE3qk0phHJmzbKamdur14jS8t5ZAC3aJMfu4iYNHYioZBn6FYSr+zJYkoE
6qIW9hjjo6/VGyn0nzQytXSksW1BA/hv7YkuuRp86DPqzHMeSmOZJ0OMnNMmHUZC
n6qBv2wykdgVGVSMYrovKBTV7VFhvXV9ZThrLmAm2HVskR8mAICYq4hZMxBLdV9H
fPYOGIKm+6jdZ1MnMWeyshfFt7fqAPx8CnDJJ5NHJshDX8U6k3Yw8Coo5sYT1aRf
yehnjmbqk/SqrA5PCLs2temxmxQXcnW+/4777tsqKJQk2bJATH+F9xJ73NW3C3FC
BXLdBD6eoejehZM94xo7M4SjDj89JJl9ukDJYkHtqgTvpvc2zez6H2dUk2KsQb5a
gqqBIyy07aAcvjf+RgimvJTUHqQ7ZxcexYIAQ929B+DMXtsvYklO5DjMqMX9EKGC
KuxX9/gNEy+9nqdVpvVRwUYBSALdFwDui+nAT551L1IrqXNpXUjia9ZtPno9Oz/w
QcK5M6yjOBm0P9uTDDi4wUFi4TNBY6TBJl/eMjIhHFJj1S+Id5Vi1zDngli8+2yY
D93nbVdd8iPLFBy6sZ00h8eRsPEvabbBGKD9IImckmX1Mb2wn3832NKgO4up+WBg
7MNd26o95yFQxuYtHXnRmofyw3DKAZcRIuzWaNsr6x7x/wLVOaXgXznFBEoOig8t
MiMOqatkQulVa2K+8RGpR5r+dDsO9Bk67IiRx5+hGsZd/9x3itibi4lvz7mOn453
ISdOP4WrI3e1C2tULlAQs4zlTbMGPM6/rS89DhWssVpomkqHIg2KkaZ5vQqGr7pB
hTmomKUR9MwO91/WpVanXAlc7JjBGCU7hC+UNKh5pOLM9bsqiAq8wjRIc+CeDEoN
aFw2lW8880F0bW90Omn/ZWcFFPHq3lxj51ewujuGa+d2c0q27UoRDavVAGb/EmiQ
FMNfSiK1QB5ZoGB/M0X3oDtwIzSpJTdOZObtoTBDVsDp1IwEmmY+WXUUUeo4RXeI
5S7HnUJzgRG7Md3o2PkMFgn50rRYuqjaEiR4DT5/08m4LRkmdKVewcSyyTF6hAAc
J59pdcVWSZZMpk4xEeG2eyZyIrBkvSjHpvS+oZ0KgXhOcsl7o4YES3Yf3IKwLrHy
zVxj+KWAZrHPQNV1AgGRscX9aqJIwQnPCSXvViDpy3vi6cdsdVWC9ZLmapWpQReU
UFqEiUvboEpeJm+BQj4Lh1EDyDJHn27TgwDKG2etw9UpOyARAW1m//Qy9kAV+Khc
ASDibgYG2vyCTmmePKdggiZsUP/rOU1kS85geUuFRCxLnYfKerZxwgdFPH8lXaJT
cvZj66XDtHNRpw7es6VhvJaHbsBbTzFBfhVzSv+Eu+qvl0wgPGu3bkMs1OFNLfl5
9Ax2O7rYoJwV91fHJt/74pVLrBwiUCsP88/tkzjHIKZMcGcG7HLRQFhaXwzX9AhI
Fb51fmbp/T2BClzuqQuFWuJnPrf6yH5VKgzvxeA/VvUJF80zH7SHHeMC+iny/di9
sMLLZKDAPmu26W7QvbQjW7ktnizt0PyG8GAWCsQgFy3Y9zp7DZ38gsg4jUKR+Lwu
FRzKynB7SEx7hUbTAya2uhWsd4RjQsw7ddCeXY3Vt4HGDJ82jxOiQNO4hIlT9CFj
r/Kw7EQpLLlYo9hAuE1ow7ujCG1aUuLiSyW/kgZofJ+1dwot9wUmeWMSmjVhvx0t
vD6FZEp8f/GmqAsnBcb+kwUbkn+quqqCOnnnEwUgHQYLi+Y+5uduIqmcfQpCUWjT
Oy9ufI9baZcRPzkswu6rXyYoxs50t4085t/rKTchazRRFkqmXC6/kk0gTf1h2SX9
K1dIo8cIzq9eYknYfHoLPo1IhKrJr41SPbK1xkKr7YUb1eiDKbRotxdqTcbOgCxy
EEWm/+fehGLQgNWpVyIiabpNlygWq5LqjGuqUo1obfkaCDR9v+Dg+f6C6rFTVmyS
hbP6aLw4fxPMpeLNHsuRzEljK+v+eNmuSOrYumIJr/IV9PxwkLiZ2lUK+/nTu+kD
YRMA00TBDVsiPX/LVBd/YfCTDHtiIXKK0vHZ+vCBCidyUCe8l7Ejapfo2ZAcwBpY
D7kR3iDkllPV2UyNNBUL+ONGC6V19JQPBF3bBIiZwZPHMv6nFBxF8NqMlFK0MHGq
K8Q/KGtz42XMcI644MdLNMsvttPmRvfKk7lYOfFXGhy/DU71vcMObwom15U1Vzh/
zeeCnZPrwD1sp1qQat2Gd9G4ZqC/mxZgs+dYi4mPCiX1pug9nfSS6m+vFe1fF59e
yipdd1Ygn7OfmMco0zogAriynk3aoGmqp5jnwyyY9g9ny1AQWOyb7qxR6uUst9vi
swpZN11toV44Ixq6LWyq2VHMu6OIOXfb+tZRiXF2vfE0zUrgCGxYXUfTAObzH+XL
PSyjHPMDIr+EJeam5dfTsTHwv/+s4Z2CgCZZU3kaSjReLswc5CYCeKw94kfICb4c
7x6cPfuX7D2dsULPWFXmYgNwqlphWY0GFIpAgeRj1wiPfacQCwZo2tqwSCrYoh2W
aKtGjvErTxZuJi2v/4FuSxOWQLE/vHRlT3R/Kgu8Apspacj7jI79ezbEEr4Nrclt
VBIHCCQDba+PtTkVyq0c0X7XMAU9tKKisxg5/1eLO84WQO6+qiMgLALqgMDjLABH
uXIovb5eYf1SXuUkX1ATn+jRfma4J7rJmR7h70o94XPdAPuqBdKa6ahqKaJANkGf
T+cAJR27Nd4MPuFojyEn9hMlL9J8gtTAlv5dJP1WsiRWeIjKVq/MedneOXa43l7X
2fOKbwKZnIyZqwr/fJ6BgDxdSxPpuCnO6r/3attHIhdduAZ6ZyHkf4LfvrcNqjGl
V8WBYcOa+RU6rKGKtQCYlYFKFNcOPDYiIrb1xOXEyyh8jtiE7awd4JBRng15/f9C
mTejidtQGRo1D0bFrjh6JBlGg6oA6qmYtfZ3hx6CG8tNTIjshZfspdrzvgbmVFZz
MBXQ6HwYbSvfFYPzdvWoC1RjKpEeVuuftPFXiP1/496UOjYz0VfUqpXJZ5FngXur
qBSiaoEv7Ut8+EfRGrlGECt3WeZbBUOUD4d84J862QsLTL4QJXJnpZjaF9CFMtfo
0lIL2C+gDrIsaoInKjJrKAg35CKCCK/KgvJeCoh483bp35lYKIcMUs8dvwbgsrFl
pqTb5+jPS2GzjWCWzfcueIOtvibnsDIbnT2VyGz6ywZnPJVe38G9VpWHfv8FSUtM
KIJZ64OLbQpyNOlO94YO7KIKNeYtVfOrl7X2OAvg514RkpdfCfpDXGRKQFndDOGV
rshozE2W3SYuaDxU0JFbvuNQP4KQ8laW6Ggt1OWiyDb1KDMbEDD/nPoA9Py8pCH7
4tYCN6S1bExg+dPmOJHM4iLrdO4UpIeMOsPd/P4YAf6cKUUJ7uvzrkMIOaJu7BhM
Jk++ESO0N7V87oxcVtvv9D/C5IXMwDxZ9xmd2en46JzBaVyt+ko/NdVWwzoslIho
dpmAI3w3e79oHtBPgSjP/OpGPuwdRSyOgBUTDYru7fM4xFUD34pZIZ7Mixk0UFg8
eJ1AmHuT/5WbsuQbdHTH7rbI4mZgaiimdJ33EZoGwdILv8OId9qZchgTxCyUwDvA
TxkO3DAh2SXB787LCm1DqSHO+5ScqUirvgUfN2veIq0eYJk/+dwiWJawxqTZ+OjI
j38zMIezsVp7BULWBEclWCYn/IpyzHanBHzwlP0Em6hHHYmRMtcyzO8cojQMxO1/
k1ofhj/D0R5hUYh65bCESBKWejyw5I1/vI2rEOKCeK2T+SZlFAlJR81DqrO+85XN
V9+FxytLI4j9hR2ByVqjQ2xsRMgiBovfaOv+3oFkNcF0h6VOKodB3N3T/TY15VvF
LSvkhnnzqgiJl6MLZbZKpYQrbfKcLTP5kYKVWDMs5NbCQfKTwlvGvUJ1OnTuPLCa
bWveKY4MxcrPePEWugQ0ZS+UAK8v13eHtwSjhEVSWRbnCo6g8574Tza7ua1n2XQT
gMefdlkpoez39Vv0cQtauTZnv48m7VI96paWZotxnHv0Wnsq0o3/nUBbt9tY7c7y
VRZjqK3N8QlBfDv39MrcroAqZAUNxdQ5dWQZxV382W7BRTG4+DIqalGjW78k05Rx
o5DKNyYmf4ylDdFobG119qvw9Bo2f5AaSks0i1OJb4e2PhyUfg0LDr12xzEnKyX5
+46yz8qZ4fejZgYo4BKFXCb/A6gkHWJZCM54/3UKL1yrqXGMIIOMJzSxaeRqCYGQ
hDIkWmxESoG1srvNCphuhR1Ulr+gEkuUgYgMD9w3QW+1ZxoVUK4rhdd1mN3bh6C1
SA3ADRukSXPCNkVIFfdjHlLOF5z6yTAzIbrM414TNtEsw3EV4+ZSa3SHhDeNuNKU
BlFNKMnPdvie6+PzZNRVSOxHrqZUGxIoLLu7a9yJV6hhIYxEnzLM0ncLR8vBLf4r
dgpVeqbYTKJKBYV3f9atC5vEzvgpiZuEFGX/adq0jp+5gkBynOnAXHS4UaVvVjEQ
neUxoqvPBymaNlmpFRCb++957X+5UCWHC7aHjXVRzj7zlXg5NywnxbXieavQXhpg
OesF7KSQooHNrAXtY7KYBsLjebKxqtnoTSFlIcf0v2kV2UP2om4fSfc60uCrM/Ou
76xe4hSE79DSqtUB/KtpXGiHlbYnqbqPWo2kQgxyhnByYBBa61xJF2XMzVzmHcAn
9jQ7Yi8SC6yHh8hZYHZlI84QgQ2/WIKe61VzTJ1oPJunxCWtLsS/wg2Ywjp+/WyA
0d6ne7Bu69M+zg3ATd1dy/2IeCVpaNKOFO3abkjJLhwVzLuPecnUBhXJ0YDTq3yA
P4CC8QEmuEqkkmHD491e9jBMFYtfJF4OndeOxm4MDqaLNFh7n04H7a58zCQ//hD9
eJrvRmREVcMX1GVCEtf69KbWWzT5b5Ox/qV0KbaRFSUPIKr+qdHMxaOnzVzwn13f
GK+RVGwn8YOY+Rj0E1/8d1BBaTAjCrLjDcDdCex4FVzrsZVX/5cR+/Ip4T2PpwVs
eZHSpmgxjF/IUeob7rmgwJ86aeyu/Kcn2hS7jhW9FHR3LJBtn2xM55E3kZSDtOHS
RSxi4RSnhNXTFI3H2w0EeeE51x5fZQTZ+kt/BkEAhTMHdfyctU3hAxZLyhmROuP3
skBphwmmLvr7qk6EZC33JGmhi0gOsAAN8MIRTAQ5YgyOIJp2Y6Xqj2J+QDH3E5u6
/LZKJVSOsaacBlaLoGehiGN3lH9vjFKujkTAlOC74rDzagZxny2XuO4/wkFsKTwV
VdxQ7ApymiI/6H//69tdQ6+ZjwMdJ6ISDyyiCT3ORMkmNgIkMO/k8xNbTyUO0kIG
EglqFhXZubjXsz6QE1S88GytCcdYJOzf9iF6osGQ6XkAisgWkhVIoMnF5IttV+aq
1IEmCaQDM8x6suC2nNwqS1aeEu5C2vuvCvz1CpyYbw9yaI4CFREFFgaXjoAgqN3Q
e7XZCqiGZIDOHBwUwgqxC3z/h/0rMD4H6BGRHcBsfoe3qeE3Z7iBtztmcN0oN2C2
yRMMxo5DbvocGOnS3jmA7J3kl99jQduEWNgkrWuQCfh1BYpLr+VZupx5qs0ZAIN2
qJKltII8aymDkP9juq1BXSXR72dsSCAxLsy7zjlpRkqfWqkDRqpi0DjcWqfmhNfk
mtFmyzkKccojCwYOGNvFZxG49m+k4g6Nfakn0/VrVFsEPx31Z9rkB+3TrN8xaNL1
e8INEG4Mo74cFIM+r2QS7r1daPFUCfgMo7rGffs4OP3y36pxCSi54hKubLUz+Tr4
MwyaXY57YHfErw4KyC+FWQjCjjHlmpUOX9JF431Sqsf1orc6VchkJ0HU/CfoWH8r
8vE6lj8MdWSEokd7nn5XEijiSDfLVbYIFDv2iaj3bUHmj3NQZo2uLp/VTFQYOC8y
hM5Y3Z0m5Py6K1TkP8+X57bUQyfW+qSQSwWcsVGLAuakWZ8MzmQxzMVM5DW4MMdt
d1FD4srvePC10dwR4YG48NlrCxfPYZJOresP2QU888CQJj6uQDxNc3FikXriWSFS
ZO+BRlyJiB+5yamYQNuSQ5U5MURDlCDM3pR00Pb3jT/UzctBeEpyiV07eVvKgo7u
xSRqF9N+H4EAVkO8hdricolXLpqsEfk/VB6LGBHIv/hzbW7B74mlAwOaEdkSzLDJ
QTv3xe80AQB3kiPDtjG9tCvloXGTxbRcco/szdmd7m/nxcAqKM3cC/8yPpnMozS0
EZbnjMrCUiO8zzFAFg1URH/HDrmw23PEeFiZ9JvWRCmTxl/2gZmOLnn+CYN4idIm
3+lcy1kxjYiYdA4uj3RfYDU0EAl7htjGE1oLrAkBwHyc8RiBp1qmoAaVk8jrz2DU
4V8mEB+P49t2evq4bec6MIffX7bpF7ZsW2o1DsClaYbrgu/lOkGOv53fUJ0zzOri
rCNaMqBNKFaJRwsv4a54t3/iGBFz1tfRsxd16WynlhT4AwJJJZ1tDe6cNU7Qc856
UQdMp7EZMrdPRWEgY8xB6GUJrPVk5+uZDUyUuWf8RR+vC/FkmlPBYS0cc8FxSOeG
bHAyJUYD/2G/ZACVt+EDyK9eRycwlCLtUXr7As4dYunGaucmOu4fBPrthwERkUlS
UwMWOFabuO1NgazFuPQzNsYnUO3lKrt7uCyQkAvjBwkxNgcfT58H3438Sc8+DLeh
SF3i8hNJU91mJA2GJQITeYTDAcVAxiaWItjHhxmrAWE1d8s6T/cAIxI39b35r/P8
MpPjDC1AJBelV3qfxhQj97hNgM01EVV8sqJvrmg3gKqjrCq9nQVMkhAKkDeMPG5N
ZMf7EoxSQmRHYLJKF6ZQWvpZFLJCIldhtfQzLPotCeiU83ilFyR7ofuoCOSa4dIJ
d/iZy6j7cGiiLCWWF7T6E6glK5SUZW/8iQIbGdZPYJfXRIvveSha4+QCKmsZ9fen
lnJfdVhbUGPMmrR9tlTKRxX0se5iy+LU/DH2vY5LKmETU8TZePG4+/BgNlsuyaEB
uy0Pec+dU/pdpCVPv2shU3DcBb/r18FD6uMy3e+0WBJxJEfyOuPmVj1pSO+2scid
/LwJ7zYbdAPzJnuBBxUcE8WCgdeAPWEhNR6FafgitjI9a5/PSZpiJAbXUWlXVNEZ
YyuOrQKN1Ch6nuyTXozKO3F/tw0D5OHDhVQ1V7Eh2gwMj/6i3pXZ00IZCb64bHBV
/1h2F1utR8bf+rjbybMKptLtC0o4E2oLumvYKBBdLDV2ar+hU3Ftiu2FUPuXy6ph
4TnDw4ZYVSPi2NL3dxxeP1QHFmRyZ5HyX5gdkyfTAecHV5gyPckOXr+fQpqmCLzv
us81T/Vt4ReWUJNhDy+RrSSnQI2d2xNHFo8IWHusjThM9/mcOQHQ2r3NM5N9DnwA
8H+TwtsCf72xkVY9y4Q14vu+EKtTNTV8/tGDlXNKNatlaJbMXKBMC+w0d+OZqgJr
gCNxLLtQMlJCEMsejPnQ8xUO3hO3YuSibhDLVm/wYXSzUwUsqo0LLx05WzKGewSY
a5JMd6s68ZzhoWl3JCdqFwjQGhQlTf9rZGw2pmngTAOYxnRwUZn3LvsKnOSS1TcV
OPTNhZu7k1AAtBv9xqFHctRHX31V3PHtSjMq0wRnMhAxUPKCNFtN0Ck/FlSgei+q
GtEuVigs5USP7YnEaxAEK3F44gSkuk7WSR4mr1ATlOehCn8WHiqxKMtCtp4oIksr
PuwdZXZFHBuP3KecE5TB6uZXCZCGm5epYJoNMDPsMCpu3/5DIzw/Ox2CN395Ru5c
YRitK6pP/1+wt/TL2POoU1jwrea5z8TYgf+gXLUa5ckRQtzJuWx4YjOUcLBf0Wq7
EINeSVFn9W2Rcx5Cl0TxlNyB6QtxYtfBv7E8Hnqq9co+op0sy6fydUfNXDznOI+j
jIyeeK5zkghPqEh/n+qJ4/lo/6AxbdA7U0fPOKGWyqpeZNdGBb5rNSIp6VFZWnXz
/4+CMZHl9BVoXHRmChtqmmf9RE18KJr2JUDLQ57iknBRlCrjLd4h1xtbDzNgQgLY
iCFH0OdntoEAoWbP4VKQ9wsWAGrhWI1eWjy/HRlQnzgyopIEvbJr6cfICd5GIimZ
c19OIl+XeQ4WQDTbx7znrWPlnQYD0NUZwCNtk1E4jPArtmkRGGHmhJAqHtCX1i5z
pRd5GeODRX0fD2J7zXyBhIR/6lbLzgnooFS5Eer1Ee9jsiR/RmzxvSFCL9lxlzKW
brlWYQmV7z/saqP58AnPHSFYyCrbOZDAO+jw1LECbVVciy4jH/ZSEb3R8fwJNxlA
9RfVEoFVJERRahbEQd2CBI0UbUK5hvKUMVitKyf6WX5/7dGNEPKB9OqpPOHwyQ3k
6ZwhyRYtuTHVevhGrfD6Me/ZKdGQx5RW/7tdI0JjTAThpvaZp2BGmqTapLmy7AJ6
EUTiie/xP6onKXYdv/tjJdAPAKUn2sG+f/+xE3JipZm+lZTajFaaj5L0gQ5PZ4nH
lojmzjRpO7e79aw5SRF/s6hRdRkR9EsINFrbOeL1kAceZG1pjasm5LP3577rPWvB
q74meLFPDABI7v3it49sHAHbYehAnG/c6S+NWRqfl87IjUjsiUqU05aEDOTYkOHa
ChBVtFnniCcr/dA1QzSYVHbsaj56QLxWE5/QyaQMNig9gc5CIcoaU9Qyh9OGIJ6M
I3/Vs8B4EUT1+FW1HJOtpilSJGMOw6KhlqzPY18ChryjSOuysV17gACFMBTsgVgW
brpaCLQsaHKzm+VGsC9EIJgKLZ3yU8xN4fjRvFoG5iH6zoOjbKXeDhnL2JwscCX8
Hg3LfBiMYejJcw6fYDx5Ij1n8Ww6irqw1GT8+KFhylVT+YFnw0Tlpuni1ymWS1Cr
vMpdDBwV76STcbTfhUwFsmp9+ROTalxJ+eqBWsyYrBFOclEqrMb1/w0tkrVi8892
NPnurM14+NS7YX475TMgQevW3dCKh16xxeEgjltHuKslPuVKYtkPzVcfg83qg37M
B3+KwDa48pnQue6sEdLUwmEhY6tNaw05xTEaCoNYREUODx6jM1cvduYiVDhweKKZ
Wpjmf8YMyUUTADejsBd2803FHAafm1SdINjWj+sZoudPAzbXmWqEpELc4qwyRBu8
/vkepbwsiy+ngBAW/HL5LzV/E/7subIFd6HwtvamBedeEj7eEphyz7DdNPNS2wOg
/ki/MC59xxGU4dNVDHJ/ULLRqC1rbCW4civAV2uRXm/VW4hAWQHuWptF8Re9nyrn
/Z0XjgBU9wZftGwCiTm4H51WbknrjDkw1GbkO8GJ69O/EjXlF2zQb8gwP5GdeRiA
J05zdJw3I7xEMHYjx4mC8xSUJC2JCyI7Bkk9ne8RAIbCwVD0oawyrIAQ1O68/UEU
GHQdp2zDtYkT0ElsvQ5U3vPJ3O42ncsE3I7yJezS+8dSFFOrpr+RqAnYLkYi7O39
whMRW7dBhJ4/hL+scB/xiihNzlHL0Vte2DUUjpbEV4PHdqrw9FDEsJDR52NHbyZP
pdaPEuI3IfsA36my7fzU+U+lP0qMFsjTgmFkZvwgaxEw15Z4Gnpnl/1hJtZpYM3p
WcDeumX2FXpjjvUxfmxSBJfUo5Xl03OL5BwKKLzlbBTPQKgypMuKEW2M4zZJ638l
aOuRTJs4NC0l8Q6ygXi/S7czBuuQNhup6WSg6MSYJlNzjF7HCewNX4Y2e7aLbQnk
TsAq1c47oGhEg65Kd3LIdDi+b+x3bjcQukfx89Is10WinSmYQl5HPoPUzJf7ZJ0/
6gdonRnv8x1lhyk/wxM80vhecSjyQxbibSHhTu5ss6dds3iynA07CguxGP30dwOm
X1bPoU2yDteHj2KWjbsFbE8asetlTa80j9d6e5liRtbwpC17o4wkTsiIoIy1bpO7
WOlgCsQC+HbTES1wRR9uncGSFDCdWLP/fda+qPo0th6JIejEGyXE6uu50XzjSgwr
k1Qq/z2gl7M1dW2xya6dsiXom9BBz8BLlw2dVnTlFT9DA5SOMqsMLX1N0/2tWWa9
VCdEKCA2SACgdfzqHYkuFWD9CFKDw6AYN3FKWVcPEc4TjBtaDgPm0o5mX2aUvV1o
+b9/RplPy3TDApuUysNBwl8UmCX9MnGBHiuI2nZ+im0x9ZTxAnOOBix/M99Lmm3C
6UXlsGsTrraJnWJplJCjA2bFns4XwiQRqzkLeSkv4iNBRC+Z8ag2KjoH9c7VjiPm
DBsNJnoAaKppU67s84cDCW4dn/7yBQRhUDMVAFmpetr4oGf+p0Ov5uLGRbhS1E1x
adL5r51DO0oOH+5jeCiX521VfjA69mkChJEI+SlNvWcnAh/w3y52b4r2rSTQUeiR
A7xUM/rLKDTAZJdfw+6s0hgd6e1hgAo8nMUhg8Xl6Jtt89bH6NiK18JNDO/R4a/4
rgmj7tmIeflQJAPxlgsoC4l5X0YdCmmyMTwgCxA5LD6mozpIlNP8NBqbrFC6xdvc
pUJWiKqFBCVksnITqZwpG9WFpxlZlW+hn/u80bcobGED0wa41hmyyFoUC+Kiggxo
2emN46PX9XW2R8h3PRjrj5PBEagRlBdfLOFoFXYyn19eWEkC0GZn/327Ug2yNnPL
IKHXhPn5pvhK9p7TBWJvGNi8CcSAvQOe5eo69BFbfG4=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eCidE2nXJz7FXCssBkrn8ddTjB/2Wb2p+Y7LeeSSsTaMFvdWEb5dDlBMFbIo40gy
/bhd/vbv7YWQ4gUQDMdXB7fkRF40pCnwHYA0BORbaVdgYwUAxVXL7Xd2GE01Cc6b
qkTfG0cLn5//OebJx5+1ipaIcXCOdvG5qsRkm3aFowsU5mALvyQWYemUIUlEV+DY
CW+lEOzzyrasxuxrBn6DLOMdck7epMhqxT9EZhDRPcQ0jylna+UnN1bCqWnsAE1C
VHWJNvv9bTpttrcSUPwPwls14jM3XAQ2nsnZrGCmsbhWWj2qIfllbGhB74Ej5UWA
nzjw/udqjH/4PhTbI4vDW8fTRp1lTQCdVhAo2r8l91lGU/6AdP0q3x+ROuHz4kqa
X9cYGJnT2wcqNyXGFdttaaGSsc3zj2DrlbLcdkJfaNlIkB8YLCuxRmHbeDR9qkKN
XfSEK5X88jSaCqNi3I/cOqIADdfj8vc3L57ByCbJ1dwOtTScKexf/cy780XPSMQi
HZnKlySbVnJ5FAg08761FgE61ZPKk0hShqmt4B2Ub5PH0q7RCR+t3wb8EOj29Kk5
ykcSn5/hmZFLRMXODwrmc1RaEA3uByFwkL3r4Knxs58i6wjT6AmWPrrn/x1iyyOD
Wrz0Qf5W7fJshsDrBsvv9Qd53PHAP871817jSj2NxJsKtURe/W/cFkrXN/ahFV+b
NlVMqV+AIE2lIgoxNaRJa2lhdw6HYIs4NOkT6T311Z1WESDi4j+BtiHwCcS6YGUJ
xQcw1m4VPL/aQx+FzrIbHAE+apBRkqEIULzokln1DB7uQLPINvdkCOckVDrLL1zr
QY4B/1kgm5ZKqYTQPAdjC0XzaqXqb0bc+6mpt6y27/Gty7Kff14oj1Uj/eeqi+cr
LmeamwhUgniORgdSBCLT/tx2//gnigQqCyy8a7GiDyQmBvhUKo31q/gqcIEwZflo
0unYzALTOb+JlriBEI8R/cqbzmxKVkn+HVeS9AlEXctKyicsP+qYfmm6MRrAnaJq
Du0eh0A54NN1qzbjzDbSRA8hxBbhx6ae0X5rrZFuJtnTpdng6VCCBFl1s1/Ju4A3
qsiXWITnLmJrPtLdsZ/CMu34yeGba9//k2Sk1EqC6FgRxsGvWcHyJLl26QNLfKL0
JdsuDDU5GpHcJYu7vKb7vGypaU4BTtvgNerqsHv7YAdG6Mv7ZGVe087hjmzeTLiF
D5V8ejv/Bfur4uCMs6la/f7dVtuz1dzY8uixWGq5oCS9kFQnMJVVxP6VTPPAfkxt
SMs7+5bqmGrFAT6Z90vlLFPAIuMcZPOW65kekV6IHNQQfl05OS+QkWjrziogBtw3
qP7EwsQoJJoXbOnrigDVjbu68LMgElcm/wgd48a1N4Av8hCkpVl45LI3j23rppBc
kxsvMuQDit7Tfa5QpJrn/G+7A9RqB2BjqxcZzEOwa6HpImzHGlNhaQwoM7OAw22d
`protect END_PROTECTED

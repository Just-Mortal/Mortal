`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+aH5lDNvhMBjOTuBTa06v6obcL40f5/DjOg/d+PfzKO3dECHLIvhUltWw2IeR5qu
h1uaKOfxD0Vr5LYWEYt5702m4m2tClfIsRHFBMNskslyekccHO3ypmYJon0ULtfs
c1YocRBN99Vr7kLjQWaPrQD76f5yb1iOHryI1/1FeR/s/FJVnFUk2egKy6X65ph9
4NonNacCXMkub4bcv0LgTC4uuc5BfD51qxKk6s9CpeQ5LXEJFUSG98ekBcopkcMe
pEWVmI3X7mnoq1IoPtiprItHSakpK8jNLBJ53S5EmmvxDHbVtOPYDlvPnGv/yOyj
qGhFEvqWJNQvbQjrStbn3U9dKb/01S1l1/mpWekrfXho62XidQNyjazTr51GO8Ag
dV3YZucHOrzAcSIHnXgk03NOUqBAUd9mP8in1NDQLv+uVqQ9uPPSMQ31VCdaSady
T8aRMysTbjf+KIbxLBItXNZ/0Viot1l6uktcJIWvSTXxTD+M7lpHLMqYG8vhmkVV
tV79ripyVgiZLjCQmqn2qFk7m0Bc7j1gPjKVP3YTMiwG7GpqCLk9Gc5ziBl8iMPn
DxaUiqbAGvwhWGsrflz4BG5OCLNz4vgk0YrTtVTDQDHWOqcfhqeYLslU+DDiEM90
H0ZrQYH/LZEK5Zq66YIzqmxkdotLw057XlR1AokauCW182rHlTKPRqQSUs8YXH6r
ZfomWWk6anfTt3gfWgcutgegy8EKagFAih9EgSwKwEeYV+QX1SmhTo1eSX3dIvsp
1hOLlMtHPln+Jt6DctmAvgBuorzZK1NK/fbMFm3wX1dYN9YXEq8xwp8xCLbk1e2B
nDtaI8O6Dyg7kH4QDrz6mV19x68r8cdy4e9pDQwGnwBuDCNC9YjqZaszEySlHwZj
1GBYWIR+yTYU6WgmP3gWjhKWZu9ISI9aIjyPHHSrfasSU6q9LgWE7ETryFmp5fLv
mk2aUrwB/0Ypdw0VK05wDkipHC0q2O1VPUI1PaP+0wtPMS7oE0yJcWIMfeb6GJCv
IUhXT0fk4sOu9bvSxRzIG8KUlvt26NxrfwxGXxgyC+tj3C7SnZzG7RFidrOt+sRn
l0cS6W/Rvnj6CnNqwwmuL6MbaJhPzPcAgF20ewZYqbmpn8daFXvVwP0vYfpRZx70
o9PPwoba6xQACWYbbtDm67d6mLAwA/dXeuOtriwGMy41rN5LfinKgiso6Oy7mbOw
sDu8Nrm7s07tCzgCTBdolqBHTdbOQBoHiabwkzxMUcSyQlfmoIScjfPZLI9GatjA
dCuMuSgDT2aHATsQS6KdcR9MSxePuYww6nxPYBkLewuTFwHGNNcgmgzoDDnY5f7u
YEwgjMFM7TI7S3M3QCCo1NZAK47bBK7q1sMpzK7kYXUjhy6e4MGt/pyLUUglhz7z
5MLm2mjVCF3vsjUKKoI7RUZ23kKCPT6ziSKZ955Lq9BbPrd5LAf9VA7twVj3rkxm
mnDFuA7yk9jwuxG8bW8ZYGtGBpzo3diHYDys19wuOr1LcHfipv1GHBomgE78LdZT
qtct3eNqSuDPwLM7ZjFrMvYTnfjW25T5vmOosIFtHAtfquEXkKZ8JgqOTw6ivXXj
MnNtWADiosj3ow+VuGmuQ9H0fBeEG7OQ/xZgUgOzcYL+y8D4eXVALZIyM09H4PGE
Z9eEAuW4MlO+RTWD+SFVE1O+2O7Bx7Ggr8wNWh2zIxEyuayPTDqvO/3C3OkZNuuN
dh2kYB8d0xMiwbgmI4SteBM9N5n9b6Nd0d5IsGfBFtyJlBbQpKYZeOpnYg0KSmeE
CYUVVbpbOWwkmvPaAbWZTZ0FLz/Uz7jMweenVP+xqRh6X6MdCNviDtnezGVsd5Zl
VH/1kif69qyBQzKMecikk/ObmsnILSPuAx71v04jg29/zJjiS+qYAK41hqa3dEpd
ECnAxPxkekrwS1qTDopnCADxktK57DlGu6dJrgn2OpDyDijgcBkCwHtyBMd8suxz
ajCGByIKFrnAZ0H3fRj4VvyT9PFCIo4ng9QnAUyys8xQTryTXsxZL27Kig16UDyW
Ai/MlZ6NPUNSymj/eYzE9ME6tp5Z5dhUvpkDd4HR+bgYQKQTCRQw6ISsj1dkr5Mz
lZawrfLYoqeigb7Bbw231SoC8BlsH12Qheo+7pvQXDS5dsye8zfiMOYw0QKyQ5nN
JyL4caZRtfBUb+HIWTCNXW4FUG/fjLzcX3H4WLiWJfOPtJOBvfwj3L5Y/XelG3Hs
Sd2oywAUP4iJ0a9zUwS9uFznAFDQnz/YCktSl4LOxOCEGqkCekIAFQoopB60dsEm
nOiCv5jVMLJDddEkv0wAjuWFLi72N5bYxIBweZkLso4TRih9DdNaip/zulsaUwj3
2ISYmEUyr1OKRf2A14n5MzCsGXlKhMnBSnvUh84J+Uf8I+NScro2AU4RpzXIgU7w
iRDaWrkevaa47P5ASBbs3Yk1RS1s+g5UJv8OsWGmm6ZAMBIjBr0lzoxsL/RXzQqf
S+0XGfaq8QMNn5aWJ9KPWDcnyYaWAtQvxZZQHcbQPu3IStP2gE+Y3MItncXUL+ZZ
6OaK6VjF1JNTQrCy950unfXPVulXhvWPwn5Hquzl/GWo8wGRyLa6o4YS5ERg5Exu
dBWoxP8Lv3WwvTZ8PakS0p7Ls0m5PGnrQ/0pEUuZlXHjGtwhsE4jAi4LbijrPjRZ
bD7GuKx/DMnT3rkJz60U30p8ERMShvJ2xlnDCBBNl9jcoEU41JJOAroJpeJKxinX
VfCKUaL8hkudkfpCX2jMZe6VSPf2FSsKeKPFCzGCcB778bQcwSo3zCQrMw7oI+mg
gffrdVtikklioUlsXa77/stn70gCczHdjXBZby778We/dL0wzrF4C++QqAVLAX/t
Zzl1UxiDc40PZI2eqX5Op298cfWqsJqDmpQ38tGCwFiySuWpVSvlXWmPgoTC5oh2
ujdAlWTM0rUycAcRMYj2Du7rPk6dSZJ+K3GLXK5gkL4pAVhx3U/wRFzmZb65usW6
kCfZRKZOrwok5w96xk1mzuAnPArnB9FEWrSkFNjqrwMwlmHPDYe5RNLY4Jc+4M8S
JUsZyUCpbDojUUyoIumTaNP6qfahamKUp12PgqGIvNInf2lkxv5XYNxnZSdG9iId
qdlBlcjlZKhybONAVV6rLm5DVm0CxZppzgL+WpyQ+/V2h0w6pTJF8CkSfA1GGO+h
BUB0C+8BfEdAW7CVbSiUaNP01N/23T5+MTQKSvnl4M4V5TnofVyzWJNLpMrDrChv
cbrB/ykOXZyywxVXSOiQYE0c0YaNqNG8um/x7/biOLDNYKXM2VJ6dQVosjFPmZX8
KO5WaCR5V3qbiVmuOf3s2IvIO3V+tI8XYBdfI5UQH2RF2+Rgu+JTiFt4UbynfCEB
yg890qAGPjO0AjMbb6LDuHJjkB3tQIl/NoBztcJLZtFq/VMrQiCPIhsUCyFJLIxg
pM1OAHxThM3eBap9KNiURdspRROvAj9FXAYYcQ3R2iuTiXYJkaAYf5RKqX6tJPv8
SNRJDymwyb8EGMtK00OLjNFln5zUdp4dD+VvCfjK00fnQmT3PVBkzhjVehvQBCpp
g6LxrJ0PrZ/zKe3XiFPf7uBj6cdBbVqUvs4ttxeWIZs5HcBAsADYDbvzWpMo7NUA
lO/JA/rO5wDsXJeznKycnWwy9yO1XEyBWstTMep5JiPs+PhlxJkOS2QGAO659cJ9
JGPJyhitkpi2NAj88JhngmaAJXIxHo8MoTUtTaHtjdQg9e2kFDBEcR5JBiB+yRB8
rVNl/od/o3c25a2bxQZzHVTlLkY3Y9EMbQ93hZ0fbpAtY4khEEw1Om6fqWTkL44U
82ISemrsNks7gimVn4g6t4zrjjkLkoafsdSQlMrqr00Msf96SM5xTLxhCzHWa7CB
O3dGxAMzamkU1Q1yCE9xWItrs1+JuMc03Fmzk8/gLaEvJHbmfwtorv0BsJlkDIXn
sfHSUXauhfFs75kJWbu9XZkhXx4zEy1vNF5xCcwLLmnyKZyNyVVic7w1nk1zl5kB
nlhTcWOKlGKfdcyp2BQI1atKZ5iY15y6AmFIhF2szlrfNY54u7ki6m1aATQXHVz7
wv3xixN2gJeME5lpdBZCHGcgTujNVdhOvhZAAk/FTbNzNAMo4Rxum66iJe0ahh8A
JhqnesQ0rE8Xmxynw8B081rBzL4NcO4LSmknU/lWSj+PejZILAUL+OElYIHVDoAh
AnXgzWIaImV3ceHUE9yiSCHdkXWa5oWqYFkJi9T25pOFEuT1vr/bwq7Cdydm49cB
WaGoDid4McTRNSND4UEJoevs5QrUsocw637eIqtw73KP5EKsr7REsFbrbMw7OlbI
bE2YTjkWc7eTeOX+/DlU2ssuQXMzapkkUCb59L2iftBoJ2kRGH7pTnGo3inMcEad
URXJEjmcY1l20ffcTj7YvHoytG13cf/u+vtSlHm1qDfvL2O+kf/OqEt06Borz2jH
SvvRGMOTtV/2QZG6dZuBQo0WzgQWAPKM5HKGF246EFfZ4gcxFDXZCDw+b7TUMh0m
Fj28YwT+HR7DT9OHGuD8E/g+ttsz2EJSswEXm1YvNLNeBxkbOOSif5goyg9qWQi/
ZbF0+EZj361keB5cNCVKMth7igPkI/E/bB4vaV/WcZ9jisd+Mreehz59TBA7H1jt
pMargwjQTZgFQ2tpu4godqmZHUq+iJty29Vp9SraDpWfsxdKgSOceeedFG4rstD+
ZiQxgooos+zpzkkcYG1US4/ekk9uhVax5hNCRUM/esnEc/RiZDN/BCdn9HOZcw03
1c/6gOOz/L7I9kkhOGTlGyR63GeAg+E7tssJce0NGfHsqTCzhrGeH5aJoo1+gez1
D14RZzn15l838gregVc0ttp52NbrVB26u9n9kS58KS+9+3kcxWsdMSlzOWaN2A02
usXl+FrsE5d434A+oPYPJ0zU972LWXEAQpYb+NTb2o4ZqwRQZ525g9iFDqFzuEO4
1go0kMZcBwaSImKV7v2ywY8xNvK9TDfAzHzR5W+qVCjqWvtAU20C6FNqdKSi/1Uz
PY2R4QQwXKN/06YwrMDGr4s4jrR9o4tjbbkFeIE2YRLqiOpU70wnCCaedl9XKAV3
NxKlXpqLA7c1oUxTYc1iUhIKF2EbnIqf4iZ2WleWiFzSzFK3pTgwA05wktbXdWpG
6bZ9noKguPWDR7CAlnOc7PpZjTcXHiOUdmGjlgiuVgF9OyuguZ4FgHYXQFO7Hn9Z
gTZg7XtEyAEwDlDj+Sc3/ft86EhMFblal5+7KcDIX3cTl/HntjkXhizLAtwLgOhu
i65aBXUyBZofDojX+YVfAQfI3TKzyZoe9eNu+Zcp17kyWnyrTYd3AtAhIPSGYjl6
sxIxp6jTkIImkAopimgwzInNxjm0eKWoZ+NAERcdxFujIyqPp5MISk8eyfiYiIQf
cTrhNjJx9vJMk6+kanUdhl/PbOFtKJFIJV9dpQP4K3zLPPByq0k6frY8NN2CnbTy
1bv9MWK8I7trDHZg82Zry/CuCx9vnhzI8xOrDpIVbBewFZ0LqBIRddGDrpLOGYcK
atrdj9ma8BOBzWZIqmy9DoDkqgKQOjCCgxbe0KBmxbR1MQMU5ZOm4pSJopj9L8Pn
l6RmI1+AaGkwaueVbUfXpdzvgU3t+wGS0VLFDIiGZ19yMr8O7itRt3heX0zB08tt
/LxnBd11FPsNrGW+c0u8L3fiiDw94+IYBjhMHNO5NSDL/VRB66iKGl4+Y7K97xAX
yP4rr9CT9zgyw7BMkQWiDlkFOSAqv8/ReJm+z0P8uVApOgZ5r1K17VmcwAPNELwA
M/6I4ZGvOgElYClqYxzxwv4YC5r2fekDDYq7Q0fW0OajhOpWEUkN1zuwK6/T0Uku
rN+DTnhbNHmEag77TPVfu0FNu1APMhhoAa6YSGXNkUVlQpeRczNA5ZN3ubEkIsxz
AJurYxyhAsWxsUvEvNn44hV+d9wU9dEY3jk8RQ/D9XhM6eQiGqkXGqsVos6ncox1
/unx0isjzXtE1dHOVdRDXvnWhWnGSVhi0Q6TP13YGjC5DfCqHQ6jDKnurPpXxXsT
VNx1KPFpzp8kEPEEvAqqkaljbNObBCHomKhSErpq1ldmwoxrZYzvxrhVFKcHYLQq
KlHkd1+KBxALPNT1hbIW/kyLHrUShVf4wnyB4BZJvkc9zIYXzGLQ14Sl1UEYjLIJ
MzaCIQjE62uCwPl6w9Hy3QYxS4IwnpMwezNyfAoQCKuk5qDJL/bymseCXhG/7eho
8ahyXEwKP3DlqNef9FrooWnYQ5Hvitnhoef/EonF2skX3hQXHSXP1GOsizvkjg3Q
jW6cMhqOz/Dky7RTOnQJy+3uEFmaZKhUlRYBk/igjgKNH5+WWUgqq1MtXInFXIJQ
JBpVKnDybMu1nIX6j4xeBIkI8psn3RJIOy0gPzZorjMo1NaTSoIGPJFO/e9LEG8q
u/zU9l8FQe01PuQkGWbF7BA9/HnUGM/5jDFdnrhPJGRlLm3azcdXKfe00Fpm5/N7
UZGV+PgRA8qmwX4fLNCNslJ52fUpUEjpYkWC7yRX0VP5QODOlLPicph5rkGQBBph
J9eya5slBakPmj5pVl7muCeMX2wMZPybjKRpK1mNZ3f0WTO7BsbM0WBw7+KFRWKm
uhBsqXxU/2OYx/kj0h6rkctsTqnosFGULgdDKueGl7X1G0MMQYHCQveXl/P3efII
OuNE9enmxF9wVZm0Gw/7WuwJ4mqpNlrV0gFZAw3q2n+oO9TeR3CyfSjzjdRdIAG8
qjTuj1XuQn7hrOSJDmMtiKO8ZNYHwnvCSIsDRBimXTg0m6q0NgGdLccf0G8TE2Jf
NQ3fs7e2zIMbkzEjcVrhrM/KWWL4edFrSxjYskedX9qIbLmTl+NnnHaotR5ujxvU
YBb/cKKcu+8gbugZfE7AstpQQiskFtmIXJ7Z6sw9iIQW/i17WtH1Bwy94ALIELC7
Iebc2Bxt1CHA5tIs8Yb6lxM0Y16HOhI7AfG9pLi6O8r65iyAXXkmFrBNBLeaKNKs
Cn/JkPjfdbcOxdvo9ivegZuOnmu3g4KcnrAN3dfUw5E3rsoKxbP1GAHsDxM/DnbK
I9mxnBUBzn7EqHcUZVxsF12e0psG8Lby78vCgMdizIBEkIfSvaPsFHadRwKtNIZ7
SpVNo/Vm4tu6ppkpcXouRwGjI2fQC9BbWymSbNdnykuexujVf0qFc8o36p0Updww
di//DpUWW7j9pZDHd2d/iKVnohz2ek5TlMu5vdLD7puqVWNN023i2fdItBKtrl+M
lBgfamhmlSs3ABnBH5vvFFJAyoHzeKV0iuzqZRYxWl3HsF+Y8YvJ1fFblwHNk62H
2RULx6YAsMKFxmNe3NQTlsRqvu2YL/fiJ37knGfvwfG3QU/FJjVGBeeEu+FDlIgF
KBdZAPfgoHV3RpA6SLDVLw+vi9VQyfPVbUt7khnV7wQBGwANigtmejeiOUnyg4dy
SUilRJc6lOk34kHj9wzi2Z/l983xttHsWnybwaGkUanBnxW78jvyX8OjHTUbFULL
gPO+sfdvEUwh/RIJfsHYAy0SWwoY/hKYa4G3VGpLB/LDdBY2Ziex6xf50elZBHc+
Nf0WhbLZzJOAz948cKQZHU4bSmH8u9BcsAFT0rTVTZ60BmiGO2IYM6cOWTgvCQKj
uNaljRhlaVswvACKYZbkoHYS/mT0CmddJOxQ61tX3z+lN/LjzazM9gnae+GLwoR5
rANtvQRg+Han/jRuZR4G69mTeOZ1kffN8Li2Lpr248FdL7/hwpGAEBPWIjV6+0Kc
g5a4dzuHq11PImDT8H4i1XoNgS9ArA+jrX/a7hWo964FMomciLVzdWIgrlPXAYcM
wiYW2M8NcEtx7nMWXmBhFtD1zSqNDwEgJoO7bIXQDheD91NrN6M9mF8o/MUyrXsR
Lija64TBxFS+5V/PMUNZZMI/6kxheCuPRzVzjaeWD0nuYV17P7NkPRsucyCGXXD3
2ELB/9v0q8Xw4RJ048+GusOMEPua+mIju0voFJa/vj1Onw4lI8KQPtZoOsNR8stK
MjdDjLvqFRBu1eJW0J5Run3VaBR9fnh4ty5k/tP4cpeIkxrjteG1vWBbmpvspz7X
MyQQz0Jy4K3xoWF3FZ9S+k+NCRuU8oHB2QjS5wabiOU4PrLioy7IFSDM9gSjjSpy
AXdRwfwLvgstzlWryHu1ZKMVLNuGB5DnPXilPyybHp5qPjbM3OT3EPdQ4aQ1FgZf
3X4YCCAM+mxvK/Uuv7WYF3EXdWaUUi1EyyTY15bbA80fndQDhTcDmgJqB6vsoBHR
xnJVpLS6WOanDBVlf4G7FYSEBmvu387h6vw+jHfiZ0gSv2Iy8O0Nk5n5wNfmuxhO
TjcY+VYWiKDLeCkE1auCOju02rRy2D46E/V6lAVz+u87m6XSUrI1MP6srF+eLrfe
HQHk83mikMlrfYi/ULHhGhpU5+xbULNeHuhd4LC2z4zLXVSAi0gEpavbWcstOT4K
dwIktCarC+Axju1idMA2B20dSSrEzNJdEbb3PmNc4jiH9GhFcYaNTvonVe6Fbexc
C19n7AjGN2jxgkrS1Wi3wlNvSztwU8d9+Ah2MebKbdEO40ZMQOyoaeKTkiLxnrZe
JYgOVfCRxVdSBLOqFxjFk/HvXMn7ARlrU+zophLIKg+VANGuUe/gcZXvWq6EyuBD
ohQZJIBGQoiiYC8lKIHhOeq/mTmQwhlQvqQJEcYm1rtbqevr8ABjr09rVuclgz0i
Rj3v3adV8f+KGCNGQ6QIrVnkGq3FMLSbst0OWq4OpR4v+nzR1FG7oWWcZnJl62V3
qnX2fwwSplANlrQ795xRKCiia4Iq7WdL908UqxyKo1Uth0lFDiLEX1gyaBiZ1nfR
EcwRGNjprBgOZ7FRVlphH8CbFCYppkfNYBAjWhawEH4+VEt2ENzB3kqdR9zlVmQ2
DOju5gIA6zuVpA5l9deR6vvGT8msiksRAIrPJpIbOQz10eif6ADmu8vqlJp75b7d
5pcTlcB3+qyAQld2Bu9qi+zs8QYEpyOCPmLTeZRWa2RokaQLCPXgBDENFMEBhnZg
MBapLRiMGOmxQmIeCwtLY8bPNrhkXlXuceBmf2X/C0V+MeaFJznoRiJpNma2pPzF
K9gw+GOYGKmEqKbn9FYzN7Xn+Nst0r7YiqvOo/kuFefGnJS+z2q6upy5SkXIiYOC
ME9g/SjVEp9NhH8M0xFEw/ayHMS0HUGi5inDYklNwUxu+6EY/xThnqBltQptOkvZ
ddn4SZzK7yexGtvY5A4BwDI6fCZ7qbHanGoTGF7ZEFwwr4PevPBs0v7hbRCiSFSz
f1/JfocjiugIXHFkDE4MSKfl8ILu33KmGLA4hXb69n7kutYDx+Uu4GsqYvYESqLE
7u/7z+wHFRqf7L5aGdOWqtzX0uAUc+Z0tPfcU2kJQAfnr4krN25Qn4z5JtvLzGxh
YvNI0HUGPe7aHbpGcgcnCdUGu+l8LIyQzyUqSakjKxmIvjxHF9iFKDYu902YofgD
QWhl+4B/nDh9NfT6dPUPZkWeptNPK8aHH7ELuvhO683+J8WOgbefBk8BBe41HT71
HxFFlZBbEDcf69EX8SK4uAS3d1C8yL8InN8v/xSP88KvZDwAbLGOT7OwQjjjQ9ZU
Y0Q4VzxALfM+6pC5k2a17+KViKGVJP79exKrtAA5GSJXvUu1GWuonDzX9AANadEc
CFNEEHfnNi+egIqE33pApZPbUKJmDfKMsUxeqRkvzXJnwLxcBNcSkv4IirzPkKyj
LmjdEwjKaQlSm9FSxekf0FdY1A9zhq29k/unALNEe1EhLzBHhhrxF3hBFh9WZsXc
3MaMIa8qX6sXAl6Ao7kbDHr0Vz2IQTgRHCM1nq5ykHPQDPVKM1wAkwST3shkcrso
KtDsLjswXsd7gELjsMN8uElGI18niobZcgkBtlcv0kU3D18WwMTM76cDeUreRGJ0
6CwTskd/jrQrDgsRj877inBWwO1TtwC/HCbQfm3OgOT8j4BGGWhL/RkjumTFcw0J
0/eahZUynEuyofhwYqM9V26qSdjwaIsMxpeWpFX6F8w7c/14MbbGU088PsP4V8hK
Ud9U9StihSdqV6wUyhAI6cqf8sKFMcOeOPz5zmDDWEd9rludjSy+zfwyxJJELPx0
inFmYeQdZSdxn9VAJYVPZSHgieruYXD+ZgLpTfEnUgbw8/z1woievcjFiU0631UF
MppU+vsKRJvJMpAkXoIVbsDo+tRoiJyvr9pGDB4rZLHpqHaUO5jk58P5/wIDB1Tw
U0crQdzK5sbHbxpTiSwtnjzDu/SybTLYv7Y1BKUy9YjgEnRxLK+A8Dcb9bZoBkLY
+ysKr7vVUKVrqNOBbjalHCheDJFuTG5eEagCMassQTPLZvBcViYcpLLhnKYU1ca6
v4aH3mZJiSUpqRF52Qev8N/m2wb5aX7W6tKBKQRPELALGBH1gHvhVafGxNOpLd/3
K6iaQ+pWeyk4z8vsTL6bI0IDmw8rt/Qi8AoTBoGOa5d1hwrg6lrC7J+Nn5f8L2uJ
6I/0haM5u7HwbQn8yxBwb5tLnP8f3RGfep6XvpZVTSI6h5BtbH8DQtxG2LdCcrt8
6k1me/cJzaEGTGx16Zqxpu/ag58pWNrEv2x5Cgt4KfEX8FywTDEqZJGsqMFeKteK
tPHUfQ2EcV2Maotjtg5o3tv+sHjEu+q8LlQbnltf0kV2ypjMxqRxc2/D3QP8p6n2
Bu1QuSmasA31ewCEEStRzuglxRwFA0Co+cdn8xyaRq6GQtn8IA8WtLBXppOQPEwo
wQtB6n4zwFS6Zc/0R53qI0kmwEJ/aGAoRkHfXaFD7VeyBvLUY4mkM2c8RmtFH8AZ
zONL8jM3nsedOiB227HN4JLvVYYIsONQ0noniS9d4MXN1Dg3wBPiyKzcjllxN8sF
rafiDUJTQBySQ3xN+YVNKs1D2QT7drcvxmHWGsa888FW68Zxqg6ttDQQNpQpRNH6
bwjQI9KBTqAbX/fzk5VV9NBFeo2B0smdWlT6fVUqHzjAHJ7LzTR+sCjriwukXF49
9BN7KlGhMlxDnojnt9fVwii9MtZxfJYZya3jG/znwFCuSrp11ftFr8slIwi0AoMW
enHdyBgjH96vilMLH6y7DeERwnvPzp9hrT68vS2V0NXH2JIXLAOuhJ5yzMR2V/Iq
1l8qaJJHBmRoqJxAsyROlxF363sJn91IBV4cJFGakEnRAzPdQ4buqcR1dhtm3jt6
7cd8yUAcYwsKLwMM4xHtimBIEI9FArS9thg31JQL97QPWehqp5LBoXsKTDvKpkmG
RUjxgfg4qmifB//RhBQUQVzF26DbRR1Yj5ZBLtZKGf7kjpc5f84L1AAVI3dJx/fp
w4FOZVLXL7Citnvw/wsZ1Ldp21fw30AkMJo36ACnEO7+M9hOf15r0dZWL2MuWs3W
qEyYydpGhtWdAdXpJqv1QCh/rdyAAkE5/doSlrpI71cY8WITKMr1Oad9FLq02Z23
mgLFQq8PcRFvu4DTANgXjSIWkwB3t7M6DWZ26NhJZHIPaMFlwC1kEVnp7KnMQ23T
008Ad191P/JRR9ABh+t37uplI/9O74YMFNnIERV8kVvDSWArhmciEhizJEnHLcQK
RKkgUrLWp/DUKz3ePTEZuUZEBJ59ex7Wb2ZwfaRCofvyYyNDAZIdWg2+rroEuoxH
aYyNlWRXBMdz2Sfago6o2bNLIpfl+Fb1YxPBqrRvGIHXJ/EXuxcN2g7cSGa7oGXB
MsiOK/EGix/Ngf53Bdu3ASoL7L+u2B7Lu7qty02hy1Sz4fMBodzsYYOrdMulDUIE
dvP5oe6JWlMSxeDJDOGo/ye9JdNYaRY/honaszQMHV6n1AqpcIbh9phyZ20p/RFa
ctcAmdQfL0jfTzH0m036EvdGkmZKGBSl+B9gTgcKv/Hg/jK6VwWilbUz+speA93c
xj68yTiVjwvOnBX7ueMsK77H/3A2FqzkyGJEjmKZ8B7yTSnQl0pwHIByWJwKiNSe
tebjMHwb6qdIT/3Qk2ESQjAGTOibbDCalKG3LRDPGhbghg3N2B2pYJr0F8rZo1oh
ZIbLT0M7LrmxkBtjivPoX5VNUU2ATeubAUOh1wJl7wd+ofhz3lq/PqWFfNJP8D1P
eL72mn1p5ABgTret8OVpj/32Rt9seWgbvBqARIUC2qLxSEXL/jU24QYLY8QCgLjd
qD+md41xyVpQfSwbz6Z6ymbfWmyKD98OwThddeCJVl72RyBvJBf7tM2anVhVppfR
HpyyXiuax1OwkhS4nHBUPZGPzjgBrRBE/ThMR62cfR8iS5flUyydaL76BNfSjumz
z8ho/Hc7C5aDSWQBOP4infmWJVsAcDp2ZNTG4QRErTz4qGeMuWy/T2NvJfeNHcqJ
0zNDfgW+9q+eZxb3EYDbB1mCR2yFleNkG0l/4Pmof42s0l/j2lVfRiHBhkWnE2Y/
ms6u7plt5/chOC7Cir59VYcsdICRo46xXFJ3uLbMp3XzZsLt+yoE+A1AK3NHJg8U
YHF9wzIRvJ3qlGVqM3AJKWLw4M6U4pP5K7223e8QW5E/bho2SLNjyXW436JgZ9u+
Bq6gHxeAmoHUya3CZ07B7XDU2zu6NkHBS1MVnfNsXJO+5i2KEFv+JeQ/YkHOryFt
v/J6fMn/Zs4+Y8+PD+tsheh/NNC7oC6LwyivJSVKHxP6Mk1TA8TQFFF7ImO8ZcZD
8+7iWSqNiug+nbyS08GTyuP7StVUGmBt/HU9yhQ/NxynUBuYslS/tIFGNtGYmNBp
AxBdeldV6RUrA5CLgCfvd6BOq6gHJCFcfVp7loNUtluAUz9GGRC/PTySktZBs6G5
GlFNL79bhkuaMacs4TZQuMJUzW+o4K1VxVeY9hpSGuXoiysNl8aN7fbZpzF1Qrd5
JhTCYcmb5DcH0zwW5Te98vW4p33RgGInxI3i4fta6ZJBuMN6gnMmdKYFQnp3UDnZ
LUd6qakrOlXbpw159+JJUpfcIwuIuXkPUVQjcSubj6qh+7vicw6gt0rsTfIAhku+
0Idp6+/tuhsgbjC2uGcb3tQqElchv6cSNOu1j5tjo/TLb/84+dANV4QEuNwy2W8n
xqbJclBKDRQ6zuAm3YnWqVlR+MP9bJdcPXOOBP1H+kJIAp5pZYUgbyTntuuYoDJX
0mQX3fpEzpGPO7hY5IHjS0FkJqjyHk5oTMxrmoEi6CfbLMVXfjyBGQyccLEdTVOW
rOLFjajjc4iBIGd8wiiD4q8pe44XlHiGsfnBWF9PbX5Cc25qu1sl2XKDGNXFMx9j
1W01nMJCkmeM/1dDNUXMqARt6CKmXxze/IgJHFjRAIquWjaTYxux7dUCvaQJT08q
X3VtsIhdbs4jGMgOOI/S8NTtUxn7z5WJhjdmv26rGnsc3jVAkOzi86FUHxMPCcRu
M7vyjHpAj8VLQbNjbdr/lB9z4oUO0fy7mKk2fRhymygYrlr8e4gC0CjhDzYtdtya
wOSiVuc+HF7BO9MLiRQGxmrIU8agSlYBxKdiNNtCpU4oq34RyEwIZN45d083uptI
4FsGtQ201hXWwOQyVK3h1U9chWmcfP1TjbXQu5gVh0MDire81aGmmz+TIFmu3E+o
PohSFNiutMjOFjJhNYFD0RtHg2UxA1bMHzuTCcTdmSHGy1mbWDZC1q8eHpbOWM48
KaTPun2xoiUWvGxr0ARhTh55FVAXZC8gEi+yUbDZnpz97nf0SfS/dHc7/wv5Zl06
OmlNh7uWxzWWXXXLnIi99VTQ9Rd4rk8vg/UZBNmUG29SLofuNiO4Wq1eXlm2lbQW
6/DblrCaUO8uH5JaFqdim63sU9up742WCiunsHB34Qp+EL8Qpt7OY0JuXMbCwpJD
97IV0G5cNqOcoIBUsXsDanI+CSics7Jd9NlOckezXmAIz0Vt84Lv6RdgyUUpV3dX
U4fcx+qKJ4PWO3LSspYx0Up5m6H9aT1kStAsPlSgz8lW6ps7BRGElinHOokxxLdh
Hh9wg1axuThYY63+nNLbW/WhGOLKMBsb9Ds+SZu2AEGblTjWRGTQgRwPiJmLHcbq
YWeDDEdzWH1iyRqwprGacQYs53+M8/VCwiQ1XyN5eHty4b23boGMudyPmkDzmnhn
9qH2cveZB+A0jk7CXDTWQ621nNjg3Id90sg3bge5iiTAAgcghb7SG/tgd9qabj9f
VDjqVyylrfEn2hCVCzVxo+lPjQQ9jGrSyC101h5z5ptuy9BMcgn01dApTE8giX0F
P/HgiWdYfYtv7q6OgY0+wbYpMmTIvDzKzx7voAaXK7CACDi9cG1AXJQVlThjUCqC
v2N7TochkYuTWA1uGfBDggJcbggHXffOfpkiCjf0HHvgFHjSVLuQnMLNF1RzuOCu
CZHC9ZGozzBSvy55z4/5haJpJYFvPjvTj/GNrKXsEOe7urFzmDbn1tKtA6f6JEcg
1hEDINotRRjGQFuurlMc6ZYPpOFHzutKT8tudCgkdb7mGlC5R0eYBqWulWvr44vu
18KMzVeDoQcmpPb65Lok/HFCtbpO1t4dgjq1QnQd6IZyo3eLOX/0lBVzthILQjrq
Dix5e0tVjo/CVH0L8S+99nhDf0w8d7EGRoRjWJnRHONHjr9Ds7NTZUIMAW5TpMSg
0n9UhIYHjN23BS8IwBxxVTph/phZFfNg4w4ZnbJU6+KWzam44NegEPah2uW/hm/T
pk0pLgGDr1Uk1jPTULSrULV13EZa1JHtHGEbCzn3lWgApBNN+3BNJGvQOZTQgDbF
E2ulqL8opaXrUpnrvzKvrYOBTUUiRQGPhDcD4zImdzPR4S/xC6dlvnpS8dqE6fqu
HmTmQGZE4yB1EnTclcWkwx2TquUTX76BUDPk04yziGwPQunRMLwd0IFAo3quQB0k
GdtdcGReDFhp9ghscsuf62ss/ZFCO1DtQDUBy711EhiF9fRsziUN9Qg45FK7gSYs
tPMWhtCD61EcQM1T9sxwjTqQmEBTUoZGRVb7xTJG6LbvS14p6tPfPM8Bfsw2x2RG
y8X6ioKkF+Hi0UI8OrVrEog5q7Du4k5IsOcQVmRFWSV0fG5gGuxcnuwPeQ0sW58L
b1VFdYVdU0qayT64z09CrTu+WigXJmCVtgsULSwJpG83tP7zSbPEtN7BA2PaRH6o
cGyzcsM26K0qEJG1mUZuKKke03RqxgxAFv7uqVkdQI4CTbb7oYwwjEIrk5HJsq3q
6GNxUiljLBOOLChB4XBI6stXM5aDZuPdIL2sTDG6ZiNVcsT/++bQS96tydkpXi41
diqxL27s7G4Zz2lZa7Z0YrIQi2Xnw3+G+JIISl0njXYFX4Jm9WnQVAcJfoDQubWq
Uesti3TWVW2Ax6SqQoPi1bduWY3Z3bWBgrfYYkBCHszxnSDDCKN7iqVrioF7sa4A
5Yr2uMgTfohHnl1GdfNCZSXNtSuVBfERfHoe/fHLXwQUpU0FNGF/3NXjulvFLMfY
SLRcvxN98d6J68Ods62ImK+CzAHsW3uTHwKAaHE5m/tLY20R9zbhCYCyWjc5X/t7
E3VWV9Epz4Euzutke9YTrXTjF+t7YozXCX4RSlkjFeJ2G0F32dPtM61iZmROSGIk
Co7QjeKBEThZpN+Ab8oFqePpg3XfgtTXm8F2lAHj0VQGLwonkhYNy9WO8XLHlqFB
mTM3K1l/oEJ97TAIY2Njd2TDELesqdRUGKWpFkalq+LJFxsQPiZ2T3TBrbMwUpQW
oQj67bNs3kfMPp52HUAGCgnQ9Yqe5hSpYp9ObFCDBrQ3f3dbyBxhQPUKokqf8gwz
l1PIgM3PnM9Pt4NrJlVZ2d9WoU4p/Cyp7+9bk2raU78/kzzkbiSU232sHNZmZlWI
uH26PDf1al8FrJafhiOFroQW/dPdg1PR2leOqhC874doqpRXd8L7r3GbB9Fyw2iH
xV5JcfRxwJs3fyp+5kml14zogZJgt0eYcN4D2pxC1FJpVWJVjVW15EYwGacUcadY
PFEutbrwNTiog0e8NSmkk8hH9VxGD6ZyaKQRAiFCNoTcwqQsdq+U4ortQxq3mao9
IKsvXUNv2JJ+91SKg5o0+d7Kc13wWXzboeXqwRuzO8Y2ZPRNlso9M0gmR0gmFtMz
TqGPhIS+eRYzyu+wtHnAjze5lFOqBsP7fBxW/Zt2P2MZi4472fv3jqEC3P1Sdw+7
GwrlLIDTnsCTEym9y3q5gFKocgOF5cKeHPZId0j0em+nYtLXe8TaygsJRmN0a6Y5
YUY0GyB2RQDRx2SJ7xYkvZpqhzbIAfWcdxhvXYGYtdYlsNYnejeAnoDB1VoR9lIk
GX6qeTueciteSLJLqwUPY5oUTFnr5yFu5pYGJzXMm90+XykecOOFQhtFupm2SnzI
eFIHWOkPWRlVTWbRce9E35YgYqqwvXSLjwA6r0/e6VO3FlfO8emVYqaBEDK9WESj
yyoxiEZrQuLdG73qbGVIu5A+fpupfW+nWjAKyAsswrnMVvvC82OgSfxZ0OmJfvB7
SovANvomnPUlHc0AHsGD9Xa2IDc7rJ7NasQppoGMmbc6Mi87aQ0qX7wXyVGs64w8
rgYMPnglDiP0F5slrB8CGAcvCoCrw08zURTEqa5V+XXbm6sWGO8+R9vmqoSWzhd0
oLEYrqkrUvD+rZtHYwvmUK8ueXlWOG22hIyAdGfx48R0ysolvYwNN+73bPpH0dH7
5fFtuvG/uG4yuX6n5Q/EPp2cep1u2So1P03xoySNjP0u0AW4BOttbTIYJa5f8WIn
0TwfIR6W6HUGxQxoXH3gqMbvVV71UXfzORSdugjWNwWAgkdVDbhEJscRwFgHAMIr
OenWMMYHMkZxpKh9qrNl4gl26rGUBQXvQHwqPHfqmIX9BtjvhMO/swLN/iwMHMsP
kCNql1YWLorxT4Q+xSLHGcu9hWbGcR+3p2IKWtzoKqPF0h9CAnSnOKmRez5vEUb0
gjppnp+3cagt52zCjQ1w78Km3oOCh++VzpNkZv44jDvbJhVK+fo53Qs5ZtkhrK9p
5cb2avi0HenHYpUh0qsyCvCQetCTD0reoa6fUsMXvT1J6niXRCxX9xXQpld9+vKu
pvvPgmWx+l1AxMtDga347iI2lBNeZ5zVTxlgcdSSt3Y52SDGQTb8NqWcGPK+7P2z
lDPTef0B4yq9HgXSrlJSLNajrLs0VX2t9fOSz0GLX9XFlN6falH4OEAon4eDXbH6
4Kh5DdzHDpNnC1OXwXm/EafIi69DOTfiSJgZB/uwkudpSw1GdWxJw9LyosDrdMWS
8H4HyxZBSC4gWM77ZgoHTDgLhJbbAnN74W7pMrhgXIF2hB1C9f5U8MNsPIt2HLhN
hmmR/OYiUgjQ1mWaBPh+Z9ZqaOj2vtm8rBlIB+Q8jwkiGxNJlMDjQ0ixk+8f9VhS
i1VtALtSzkE0ImeGCQ/aLF0Jl9Q2GX6sRiI/h0QEDaXwPMm6YB+o7BoZ0Eiz4WVk
QBBL9GUAO8F9ztShEPPmawnufim9SZRGKUfOd7h1ZDGzwq9PTBe9gKOTdDHjy7e0
W0NAX2mhyp7fxtjam1ipqcK254o1Za6+mz36hjm74bwcRD9CK58bbUsJ0ygVYRSP
k/ZCMDMU1SLaJwvP4U/fWThZ7naU8EyakZhecsGISj2R1URHiyRZbejjOgdh63zq
RDIyoprPMstwJTEGJI9MG5fwov/ZozP+oh+lP5FdkY7bIGWNOj38nPVXPv3/VGEx
ftsmQ7drziKz59+ZZyxkj7Cc/cv4043x96FN3quvFAB8b9bv2RwVkUkoMuqK8y/U
i19SkDpAdIQUqwA6mho5SNfuw7BeEdj2XzCzuasp1MainkCWdI+/rkSmrbzSOdF/
cdVJ0FqSxtQK1dAOwDNLve5c83uUJ1CWis574Wa86sg64SdMk/hdzqd0O8BBRLBM
82xFyE/JRk3vdi7sG5o8A8j3fkgVTWCJQVpH+P7X8xQ2P7QmNIuvgMm2CSEwlzRL
NuGIUIW0vkJlsWXDLCCMiCBtPuBoQ4NOAWwodw6vHnseVOPf4Z7bGWpwOgNg+aSP
lVIY8TxEkdk8VJ7TAXBBBr2mzXczZtqNt448XbKcooJ0axHTxGiGn0yL1RprfYg0
mgGeowlqKE6YeNEM5dWpSYSlQIz05eHcY3fq1TkoNnhgC665a8S38wUYepvMIlbu
H9WxQ7N8Gd5C6Pz8WUGSW/3NuFyVr3Rhzfn31WtnQLZJK43yTYJsLUYsR+FgeDkL
IxepDCBsI1JiFFgtwbXBEXfZ7DxQ5bdftyJam5C0Ae/T2mAPFB8ZuoVvJsvMUyQL
MnP6Y8/sBec1vny9JMPiGtupy65pIQBZeaK50sFeo13s0aKuFlgVE7dfXsdL//v6
adYMOyWCnoAOiqhMpNTQmhG8xMXzcM9O7PSMi+Mymh7I4mSTMVNtiGL6AGa/DO2u
j1S1Rr3vlqCrb7PAhryjQdgteXK+WxxgQ1RUf7OzHCTk9ppjr4B9B8MNCVKt3ENw
hmif9ingDRD5A0EeeBNOEClPS9wWidhyButNnTjunL2M5dTBai3RI8Ng0yDW0OI4
obJQOzgHaJuDeWbM1DiV7xmouXuEHizPxZxcwImJLRZ4R14M3WLQE+iosnLjukC9
aHrlxRucfHkYu26y3U7Ul9x8ZYz82/Vb2zRc1fWSHzKFGeWRKwKGC5pFOn5wo1Ju
7JCMxIS7vNtNSy+IWJnAqQ9AZcg8KnInPHHPnuMdaIs8bE3Mkelb78n2HSxbF7lv
87uWqWnbBtgLcRUTVMeutcHG8IakN+Mf9INWOIhKEOhaFxCXSO8RyF335KhZzC1p
5duh+yLmSo5yEh84iTxrid2SK3Z2rHnJAoltVjixG0OLT2TqLuhiwxdiuDq8YLr7
EI+qDLrZcbmgGUfPMAe/k4Ll8RZbs3D3VbtFHzhlXbQAtLgmy4fkHF7Qef38eohS
kVRwvEe55RDqZmEDWU32IE8zG+spWFPpn6jJDiofERw0yEVd2tm+90XxFQibE+FH
ADMSpk8RSC+d9vL/cZNbUV3NKyDh3kQKKwYL4OhDu+SNbS/zI442wsqB3xGVNI1q
8ZhKC8WaLDrzlEj42E+r6PWxOsg+ZrNr5P5CLo3NwX66BIMIShyKgyeEjKb/cJeJ
6GbNQ8vNfvlrlnMzpt22X8NYXVCHSBkrJ+s4FZJsS/BevSjd5lImFTD51GsZlr5x
Kyah7fkCPVCnBFGzAjAxwwt2/+Gzv4fl57hIe38opfTNCK7ajhdbjozJGpbm9lHn
rQ5imb7DaYj0hnl/FZvZgHsjnLMybE2eGzcBxTrzEUheY7QWEspKztBls6k3f/HR
dZVRJ9VdyFspWkTFSozZkXSjvuynVGgrc4YspmNnYW1gVG1NKtMy5p1FYgZp2tJf
uo9plyVJGong5s/bkeF2nCHGHI9jKVRL8c05oVXVppvFHwuQkcPzbDlOL+A6tNn/
9IOD4g0YPDY2SFKewHM4qCwS2xSzBh7h1mpje/69VtsyhZX601USlwsO+aHtoH07
c6Q6fSJkqYjX9RqvGgBVL6IsQ12nj/80qEb9bNptjUHWBubmdoEaxRmIdOi8SyQH
FJE2YbYAUhOOKFQyF7EmlTYX0AV/vqcItMV07rsE0b856JR+vzXrGSEkUBZWDTxv
DxPedSMMGvRfaKaXUj6mTevpChOjS8HpD1MK/KmzAPIglrc7KJAwJQpGmVoBv93L
oMVAnvdcGTE2GpL2+WHVW8lG6IVEmbSiA0yoTluTinIMAaAmgmd58J3Dev5UMxbu
C0XZ2iE9K4hyTrROZn0neiFM8XucRUqONAYQCIOrlWQe1wxxApIFqGqRfg312XzV
JjmcKKTKn+bKLbjNqmuzK0WkZKevzkgVcrAEhugt2ef+g8mi2J62KvHszKzGXzoD
OpvvquVmHx2gf/xIsnmoa4tfHTOuTq8fo+sC0BVfMt3i7OHME+A+BPYUH+5saYpA
hvXaEvlHVk5g+T2HNeap8sPljIVQu3MDarClfmXatZe+EVgHbNjOVLQ7y4HnrdXm
uH0nt/uoD9Z7PXFhrjTO3CxZjQ49wMblpkPZNuyEKacRWBX2T0kbazuyQgszLHxF
20WsqS0+8ecf9qDQGQ5SjjcSOCfRYsbE3Dzj3HV3fkTzqv4JhoGZdN17iSd0Gax0
GPns5pSzDkM4TobkXzAh/Dpdl8jlrVrCETpebsdoLvPkL1P5psZcAlYhiQw1hzOC
LPplgpB3qvgLvTAObzxjgjxUpa1ZV8Up02wQC8HPOja6iyEmNRZfeuWk8YcUmPHa
kz9kj9fRD6wEOumGYxxKvm7RHT1dtDGNiMLMXEYCWs9MFfIYUVZfuHMjlIE5o7dh
Y5J63CufpkfGsq/dBLZSTi/kvMhqaZxYwkbZkEE4UiNsUsuxT4x8LFjy6jd+itkN
oznbkWbnM+fNHl3KT4zjoOyS5Oqk0Ml5o1P0/VEh0bFr0IpfgtE6wPZKsGzMgFMg
4691HNI036WTc9bh2C4YzrPR4CmMN2vByWrn0FyaZCrs9AXJGdNEbgjSoJ7lLnEr
Uu+dMev7ukw30CCdaoo67QLUPs+EP8UpM6qfqwXik/n4TChyPijqPd5oOJtbFnw+
NzPXM60XOTiBRgeDRetTQ7DZnaos0K5cdHeAKSYwJnI4S9H5ftHroJn5ZiXsOZTK
awqynDLW6Su2h3nYWmVsR9xp8j4wx/7yKW6my9U4CeUk6KmZ9/R1YBiuyXA2r/SX
4equTNMEcdhU1/gcBbs94tfSUYmk5v/JaevDYo7E0w3MUUF+WT8WM1R7Fx6Snasb
Cp8wL/gfB5LCm/kmnKbE7g0DWoPA8kQo1nuhcST5/eEa6bL1m9l75PwY7paeKUSY
k29VZvXKcDDjxgIQxsHaz6e9L/ZlAXSYyffQCYgdm18LVfLI1l1WfVRF7MRS1u+y
awPJAn6W5BCoWShxAdtklneNuND7ZwopzCw5PWxiK293C1/ZNe5zvf+T2WnQ5jn8
QNoldgptaSUleJcrqK/7DVNDJ2qOix0/W30hYbkdew81u2+lQV3n1fyw4y17q5M8
8tO/+C8I1b6h6thVhRAtQ7Go0bAZUuS0pQYdfOp17skdJ47gLldpNsVddrFBZyKw
Nl1I0C53cYDugg3L7OB58xnMJR45rRXKSe4/kc1XqXjjQqxpiYL0mH4FdKGpo+Bw
vA8onhY9ozq/ENn9iughy2WqctqVculf67t/o/XYI27yCWsfusmcJRLlsNg0yaA/
cdK/C1GSV+x9s8Wj/mCwdLhui6Ou9NXtHvoyt5mOUiSsiumZZAyuUBWW1VZGX5Ym
NMPFVbI36vM+k5ffliRVWF0Gjqx+ZNSh7KAWIccyxMTRKfAhaJ8tgS0Ra4V5YfPd
P5Agn7dtSGer8C3QPshr22g0CqOfhwlkSYvYy8zysnM+eJFwrY2l0nG2c65kQ5cQ
vp7DSS2NC6cWeIIuKBnWTSrRXRGSX8bsfb7z9OkyDnZBeDS5B1vV873cJoFATCta
KETki0Y2+Y9gYeiNij+aoPefMnsbWxaPp3Q/udXb7Y6vOn4omW9LPiazgAAD/pZp
tXf5JfvogDqOjeSncvz7Z190Y5TB1X08lzXgU3wlDJhnb2ng6gpVGV8u6oE/+CZL
kjuX2dVVyFd6k70EXUGp83AGamnehfKigojxe4t/gdmgziVq1uVtIc35stcpnS7U
XkpfZ0uPqogkRsr5Htgj4rReHzmQui0fIfvS79/04odrTYyTzakx2cWkl1rkTjAl
nC6Jo9zTgkVQMwFTnYvrzhRx1ESzevuUn7QmEyTN9FXXwTbGuuN+6TA8yXHU+VG/
lZxy8vUWTD5td3txMQ9l9YDcqqNpcbakpDFoR6pgDiGxMUi0pBba9lF4lvyNk4PK
ITNgpqKqAgy9fkNiCAUDWSYBT0h5F/sSXZ9ZsgVi5v4VcCojdIPB+tbwgGiWqTHC
EhUnjy+ukttjCcAqpZM3+5PKEYyoY5Z2x81MGxKkgyAud5S5APLXMeNV+t51M3p7
lnd/knq5zcOpZkdePWX78nGV6PMn//CHYw56qF+dQlU6sH8qKd5cwUm80fYuPTZz
bt43StFrDKqV1hiDiMuT6W+RzTOmGPI8/YrU00faMEh3MkhOCVl4BRI/KqE9H0Lc
mebTTc2Gq/zfK3ep64XVPjC5P9mOk7ReOpLPsRYp39CGXbUjkg8lc8Nu6IP9jBNs
yzJBvTMDFWZo6x00xLNuzETSsUTRpHpqMR7ZkCDVan/8yMkpbwJtiIDl1d2a/5FW
+HaJ47KGzoE3M782J3tcf9ETVaBeq43c5TED6MOS/fgMcxpGaKFltrxB+Oz0E/St
5DJTVtKNwcKa6NBIlRpjM3tEmSiT+fc6rCtPK3ClbBK4R2QMRNuzeD7csyGB/e8g
cHG4CMI1mJV8HuvO0F45XWU3Z7rBXX5mlliStqJaXU3MuJ+NVwxpupq68WVgssYK
ot2QxrxGZn1g1VjgXXqFpfd+Dp03KEKvEdfPABWvTNZMWkwoWfexDvoDx+iVnXIb
lLWuAjtqEu1i7MvcJ4Oc5aORTdsjTEzKVopRcFRcodTKXP4gJpVhiBupJV0TA9NV
PyWIKQEdko500LcHtWjhgEQN8RnRiZKOXaRNxJ/TJAVZy17H8aGiY7XRX9KbieT7
rDOJPoX7TnMi7crusJdAET9KRhR3LLoykG8d/Z3Z2V2pdCYBRV9InDmxvjhrCV0O
nY8/KTtLMRhRTiiBcdRBNZRL2Y6m0phL7rHwf7TkNIMHkwpl6yEltqm/S7/t1mEu
g/alzP5bmUL9tMJ32n4dNOxlZ+c+g8WFX0IHBoE8LG65CQV1m3kwas9Su3vihnLy
591fTgsDi7hMT9+BkzykygCSG82YkoxwlrGXR8f+eTN9IaScLhIjjs74RbeDnXci
s1DNeRI0JfpLXmngrr9KflGYo+FgbDHeehYlZP+ibu4AQTMSZLlzaEUlDLuDq3TN
3LotaEemQQt7+zwHEJVSvG6uJLazptsgd/Jq8RJKK3ySCCRV/2iYZ2b3x67xx5pb
LAk8y+ubzV4Dkcorls6m3RBYzzbmEqHjgSHocP9EhK8g1K9V2tA5eQdqaXBC+4Od
CvTjWKl7+XnKBX8Qufw2hiw27whWX0X/cATuYtpDQGvpSOMzYdgLs4XY1qXtecEN
1TweDBAbowgZ3AtGH85V96ETobZtoLW+H3l7uUL5Nrpb0uSgP5GrnLMHT2GDcNR3
T9Ae66X7fNLOWsPrmnlTv+j2jTsozyoBK8LvnjqJ4+GJcyJEcx4wEnNayXB+uPhC
WusVx5Nf2fy0BzKLCdTW7EMQ97q+k5Lz7ttwO1ppBXkdjPVqDWKmtIFHqDJCjenq
03u0C4O+NgoOuHrHvwMRDNJcCjiqb3KiZoz3scgDU5RNhC1nR2krsFuTTvRs4iMJ
dGi/sn01bSkkneeUuLJo6TmNvUoNu9huzLCItI0A+sfzLcCwOeHqMcGqopDAbqtN
YtG2mqlthFT2rpiImHiznzaq0wCuGb3JNQSnI8o+39yUV41iZPyxz4E4PQtrUiTc
G7fGq5zvs/b6/jI6bnxmzXaDKyyo8uuxqYVLaq2d2AGEEKYJYVMe3xIY43wtYUHd
0SOXBtdnrULbmrMRVDd7A7LWvmVY3H41MgEUSoBAnDwetKtft5+EL+80qjYOi8SD
oyBD5J2ttATP3RSLID/GqweRUz4w+0DNMhcUX6kLSv36jLfPVM2HHAEecMJwihVq
IFsblZzOrarzeZpMatAvNy+Qe5rKaZPASDJ6rTaGl4Tw8Pa9bHx3mB9CIsMvyt1s
KvyxKO1QDLwuguA0Apj/FyrcriOGI1xFAKANTbJnlGEFFNBr8zj7vr/E0iiEeowM
sO7qeBg7zj+SR2ZkAl5lalsMCce7mijw9VXGfavhVHETiT4LqtHD/x7RYNnawIKE
utNLFZc7JvF8NOBRHlUKDIQKTFu2ONmzpQVri/iCrHsYMzEV1mO7fObznArvpuN8
jK1LOTunobGM0luROTP71cF8r7vGhwmK5i3rkC699oCOxnCsAjB10SA/nMm8EAxI
vIe1z5qqJ624VORLQvC9SOlURNfujWBAgDQBtjM8AwES320P6tDzlWfiMQW3zSc4
P04GKZbkpS+/+FkIQJcF/b/4JSJJO95R2bJrQz7q8OOGYx/wq5XTy0KUGeG+Eyn4
Gi8+5UpN9iUouzGZzbp7SDcq/Uhfs+EZOVonLxlnxw50FdrJ294eIRs+fWl/L2gN
mPyGzBkMpgrqL1Kv3RIUS2zwL+zFRdTDteCCEP/JrgbzpYI2rbFZJSKoSF2kJdOU
dgijutZtjYygQtCSxYl9dLJZM8TfdfOVFA4srPdO3kayXPRg7zMbsn6wqp4qBw+1
A3Dm7Q9V4qfz3huGo2nSKOO995IC1Peec2owIZ8967Z9Mn3yYGk1E1uhnc1sFujQ
Uy5pEC+yENceWkX1JfsJEu5lATvLe5PTa0dH2R/uGlJdiLztejZmV6CY1RLDY9wJ
dQ5Hpo2gxNYxF0avL/TRlXd4DIzWrrcn+IZR/dKR5U524luivohRWYY4AwaDUljR
MTMh6nDeCbGprolDBAaFp6zzg8dSBCEeQv1HJZYIT+2wUuIZNvFOmrI14XGgfm/R
CAIcjBCH/wuUm5pR41VYYDk6bhVZ+XroIFwDJml4Drxo5DXwchko5gwg58ha+qNc
7O+zu2CGjJnGX7GCExbQrBRKqVre2D5dJre2HcAXfy5QhBwehKKSO+W33yP0qqOx
uKzkyOS4eY1sz2wFvxjWtA5CA1sd0dPUhuXSFXtv9v7iHzqB9WYLoWOvVIFyWwgU
PjAUGlwlg9j1GM+t00EwvlSW6XWy5p8ijmoDUk6gKhqUY57Ae6iccWEtZ4lLj7lQ
jZVogOx+bMbsg6zIh8MJmqIXnN/JMy8uFwhnU13w2qwhh9a3DGJw2qlXKmaia+Ag
CvPUA8gHgWi4ldozl7fdWxaPuSk+zzV6m65bxnmUYbpiGaptCGkUWjXEnA8nCfUm
tWo62Ut+uRLR8tpnzMcrOq59qV1bobs6ja+04vsq4e2OSeQyLsPl7SoqaaVRO/+c
7SC8W3U97jW4cRmoLqUKOea6oyoMQmf9TZnQaL897zGJW0SDS6kYvSLUcoqtXei8
/kPDE37MU8g0t3VP+uyxsw1mo6Bs2CoOal74yDhT2HC2V+Vayjbtsmg+Kd7EUri8
lntHMqSBM7fswvEScXNK4eTB+qZr7Pb9t5eCkH68UXmCTi+YmOiJI2JENZW5uBJe
HpOQ1GsxkPCjT5rzP8Jr9k4Fh/j86i1dh26an6HtaOlp1B68BbALMkj7sUACJKQB
z4rTa6fKNyaIAmeMkVAbkQEqwZstaRTskLoDLq9Fjb4acOvFfPSXN/p+LTC9r2/Q
MkvSJiD9ZXBAexrQxmlg8bVSQPBo385ltgY8ilCwIVPlI2aUEFUhX/BM8ucp/aP/
ZIStRxniNPwKdUFx0rvwLGoV/FpAHOkItDFwsX6tC/tOAIfXAwMmb/2hDrTzb0B2
7FV+zU3G9rISFRB5cogkCDwMa+Yn/uYXhQPmoMwykrWMpudeVp0VyYrrzynjuJTZ
inZJCMm6MqQEklCxeFMvNczf9M3cozeqWN50iFcsc8lfIbA/xanfxJG447tPxsSS
5b0iH4lS8N9FoyEiDu3QrResvfL4apTr8quDtRIAIecLwn1sVA26Mn92rHAHDS7v
nzRXkGB4n6OkrYxCYV4MZZnHZvfA1jWPrsAn6mHXRxXDIoiAmB/4gNqMIyAw7Kl8
P1o2cmke7Uf1YsU4+dD46Xb1W2jaNo7CTpC7zEf0IG0f8LLFnbs4iaMZ75FI0kRE
UzEz5DmQpGEIfbG90DrqMw7D5TrIuzLu/P6P9fJ2GiL4PULhWYnfuXpoGkWllTkf
3B/MwrjhcdqO9HPIXt/0ajJvMNlCr+ImSzy2TcYj42JegISD8IimS5z1X3bXX1sE
aT+xPT5sLHdRR01XZ0uXPOmWYcRJgE6byK/MOyY0A6a/9MvdODqaCTpTuFp2DiQ8
spM0CE49ZwWvCStvim1cPjxcKj8m48SSENHb09CsdZ1CVUsoyDKV/LDODssDngVc
n6tnRNZ9tszdY9W+MGwZa+CZ4/B7krTrORhl6mPDvzrnAq9uEDDMkWTys9INWqzk
t94vjcgTF1h3a0+IR9GMmPRdMlx7xS1v/YaBAUq++6us1MW7Jp/XHhRnf4i6y1I3
qxobAnzgaHyWETAyQnZ61+yEw/rC3yzxu7g7k+M49rk4EgQHkoNqzwLlH5bfY7/d
wFzea5dHbXufF1jTOXdgI9IdxMpwCdZl8j5PksVLZp+EmF1vXvLI7lqJfoxHiAk7
+QEwv5LtFiOFmtOKT5SjBIV1rdfJ60mTyYSVsl0M/WywOlEwTwMqyBevDRZou2gG
vJgKRI/4Z/rA87/8OaQvNoMtGb8ESbQ6u+vckpcwkWJ8VkvR2HTW5pOGeJpUYYOr
FjJqj9UH8ULPVE2hvcXLDkwqtEalrvbtgbw6+HikwVXxV4Q9d8Jhr3z6jfD1EheW
oUJjt8cIQH2rVDFTrwePqn+pMAo0V00RT3JFRfpcsPCO7mgvN+FVozWctdgFUoOL
zutRA7+aLNa/P6xR67HwRYNdzEvBgFXa6f86rFr5K9jKDT/BYxzg62NE9gTr2Mtn
pK+djw3myvJzqR3ZJtAWPEEZoH7h3zUf0UbpMdSFyp13dQFyg2hZeyh2kiITGhjK
UcX7gmncBOFaLgvUU+FWJegSnsgyh0iC0xo8BInPIFjDTIh8ualgpjgXiUE4qsVc
gxK8OZ5W26I505obzjjCnO62LfQS3AtGyVOg0We51wjXXFCHLEG36VdAH1wZTL3p
Pej40eIx1sBJ4PpYcDCDL7JVt+q0q2yx3aqWfS5LGs8hpV2aBOcECmqXzu6zabZv
gYO/2Bz5cyMCPCH4nZ9991rC3Fw5areXqaShuCpRWV05pF2Tfl+XO54o2mbj1MSC
2MNWtQFdrkuYLEqiuEer94ZBnixZm/elYLtGLwkCvum0EQSOs5ctPkFFOJmkZdiZ
5J9MiDjGv6Y3jNMQ/aUsMgBdR4IL8sAPCWKIiExbpm3JU7LDeDsdhDOjbhsch4lf
8uBUzNm35R8g41dtYhT1HTbNNdAYp3D9phaKenWKfYlFmNs4JWj9xAOoowgYvpa6
jtRmXyTgfOu+L6WxtOiBkSu+jhrGsqgA09bxYpN0REnlpMKkJ3a5AHO3QWc8eaYv
Dg4CsWERT2BT14ADiwkq+xVrMI8iS1JK3AQFbog7No2cPSR0JNe4Ntt/kct+ZSuJ
WkjBb+HnpGpOUjnqrzz9AOiGbPs/h8+caBVrFelRLB8k1fD2c3aFjh7Sff7vM+Ul
3xhzPjAoJoEnMTNeoCzb9+GgwbS4XqWM2WtAodb8jvopMkk0GbERAmJ2hPrGzTg7
ADizObHa9cLe8fRhCCHSBzY728rG1dIedbk3UWbfP3pZTkdkCXgnHEExyozzY83Y
eVwZXbP3QaxBHOfN9alcSO4RwI6VpmB8qoXSukiHQV+Ye1eXgvGpx1ujhyaUcYKg
b+Efmg0m7ei5OY3+ccOjd/QiTp0lPmsevHfuxdLN3Bxlumugg6OVZ7y7TgcuH/tW
NFRmsr2kuEOv4IEbyVrE6axRRCLFLN+UF+zYPZpOEEp9E3RGIeHYWR1GtR3PCyus
hxvaoqL810Ew1xQ+87gDWqAkmZ3g7Gp7komtxWh3sO6f2eG1gOs3D0P4e+M/ObVJ
rpM/j2KL+5/+OQ2Wt+0pZFks6ww4Ott6WuVJJrHwLMGrjsZmN5WI7vBurX3+9wzw
22WFiqbhdgEQH7wRR468Ilf68jZpbwp/z7bZitZUKMBWsuCRgLZXQjrrC9FQ66FS
wyNgaIb7PKyKMxLQt9p7QcBIVq2QkiydhMZvb/lCzF2SGxR7QZREA04Q2tmpvjWR
czgRI7eimZrrEQTnj/AfkzZjjsYrpq4YFSwUMhEPUDnPb/TlMsp1qJ7Rb4aRBFZc
lFyHCu61C/WL+pvBlZezmceeuOok1eYcuCitA9WbY2/xot1XbDQkU0LSTTSAXnnT
aMoUwA8a8CVsOPYrONaokjrAlzt8+tlX/5gMXglaS11wKXdoFuOnENgzM8VcXnZH
9qJQYaW9Aq3ugaZkP/VvX2pntF0kMFQC9UAdtqlXjk23ciAYGkQfjJ4AgHP+ue9M
ABPN+QWRI68yka1dkmUCFDY6JvIfVYyp5sQhW7+g8I12+9siYB/m2m+OpiWGh1xb
oDlBdc0WLcSoj0IxkelcSLOjCSRTuCDhALCBe857dTAleSa+xMbULx6qgAcGC/+I
XKRBJ1Un4Ecdn4uZN7ZGfkyObaLD6aeO9mH4pgmYA8BARVmDtZW0UZEengWFXndn
6WfwQ+SpeR3elo/L+hjtHZ40gcrE1CUF29XzHrJF1ZowkMxx6NH4R5jylEe99GND
dve89oJpnRkZtSKytwUJamM0vfvLM9cmCcTmu4jB2hxVCsIbLicibv4WvY7vKfuY
vCeGmhLqL39WEgbDIwS8Byuk5CznIjUcCijvLVEgYZYueci21Vv0oDiPpK1pYYJf
H9nQGr5bGNj4lGNZ/NxZIfssV9dOwtFq2e/edmgf+oaSZiCWHbaMeX2HYGLvM7hb
AUMQMKLy9Ixh6UKaXfSG4Mvl7sdgqMQ6tHNbO2vmL5IaPmRJtegNPgg/XKyc/m10
GKBjpQ2uHr29iMVZVtxhLm6uXHT00t4+K6bz1KqacjLA0dFU5s+7MpKqKgAXoH0v
oMymb5MY+2G80ImS0ByBxlUCgfHNw6iDiRbicw8FyRWfW5y3dwPQAnk5AFqkCtVz
9anJCqb7u4PdbOy2BOKOIE1Kk3vq31vWzjbBniJcpvfmBysJv+sT3rrubdyjzjSp
3dMfravY0xcd/iK1m/6tUWBOq6YNvhVGpTg89/+13XUomeFM4SjgnrdgmEE8AGiP
jL2LKlU42oczBT3uVdIyYSXhSFe4UOQIuzJESGhV+cBWPuLJ3iCVDoJLMlUPiusC
8iIXWE1zLcDJ3500o7dAdp3URl3R/rPjrYshEfwnT0pJAJ90uNNhwMbTcpM48Anf
HrCuGUJhKrKvv9ZsC/W7kumihscJwj4oHItTZ9q2DTaGzKTp0CVsAywQITF+Am72
RZCdzXsWGMbBzYuRPKYP7bu7Yr+zWDtjFiQdr1SnmUzVe6OlgRP98YygUWwMCqJW
W3GE89ShIl39vW/5ZD8+p7YyNKPDT/sLUqFTYAt4n3oI4nWm5/eo536xpUd5B8Tf
E8rBiEl6/Bzc4eQxUaG75yeSMpoMupQOh6catb+JQizgNOIybpOiu3UuUbCc7/kv
E4hOdoSYWEUSf2lU3oMNrFJac0OjMbM44DAurxHfmuQDc3rzQjx52mkw2G3teTYt
1jTverc/FyfmWPWMaNcAuEomXnRKj7CZWRx3crrLTFoPGGBaZ8LRq28fWe+2GbBx
6BOPS23kd/HafjqxJJYG8VLR1trLe7NfwgOUxZ4iuvCq5dnT71kRogRAafykzRSD
OSHTpvE3wUFsYaCZwUwflWHcXMhlFyopmFjm+eUEoAyDD7xwGDSyRCsgO4BPZ4HY
2cbgwVCiwHste4apElvXgXGQElMYPFuSa7xE4r53N3bvul04LeK88zxBdUiaUorp
x6SQYeFL2SL6a88N2FVdz2KdcnzbPoWwgDynr7JCOS8lUcWZf11YD6XG5dem1dmS
XW0r66NXhEatIWIdRc/0LQ2oEER4gcVfVRP53E4qZYUanAY48oJ3D4VSw16tI8wv
GE8njrHDcTN6jzxPOMFoFeMC8vndasbmfK/b/RQcu0Jf3qxlj8kTsr7jGJyzZFTr
+Dtv/pQ1WM0iUha2VUhVpfVVvlY3eY6nuhUbbu24giP39Fnfl4u8qP5Gp/4LpKXd
zOs5FEXXIa75yFb3I0RLS738l0uzFqNtk/RMelh9dA/V619Ho9zsZ8GuJJuB3WCw
UonxK0fVyWeSwlv8wzjfaBxNhdw4dTAvotZLF/a4pKzeDowDkgn4+ubtt7pqnkXH
wXqsz6sItMwic/B2p1ZpDKZdMTq9gNZlUZpYVtlKi456GpDqhVFi0jYl+2nSB3e7
ptn6gFOTJtzpBtzjug917NzI71eFro96hOQhnq9x5wTvmEw86k/xTxjfAvLyI+Nx
JteP/jA9jV20jfdoUlFlDHFgJAvmtRhfezGstM7xuFs3GNcmA3YeIyjvpspuaxWR
nLX3ODRm86KBIZCxDMbOJ31rldvVNlO7IGjSwzE9qthd45l+YXKdH9VqyRZhapiG
gCfnYHZdFrXqqp+vaNp9MdiBD3bXp4IcDNkFdyd/BWCg3ud/ul1XPHkTz8ldMMIk
CWLVd+j4r6MhQv75FZoJ/JyqxfrKqm7HWEyMwt6EYtZdmvIz8adiodpFyeevhX+j
Zd9AGcJRCmgBdQ4QibGn83xO+PfLcbxgpOAildnYW9x544tzMhpWXuPmmJCEsCSK
24d8rwgaYDTctZSsbe3tSXxNAG93hQOdB7At8igaUwNkMTpwfys1Wtm4XSE+MVQJ
03v0n3slZs3sVXYSeopC1vW75LCLEUj9SJEA5zN338FrLBbIHk5Fz4NHbbTQ33Jp
6jNkFx6zdZsasFNdxyKuzQO5nC0Ee+8UfVX3P0a8w6klTNIO2ij4hfe7tTHhEaJf
Uh9ZG3CdVzEQC5z/o7zaWLmLMT81zmyeaazsCx4MAhURZU1Pc1oneeRNcHPM3Luy
L8/BoRfh2u5+YIhOlEctMMq9OSukcTqXvczY9V6D6eiiu8/EbLtXyFa9CLGRTSOj
GmZKaUb5D4Q3EBrw2KZpngNQfuqaLwvnws/DjJAK9/xjY8y3ortbx2mE9Je2CP7g
VgGWYTWTmMdpA2eGfkgMpbQja3wCfufxjEu480cs/kgiNL+ImD5YMKte4RrFgCeW
tjcxojJgA/w+0iuWmJ7y5kh2AGh4HoaqCcfZf216kZWAEOZl0C9Q8kgLOrG42YpT
Fsghm4YigRco+jiU1iSuyLRN97xkRVurJeGpMUzJhGgorq/yTsxyEQHg/53XCDeo
RPbP9uRjIDjjk58bWp1BPJ5rLiHx4nhL7Rf8pMIOQbKxKP8dOODWadA2ZidZfp9h
aWe8s/kIiCuKHyVxevbqN6VneeqaMXtactP4bdlkGx6FhmpniYlib1KhWjOdTphA
sCeGdueXdincyEN1+Z1XqUKOvZQn3HWvyLd3UBY1FHFYCFfikjE/B87U4I3tDcZX
OccxrTj+sZunAGOA12qp7chdDfkCMCn68AePLyX9es4XNgzfI7mtnb9LFaN0sjIa
Dzbtc4nRRii2FiDuVpdyF4UQBGBJTX5XFvSWf9gGLNnUIxbAkEXO203JE5PLXBZ3
4s08wlyPg91fUbjx5KWpbJSgmq0ETXt5AvFz95hYgt9qaFAjOPWqI8rQYX7idle/
oancoVQcFWt7qxhIrRLhAVWWwg5sBF7bKshzSp1S/a4I4pd3yS3xMenhNrji9wmF
958Hu23F5Pkm4eWRLOekWD9aTuIldiF5ffVAOUHXGbaZWEbxTdiQ+qd5hEmMgCob
i4R+ThjpZeBf01qKj6TCC7cxfC8V9dpToffP1sU/vjr33kBfWdvRVhOqq8H7Ukgm
rrMsC+uwgq3e7uhI256R9ulkHhPbgw6dkVMqo6y/m6U7UPlclD0klG4kQpps+5SG
iydJBkzLbZu+TUu9OX48QGI6YKQUJOEO6muNXvKDPRJAaaaViwWwGl1odYjsyZCt
vafGccDSdvQBwf7L5sAsEuzHhg/trHv+LPHPKKDm2z7nGY032ABdMGcyyMnK4sHe
XE//ty3SOrKJqfyoUOeeJZz7L0umnaI1tEJ3z5pF7dCMuqaob0XfxEvd9oW1O9Nm
Q5cokzdNQcu+BPTRkJh0Elv0e/mZS96l5iAYjG7MrhCXMxL/IaYJHuApJxBN6sdu
gQP9AHhP6qWnRbr4rsfyirSzRtuT5kD4jCkpBrnjycceOvfJfeTgpGM4GE/qUyGJ
tQ+6OAFsKTqlyngFswrENnoErwJIGREmSXhO2QhVleO6601B5lpzmzaWAwUs/Tkt
AZvnkWy2AIFx+1S3VVM1lG90KFx6DimBhvRXPfi5u0mm8NXMbrw2hBi3+6K6z7YR
76oL7YWyzVXH0/8TXpGCmM6qWL3PlBr89vZuH+9thBgbyHUBsqeNwfuz/KM219ID
XopWU4cF0/8DAmLeuI3ODq/FE9eMDahdrelzw1Al15GtOOF1VylJxa7ezzbPit5M
opjd5roPlBDzlo/TQUtkJ2Jz6znrCZcyY96zPjVNxcFNZHN2WmKagasrEyV4RExQ
bmb/1e6MKNUZiJ524o78dLUaTcr0DX+u8ySFxCw4urbv5iUM1ibyKahDbV306tWh
wDtaBz4sEUqBtERmohg3GW9rWymy85S+3HEb/HSZIlFSbasJlxDcci+iBVtjCKB1
HRaoTyk2Ys1z/EeWHzbn/y5rGX+NLDBYRD8a+EgQnWwdANkAcYuP3KzjCLrCScBQ
nS/VlqztubLmTZ/qtGQ6ePHHh1S9JuEnYMOewHjVCQacIQCeX1D9A7++FtNd1jAn
HgiRI6s5ynhlRTN62p6epFlGkN5PhBxlMHxQFo3wWsvyLzWcnqWmWk9WzkHg7JyF
Wmn1zAifp/tD6P24cbhg50q+zLnXULOi/X2Ce8KevE80h/YFK1J5Kb8fxWW138VX
O6eQxqEKYWBm4TS4ju8MNhqvm/oQdaqdNmMFGtLXYht5+sy6+PtmKFCNpI2STq69
aZrvy31LKSFGniAjg4S9wgELWdhoCfC9Okl1lURpXX46dCu6tAVqDKlOcCQ8Y8Hy
m4sOMeExD4KXDVipC96SoRGTFLvq2VeN7G46EuWJY7SJmeHO6Rs59VrkLIaqHHF2
cwRYpkJpqq8MIy0wTlfuOT+DzFUt7vls6YyZ8dmeY3+n2zvVTTUGSuRjkmRRAhhi
k0IfFHLtGStHqdWQPDiCleOVXtvfI1DCNbXqsml09yo1bbhB6UpQuXkoGM2dLHXc
59r78q0O2DXprXx8IAELA6IGHFvWA62LPIyHiLkOUeWrLTXOxPuLgZifpWcHp2nU
3bEs1I2lsaHedo3KZk0m+okg2PmYbRRi8sXJXjEnPQ8AyW6carJvIewfbDU81RuF
Q/Js4zRtldxqIMRREjWXw6eaHLGLg86wHMmfE3yHCFDm1veVZ+SW8rE+IKWn6qjb
oxbX32xqGQRe4nAgPnFSyJMnMeS+aCrLWrFQlW+LbpxGZTV4OIaADiFKHT6iOqlH
Lt9yZQsdj5Hr3x1p5ve1HoI22kkDD/MpmLN8mcaw4CSVQwo11l66imWZW/vviCw0
xoAvb7skS09rWmlTpYZb6ZG9zswHuSrSrMuuOVmAZz55Y4o9QNbmFCbNWNxhg/1n
yPZnUq/8q5A3+9h8xjUrG1V6CxYHR4YhcErBKPO7b9WoCJ8JxRtg7KhRj5s2GXAT
p+sCHzRKNcOYy5NoQJCK5fGVJ38FMHxcjBwhd5IqsRFMmb1lO7f9JYOITfqSipgo
3OVnwRjeyJdtUhn93HTBdeAqI3Y0N0YFQ3MprI82AVb9qvnQfMztS4lO9JXoUn76
GYuYNuDfLGG0jxGWkGVEgyE6JzxCKF+vfLTxhA4/yKtUaIkmYPC7/fZZv0ssg85O
AXV/abrt3ncoqRWWrQqBd/pFdbFRZ2ahPyXWwbQoFjOQwIqLDr86m40RwJJQtMjy
EUI7HQaRWX5bAKk2xMffcldAQRTJhQiC8ClIb5Uyi0OEoCHbVHhS/VYKq1ZL4d48
WdWhIkUDYjGjih+6HnGuePve02RSOTz6YwrHAZ6Di4+5a1VPS2CyHX4tTqoY45nx
ZQtzcRnn0ipiUWK5x3qYPcQGlYyiu+md2skcxwDgumSCVDUKgFF28GVSoYD9Jj4r
HFlO/rgqDBqPh2OG04fpkldROh4sCzowaYbgVLw7uL5XkdtWhIojRhd6Kd70TxyK
AeF2aIIvFwV5TKNaYPPfcSLD9QGb03B0jht3OYJdIiCChfqFMrIIxeaJGCB36IcK
nBL7UuK4YRh365DQ9joDmiklMRP9cbRLHouzn4ktUyeD0D8o0H2lAjOgIc10+5oL
T2F1lgJLoHRQrzJ5CM6eSr4RtPbwnvszXlBsmnF88JSjYnaB9nr7s56QF2JJuSN7
vfRRLMFMi4RI2JhTU3wd1wtW1DQvmSPDhcXbIWDOMGUAjQykZxvasqbtYQDN4auX
b49Zlj9FvBOsH9T2bGZA1Id+THjh8AUkk+Wa3Gxw+/jIVPzhztYpN1BJxIIFSxun
z2CHXoJd71PUPclz4EJ2eJsaXJC/KWo3jtOpp9d6EYkichq6wkuCXZWNYk5itoBF
+juzCa5VfecQCv7I4AzYc9naFEeX51evIVqGLRBi3JAEXp74yTK2IxYg7YwJ0mR3
WYjHs+g/5DCLYkrJ0wdpnvY6OWOK1MUTk5Do+/I7qffLTxIlDaB5zhOTERCtbg4O
lrPYvWx82xT1eiuCTHh5MidFBVNrYtOXTI6ntDldO0Yb2IFW3qvrQXSLmMvo5K8U
CRHiNcVQ5CCVDL5r4cxQmO+H26fUg+AgC38yelCkVy6gKjafGy8wg5T53CMkVwGz
7NbPIrBhNXa5IfEuCUUOdrXqN2HnF2SxP6PIB81TsRkYHvfyg7g2SDjx2ejSOCIG
DOCtnZz4P5wr89GZcDH6zyMBa7ENpi6HTl/GXYROg+UzQPuZNbxsucTRB842FATy
nWz463y3QEQdln7ysL0CaGf1mRTzy9M0brosD00PFYb1fhp9w7TveHbE+FTmSEwJ
dijnvg7J69lImfj+MnM1Jz16UaKVVqYH9LV8cV4IypXZ8jlV/Ue0e/zw5K5ewxw3
GnRbHE+0AfcB6yUXZ9ROmp4CGB61s+L5T7OMTwlwx1WciD4ZzCTEvIjV91ncCUll
QIDNgBWMyP53wMx9q0gz5uDpiiyILcnx6BoeUZrb0JI4kxd4YbByj7WCrYwsLefP
HSsGOtiULPphX8ub5RJbu79a/icBeP3AVE3rlXEdWeBAaqnvao/ZJYV6RMztDcyl
Q/bQumLSCBVL22C1mCH/ywI5n74ANMMlCsObH+alKwgVhIG7sY86LihPhBwzNfyz
AnOc21HypNzxJQ1WaTU3rK30X2myDBHrFCHvZ/5bn2DiPSHYKfJ4EARF3nycBTgR
hitaf4/tgLPKuZalNM6TP7qmLNL7Af9bkv+YCerM7vZWgo8iJ/8G9yfwJoruqM0U
Vnjg560UvMnmajWXZZXC9AwmcnLRTIIyytlWgS9YlerMtQcSVnyZ9+nb/eIqx7UE
3g9CV6iVq/Yq1dvLAXJDRvKP/3xc3yWlPPTdsUPj9452yJZ/P4KEK6svNrRsvztX
A1i0wqHa6eiTZic2safQoKTw27Ua2PrV3Tjmvj8Q7rzKHurIj60jOx/2sOq4hfnG
tpJA+ByhfXzVgq5hJVwH0FxP6sR1fVi2CmWIjxGo20l73qMPq6oIod9RnufNyb7N
wyKpUtkWoQvpMHPgQzI88S1GokYafE/qDgZfA1fkbPoJT9GjrcRLtSbyDm2ls/2a
21rIATDgf6ji8KcutxCY825N488hFpIuafSr/vZYojNdoHCycD4OJERZd5eGRmjK
eRgjjq8bTgQNYt7ZikHe4YAIOqUyWmxkOz8ZoAxT5ginAJnG+ofUfm78QfNjHnCW
ryV0dkKnPeMp9O4bEN1XJj2KePFtLomBjdh7yWBxj8pIsXrLWV6XqLrZxyDikCFh
7+30xOyJ24jS1/wl16VVoFrOCDejDga346xWNowDrjQkhFuWqccYiPFZhQ/X7mwT
AuVYiYLa8Tp7SHo6RawGHa0XIG3HS45x7IXBFV2ih/X0+D2Yd2KqPoo4ukhJMtPl
QrdPTOkbHVqDvTk7VlutmJhyo0XU7VOx/xA/DEdGKxsemuVcfIcF+WNlA29Tl592
JgbtbHCZby/BoNeu4Sva2L8CEQa4kAksQMI0RCb1nIEuSrgY2MtyMitdEYm3J3Qj
ojF6NZGS9Z54tbo43XbPtjuM2bFFG+J3tl1I7ydw014pR34zi9cGdXIf5GVxt0FW
qovBn8zY/Otiuz6Qs2QNLsUS1qO7Ro26AwKEF1TRgtsHhJL42uh3LlOTsyhJe3Jq
FprpYBkRj0ZHdneo10qdYeoVnd8bPO5WfARpMdoXkDecMlSwlaHlULiaTuk4J4nq
fdhhjs8wt3hc+Qquu3+IRK8MroMTL3Jc9PtT/yOdxZVNczJaONUv3Qtxlm6W3nEO
ijwPpqxEy1KWzANcr9hce2MGnGopYlAVJnB+xMaym5esfv22AT+IX3QcmNQ2f0Fk
0yp7kRBs2TjZghlbC4gSMSMduipvKE1p0cAMVucJQxslINF4Q0WLV3Zhx/SBvSra
K4k1jsJx8k98VKpqZvY240WRhQrJOcj6UbBluUQjxy22Edi2NF00PHs/tjlsyYbJ
plJ5O9zczz7OW6it6SnnUa9bulB/Ow4NW0bNe0fquq7/wuOOjhxSxwhraRd6LuQz
1UNeMRqvEfu5AqOPBy0fY36CEw21X/zCPsbWq+elBhpTQYHb5r2NdUI68agJExqz
N/4paWqEwQMykucZRjolp21Cs+7Q28qntwhosVhPuOJqi+Dtfz/vxVw0aRgDrZHe
VzAZLvWswTJX49cs83Po7WL0dNSm+K8yYqh+FYq3THo2NYCM+i4qc7dcIABgja22
FkU5P/BVtYeNq6G8OehG4NRNP2IG4CKc0gDytCR/abXwUFLmwgKn1dVNSZa4yzEb
5dMEGHuxIhwX3/PevCB8jOwNzhEwDF7/sz153gm5xD9RuWDkrvPsrE6MbtIfaBH0
AnJ/xJUawHz0SJS0sYZ/P5mkHVCMqB2QXsLbPG/cEhZdxp3CNOW17nl53mKjXQao
CFQHj1s8xQWFhwnXWxCdjqZHjzg9G1cX+6GVbVRSTaTZH2oex7WBVvhdyBToORew
CHuAewxS4gztvFaB+yGZJjgOM6zadRHccTR6bzBtto4xI+xl6HCtIq+YGXVE6B6p
3RaCOJipspqLS1Fa0eGv/6ZTk7prykglGk2ZLJKzhh+zVklImjI68hVr7jna4Eap
OfM45kmkYwVU+AITjuxPhZHY3RyTcy7VLFcPO8dCUUCkaxveF728n0OEr7NYo1iA
01lPid1kVBj5IiRC6QmEdi+feHgYGzFyv0acm/MyrjJuVmfY+VGrrtYgtogVyYOe
KM7cuoUcFgu5kmEscsddtCDC7D5kztXyAjdDvnFzbVAXJVDcwYYY0uTCVX1VYAHV
ikMHVbsXVWEMUvjt9Z6NX4HLAfXmPxbCMkXWQU54QdMAZO9sUXgQTxmZy9P1Blme
UeGyIkrFayWa6yiprQbbsBmOJuCkykPIPY5tJPJ7CsPes5WdYNBwelZDcNytXRAs
jfjAp3Z5xR26M2AFBUBFD8ei8zQNFcdnNQAUADQbeYPWlEj045STQKFqcGeky/Q9
S7QWvN4dmjRuwFUCe0Sc0nc1T5pSlTIUteIn51yWfjxjK40NM4ZAdlv9e7/On3Hl
JbQYBNGodf6T8vZoUwUKTHDiDwtgdX+h60R/BoQyuoT5pEVgld/PE3NJDX4Y86zl
o6kMUbfxm3OZKIM0qaWmUnP75c6ATmd6gp1+KMybY6eEwPFEdOlFVNkt3kUcnXw5
WVk7ErvTeQ/QgNbhGicvZwhJTCbZvpTGKmNACVtHcBuJ1lKjuDN0cmH0guB81DFw
p4s5fl2z4eNrY6fJJUaM+06kIZaQY0asDsWr1bdTtLtkZ9yXFqDEiex1ElpdObmV
cXGjBFF5p9S6bpovk5GBc4UeMdONMimc4ct21seORAw3sp4PGvTIYpecfxJOsrkI
jE1i6046+UGCRk5iRjWimYr6OG01yX8ZUR5kYUg85/km12Wfrys674OnYQTFge9/
PrIVyPXDF3lF1qaDldWvany95bdaA8VH44Vuz5epLHWVY0w6beodRxE+yOaErqKn
CDOP/zMtYgoHIQ3r7VRxSbJkqNPylc1M5P5sFO3vM76zhpaJSjnhSrOYOpgu+ahq
F22BnedBPUMPmkFe2yFqBjv2GhTXf6fYnj+BTzuIP4wdJibBVSJD70qHU6pM5qjr
kqIcJzD7PWjqW3a0vR9HViappraS1pxUSecjTyQ6ASHpkSvnK1RZAhwlWGyFf7j9
G/qNTmCH1oBu2WBZTrSzH8YEMGpiw0542hHYY2yQxwwZkxiZlLLWiP64voxqVNwS
/ROdBTNR4MuMF/8RciRySjFhwTMzyvBtF+WKPsUM3tmJU2hKwPkVQI6fPsKbW+JB
vdfpxBGToVfboH0IKMPD3N5NAxl4fKCAp/ol2waU5xisg4EpniZu+YznMea6XHmS
djcXbI3zac8BezHMLnHVM5wNau7SUISrT89AKri2DY9oGAUss5w8cyZOwbfr/iBy
nZw8QmixpmRi62016GHRfYpCDH9mievL0t+AsAW4TKmve/rLsDuLGLY1B8HNXUZ6
/X+q50ULD0Jkatwq2I62h/xG+Axn1hpCtqYvusavvBTb3UpJN4tjtepW0eejBrLh
VJwUpYjp6V5jMzoukquo48rai40KmiijJlNe5n7TBj/iVkNGnevDmC//sSujmKyk
r8wEjzdeu1a15ntbb58Str/KNKbdWr6qNgGtRAb78OaXYX9erUVnsH8RV4UnnutT
+yhBCl+3wQVTz6Iw4ArnBlsMLvpwW+z+rgEo08xG88u5NIFZ7Y1j/Bcc3+09cFC8
NdneCGUZxg74WHpm+CWuFpL+T1JLNVRaQ8B2JF+H4n8tS1mxZZ4oIrs8963W59yk
WAaGQtJFoyoTNSvhLhi0xhYBijNydueRC3AdXeA8USajCVzVC64w3MOMA8VYt5xy
V2hsiIKn0ZoqjO5310vpn7+5+A0CMc/hhLWVmZ8Jg+iicZ3i10mKhxAQFZis+SbM
hvYRyncsLqIesehkZ1zPa75jEwfkJwNpR1bIJcs6CpFc8khAvakZFjtt0hC2JqQc
jILHNqcm8eplIDbO2XW9j1RBtTF6PDJoHwXu8njAsS+d4PY65LcHD2ue+PdTvda9
RMcaMjHMYm3mtpOsD+8rhwRNNhkrbNGm57oP+20rHEfHDslAhpxWAYQjDpZIlRsQ
wx/Wi7+kusN/dbviIkuTpyU6p9IcT2pwJCfce+Fse8MowhJpvrg81nmcyGwWWUmL
5VptWISmetqB57m8E7dqu0PvAyQlTBwbzv1kKalfvEmZGss1XBT3AVriB6UNi5jW
bTMr81MeUHIx1NC5Q9g0OvpMuC2E+8SE6gB5Ybak+5pXALNcWYsyWGZh0iOv8jyi
4NTqFRe72ekV85TIka67O5ZrEF60p+lovYlY9s1x8YW6AzZEmSKkKKKk1K9Wj/ke
skC8BxjBez7ZxD9RjJ2JAfauQpPSIwsAp8yT0K0VD1Zl20MKndQFBx7/c4FG3yr2
5e1v3keEhOULkjVRx06RVpVGRknrly7vuxdbFjlOBYkQeZfVUr265OEkde1GgxGS
MfhtDM3M87ukARi8HITZ72oewJLc/bfw+3r7XrRiYe+mU3h7vPQI/yC14lQbBJ2S
lkBkKfbIeQTlappPFiuOv/Yq9dRgC8mbK6kbkT8qTmgBFif9PXCIUoswMoubkJ73
V3yJ0GLoZPYC6kstR/h3XD6abGq/l30O5gxIYlHvwjv0aPJgokbOVPuNt8qxT2QN
7xAbkEjI5Ze/kgU9XYW6iSBzu8pg+vh4ONXDrL0HMqN8UThzlMXZqING/K1/m8Dj
6h9ZfLIWbi33gAixPLWp7e+O4uc/wrzNN+pRRVcId5PRp7XBrqNI6MIpsCcL+58R
V2VPuA44D+oteO23vyYdwpPgvGn8Nj3BRghFB3Q18msGWOPeQ2xa+74mrtPc9TwI
GP29ACMR3LUpZcEqbd75tbWXmoG9PdGsShfNHnZoqsCHoZ83dND3Epo2q6amuwj6
5gKkTvbYh/LYa+xpVJlgIMMJiY0DQCCZHJuz+Rg8EmsVgB2ORia3HZ7uecAATI0X
LTyDpMpIT3FAibbGvEOL0H4eqpsULsOFHWMzM61Lkr4jiC7yCia34iyX7O5upKkq
kFQqQ18rYAHYtUdRhvvim+Uy8rw5dVqJL5iTv02+lExhRO5YLOYJn8Dv6cPbZnuz
m9+GsguZjKvLaAI1Ig1tumLspgW5PhP0A8XZxKlCpeyQRNOLJM1SucYZS/9RAKMT
nhrrypRNHSMHcbbCfqOEMhZA1YgBJYx56Kn46xzju+Rrx5rOSCKS/LDYGUlU/kF9
hYzjR+3tZj01Gv6FR6snKdhAOcail0MEV3kGNoNXmfl1/gTGlIKdG+Wa8zvvS1aj
dE77HtI7Bni9hTc8ynGBpWmgsUxawjvu/kJ+ZFMxrGGPFvbYMhb7e09wlhvF/wnS
uTUvUO47ii6zve9+IVV44CMN9f1QvsxO1JK3rjp2uDU1YJicvW5VsCj12YaFdtIT
X6raU7h13G0ECjFHelUnuOQedrap+NUAzWlCqN95P8Pgus+w15o+1XgdKwNkgrxq
ccK0iAhpW1xkZR5o/tU7QCdGvbzqlMKtoC5UySpAwhPqp9j4ueyhZmnKG53M8viI
A3hzdFS9gtxu3frgTaPiELt1+IYjYdqWc1fvNLXcL+s+IVGjyYWSVN8tYa2iSFwP
7Su8L9rWLJ1mc2M52z3eNuoDnFIFGxj9tWfiqhKODQDwcYSwi91RmQKWxLPBKN2E
MYF3TWSDwOIMOZEP52gsZ60GNZ16LPjr71YA2J55rSQivb618e9YisyV0gDtxsBL
KXMNrnn9k+qoUleK+KEsSLfOJ4t/3q2O3dNvKdrARKpY9+ed6PCUxJBHCJeHonty
lP8FE7Ddiy7jlTlyga/xcrCuKLxG6G0AR5ChHh3ui6LEuHdBS+qzxLgRHDd7z86P
/dc3xHDKjdLwMfx2lWdyH9Dr7o1gKi6vVDRXQ3bdxUVbxlBod4Q+G1/2OFQ4krBH
8TYYA/Vx4irGP0ZCDVck3WNYnqyj8xZSK5IvthHvbQ5gOSTPG2/piAuEWIqSKJ3P
m9QoWS23Aj3m6uGWueJuDwa6uW0jWNhv75RKZcW7CMnf5AARWPPhKFNOj+RBNn/F
VlxCMs+mvbOzrMQCRAFhXHfp0iN3XB/sKXcoCpcgcsXDx/KBrrYQD0zm2ZeALsUu
lkl2aiiKebk5FJrloCfU0nl18Ji+hkAgCzGy/IqU94Mzn/UMHv7c2Om4Ys7FkzzF
jhVsth02AzVQquWs5RE6wNDEzlHP2amDfl4I5cf5qZA/oU7ngRzjiwmGv0LhOle9
e4mBe9aGcNC6b6Cf+dD95t0HgJ8KZe5I90jP6Vc8gU6ObacuOCUEFvoNIewW37dL
jE0LCjt82cLY9N0/oO/6IrbrmuBEtANOYAc20km22AVFPF0wGMIC9Fx4M5at0tgY
g+FLe8KBTvSSqd5GYQMot5wbjyNXnAVLq67CN+8AQS7K3oFXXc/J+Dl6MO5wGh5d
uG6j8ViIwhXkPyYWw8AAV8DpSvSlvDLHfZAZBp1SAdBg9oJG3UxZt4BXmaPDREbk
E5le+ic89+4eVXLmLvn2ezC8fhEu6DytPwTyiLuTjwrsiWRdqKokOsU2FrgGUO4s
qeLa0RK3xN+/BChUGgGsSZKrrO/O2QFiel1B/twNGGvBkyd1enqGHYuPWszq7zv6
xM3+E330/xw4d93tcwvfm+NpCafhVrah1PB09Ko2+mipixvlL+gai6QqkatPOBS2
1QBc24cpc/LDT3it55LqcJ7MSzGqUmfWJpAcn6eEt6IcRC+XvtJDgONGR0S5vpho
d17MDr3d+zAywdP29Mk8f1ZgTxJcj4nISrOEz7cvbJh3GyNuaQ6JgjcTgzV9aMEA
g+OHZh5lM+Js8oTqXGb1myWDiDDO/w7ZgNxKtYCEELT4dIN9RUYQRuu8PusLvwo0
mG8bgBT/ObLBqIcuamWdZaD45Ppj7tMFnqpx0w5KSc44n9Q1tCeOVPUqbzCmTUO/
9IDgfMiFcFv4Y28FwmX3mmtj6Enaj7TYOSDbtHx9CduG6E5LswxNRfAroiaIB/nN
JppI1v/1tSFisB2IZuZO2Jdm3CvG7k6kxfsOlYThfWi2IJDQKW9mLYHqDPZjdNZv
Nnhkd/clZ0Er1Vevw/S6wLFZohD50hV2nyQx0zWQoNqXINNgnJ3YCos2vfxXBZcf
M2M/l5j11ydGs4ULsUdZaT2i6HhQLZIdLis16dloFywIf4ML67BW4kbn3y61vJvJ
r4ha3MHiYp+nuAhLixuqa6vIxHJ1CcLr7C3YrhGfOo1UpLsAkrgJCUFHM9eiQsDs
fSPt+tNngH39mPWjouPxzvMNVA5TuHstHsSh92JiMnDp1iJb59S1+odX4eTm/7Yc
r5Rfs8PDRaqWULb8s/HM1LaLoA/EjELGqFbBzFKLdPdYSbhQRFmF+qOBEjsg9I+n
8pe9+bOEU3Kd98l+ISEpP7mYaVJf1OZQiMehjcLhAFJ2IAgKqI2mOqKq40JjawCy
U602qoejgTIWHcRzTM4pTaezknTMvV0OutDUvXmMBCPB1+b+sIWJhVogNpWiQwU4
cg2bcXxtFLMQ6/Yc0orH802g+3IILVClUWN8NgzrIZHlnwMjdMk/7K5z35paZH96
P/hg7DAda1lA6t4Ohe0JoYNc/ajeUaAgn5vEzCyomuBc6FmA6QrdrHByWKo3d2+D
lFnuUdKDlKaa8IG3XAxUQATFq92TV36daDcq3vlKJioWNdBtXJI2Q+BNNsNiYJ5i
OuEEZ6Z5CL848fhCNJRM0zfWFNoF1lEZgAezbt9R4WWmYr1/o39tFshOXAT4gCbl
/95O2aD96wc20FOT3liM4BhwmPtylPVAy5wu1j+buLJoNwLA3VDlLg1upfntlJt0
Y39dAYR/vcmEIphJ3zIdz7O4bel8oC8aW2+BEm+TShUT1DJvtwo1nBURcdVGoK+u
tUul0aLJi0uLcVSdeSA1jmgKnqitg776RLSsEKg+1FieSyUItoIqBu4vsxHqNQup
EZiebC0k8vUv2eoXWvpAvAu3Xo9rnFq5cAEU+pOZ71dO9Lt+a41wnBPdB+h5KpFn
mHlnYLmUJK9en0mvcoHVkLGAPwqJ+bxcz+aEBwkEtLiPpxCxteIshEYQ18+562HC
MxkMmU1O2A3mlOr41H3LoNTenWyvUP+VZCgdzrufqSlf0ouQuhVzs//SkAfYuuA8
mtWGUWDPDW6UNaYAxncPEmxwz/re4xpbH7rC6dJirVU6SbrTegSlOkBvPh+AdWx1
dqwFSaT+WTawQVweBhBOYJ/wM85sbFKqlNB/iaIiHeINPpCtuqWU5HMXPWpM3PK3
0E+PPDCrbpjw4bRQuSe2lxgGRo7pr4X+Ku3FZfnjZKIFv7zi9Rrzznsroe29s799
dt613R2ddJWEoKVWR7hPGz844IC5dzbVsYYZd1KYBOoRdlsrUENDIkhGqH+SUWhf
bmBHKJK6KIUHwivlD9+A2EivH012GnMC6cvnTDTgU6UJHBitc/QZ1D7lFOcRvSTi
EA3tY83Rnka44M7JcMfFk1kQrqvoJCyaEsmodAYdmbv7EyxkG8P/5grOo8B4isFb
MrOauzo47QGRXaEQ0JxvR+EpIYDQ7vwrijNSxgpO2SKxXmUVa7eSBivrX5MqtnZW
ImP2suYS4Kfj8U/gfGZiUeXRIzOH3QTz3TtIblQ+TPcBkv/uOIV1qi9et8XT5Efe
jkCjUJVwribKF0AShpF8qFJWww6a4haOkZh/34H6EoQisKbvoyDpegZatHqmRMIX
QjXBSuHXcBrqkTaCa2fboWqAZxp8CNCFQyMlxBqDq+aVh4dGTzTeetcCj3eVLif7
SH8byiC6fSY2jVB24ejeNvXoe79kdVwXLqiIGz7hrfQdsU/aSch4jh/G58bY9pVb
+fzuhwpmdmm5GQ8do5vm8iS8OPLSM1ZyQDTPO14cdGp7ePy8Jwva0hh2pRvjux/y
OjzCvPkLTrMJhaRTZSecZnmGARHfDDuMBG2MwkvqiHBa2a/QWEvcyQl05OtFtNL8
N4z1HWA6U18v7ZZ80HNAfakJvjCsXIITXlfQfY/lGvNzBuqGBIsKJs5ZgZESbeE1
cAzhr+xrBuKzFQecuN71Rwj5WDlxaXrAynh5dDBotmoniUplLh4VA3yj0K8pP/KW
6fo3F5eNQBS4ubWRTz//v3ZKJ5sq2XANQIHa+wbfG7JByS3H5+y6Im3acTSslvB2
jDGypvxeKUHs/TMAvGbW/ZsO0qEAK9Ex2xE3GXv83IHAp787Efw/bUqafd8VrLke
tmJb54W8AWGrazRDly1EO6gjf/F7eFxND3CfyHt41wU/+IMn04UNy4MNt7Uw6ox4
ekDd2cTtF7Lia+5A2rw8zV69IbTYS0cPVrRndxMltXvCGFg8wLd5aKw7h1K3MJ9E
kS0MyOJbCVcVQMc6V6eY4Y4d6/QxJ0MNu24ppAc7Hq/CfYBaitKtSZRJfFqagqd8
WiIF8gWfOFSMY5Y5MCwBvyLc3Lc3CtmSkwYjYZZhZdb4DV+Mw7msMKa8Ejj65O7H
vmXoySGRuR1N1yMr+sMk/ZtWTl0lGPtbocqsSFebYOa6yqFkqzZGhfJx1+F7PCFB
S9t+hfgdzWXQpRFUmBeQnGjvesKy2opixGAWi487Ay7pZxzkawhdmEU2K5AqKL4M
dxN3xIa0BruzTNc6r8rT+rNzk58GbnRh2hZXVwXztrJZoEDItlPDcod0QcEJIPfp
VVvHT1+81aNrLWvlPQVIISiNH38ztLKOLflEPJj9BU6coyiTT2LqVAom9wBGH9Yq
5cFpfBWz72aGJZ4FgLfDBb5c1ox/X3tGB0WVuAhILOt34DieThtiKJlPZ9kd+6QY
f8Mx4mZvc17x+CIecBAH/EqH8DpWBHHAUCeAH+iZSEKiR2ah+d18PHtVBz43Qyqn
evnuUEtFL2qV7KGahIJvQG5S6NZRcK+cXBOiCkIXQCmZOusZq91v9B44JsGzKSNp
NeeWhOShFOsEkyqB6KIK3S5sW60VEOoY1N2qFwL7Q3UITp529hCGPKyIYOqdFsJG
M88cQFPrdoZeBgNxIbpLYgpIHi2XPPyVSsY708LD3fm0To4HrOLDYLzt45t4o4c5
7FnhFnnyXtC9DBWs+8kW28z6F57nKFypyT1gDe/UKSykExbGeSzvXUeSG1rvXZ10
NzvBrCC/MUdZlSMIbigRdc+kl1OdF7NvddCVm9+mg+Dfp6uA2z2my6x/WsVO3tvV
otWx+zHHkRkwPebTBIAROn0hZe3+tuHsfj1krQ4t/qCaBaznJqtL70GGlBq8WXNE
ZUOBtU8zjFnb4184Sjl5nyqO45vD9H86+wYqNOdLHfLzvpWxqOiE+F6wxpz20In2
V9Z5P4rNz9mQ6WvupFUvvQYte1Wra4H6PzRdcsToSHNMI7TxOmo+5WW23tib+9ms
Imw7yrYlxCGhyH5olm6BPxFvANZJp2kEiSrSm/aikCM3jhHlsPn2WEpI7m3K/xzR
BJgMKNX25s0GF2fyL/WRKcIYJxEQwD7QJ0LrGsZIUQj9GMNLMrir0spdvHXa9Vl+
80FuZgz8RsCsjpTIfQlQBvDJJt1wa8zVaopAIqaAPfhlxaBJXcayeOYXiku9qwvZ
twtxlhEqGm+ClSfOuLjgNUbEczf0oR/wxhOqTkZDhPtS6ySYZ9VQ6hp92j07JvGS
Vw0iZ5eeKqwK92zSGOiNWc9SDNEloHRaHCkEZ0k/Fg0AvX+mOoM7lSRdgn0Gi7kc
BK8vrOopN8F5BFl2ft/X/KFH2HsPpq1p4PhKFTJgvJLQ4f60byalo3RBHaz0bxJX
Wo98n4ic6yWuNRtIQ8udPpLwVw+x48+6/eZGjQH3neVefCKmZlSBRRIW6vpbawAf
+mRHhqU1hdSy2gvjr7vA4fOPm27OXvs7y3KJtFWr5B1UyZKeunVmawIO8nTmcpyB
ymEav8BSCw3T1uePIqOyR+Vfemcj2m6824X5xahFYmeliEqCdCqKm83TQ4Bs/19g
94w5kNa5UdTqThcK8bvB2ypJJLkfjY3HQC2SnsSYmagPYm6RfenUN5Rk3Mrvm0Jf
f6ahERQ0y/rshcEq6dLW+0eUSX/eePPlizUiTqaxcOSLFE/KvCH8YFiEU6sBlP3s
bWcNl8UGEhdbetRDPN7d35qv3iSzM7k7/XNNu6gagNR0qDSDJaDYUxBMzwIrs793
Y9OBz15qkK8cs+/IS0H9aQ2czvFbXIPD1HdDIxKPAZ9/1YuED0F5tvSrQ0L2UNG7
gXh3ubDln2q5aM+llCKexR3LAhPy2fFVCSmlUtu1Yc+Bd2zuOa5ggD3TcXJXjFEc
bVRZgWTo+vg/dR5oNxm3Pd4d0ZZMg/PAmWrT1S98OyFEKwXZbwb0ThQMQiMaFYHY
+b8EL9N7NGOb8alCIdx5+c32qJpVOEajjB2I/POJD1JKQmoDPU7hnJxeZ/1DFGRN
u4rJa5NGXeL4uuypt+zD0wz/PSjwkc/hygCUizm6xbc5LQtPA9Hp7oSDHFoBt/wT
QNsFa9rFTS1QPEJsRCgxdvRN/poqAjVx3crQPlG31UiBUp8mqrKoAXvujvuhrtG3
+hvCPlZCXcoRaSIQcBrozEP2d/G9zRmthriBqPJ5269q2WD7nAg8Gwq9HpPBssjW
Vrsdsb5Fu26Zloud6RMIwbNHeTUewDhLEN9HiS20DARhBNq156ykgg7wYAR7KNJv
LRcUFWkqA3KF67I9jUy+1djoPB6n7Ty7SOU3DnxN3y92Gc55N8LOlvTtUf795/WE
FlYhxBn5eL9kQ6t67f3pDTZSRDgxsovWYucxjVcsX2dw/SyE/rGWbX+AvfB2s2ry
kKWk3JvXGAR097Z7bBLgtxbKm4ltqMEdkpr+KQkiXk7xI5KkxhSojyZdkxFhlPxs
s5SXlft2bBC8+bLQVnjF9HaamNP6MmI0gC8GTXjAVM7nwgrjJnycIQSm1nvvgoZG
Wxts+gEJMfA/7TSPeSCufrNTCIHlVbytxhnO8zdSQdi5v6hHXw9yq6u1J8FJwMav
U/KMUXBZIHCCo24BOQjf0URABRAhOBZ5WVe0KxmvUEnxiXhKJS8wXKyURmpSRjkm
e7z0c0ccvazH8seq+H0gjPqbpiywqUMc8Ol/11GG+LlLfIFdSj6Pi9Xk4Iq1pPWg
wfojDMyunQaNVRbgp55EmZCAh5bBomOh7ADFd7k08yPoznNwi+y8f7DcCKoXqK5S
xe7JpTUMMYOH982IUsI84eS9cS2fQq161MjT7SDdhiFVczOXzelteipum81vffoa
iyYyfGZVlxdi46nGs3Uh/rgMsrn5sKtGcop14PvW54sxZ5/c/mObuUpc4Mm8oI4W
47mvQOg6OkKhxXQeWMey8G+bXV6twMmviL3E5XX32BjxATVXS1w/M81m/a+N9iU1
BIBMWgRCbyI6EZRLNvHqAgiJLXUnzCoka5ib073y6LPxpTVadT+dOjV/EKS7DmS+
GO5a4Zc26BD4a68S/oXKivy4hey5D4dfOQviVV05LgnLfHComu+CLB7bySCNnyTQ
/gXpxxVJzW4l/d10rqmZVt9AWHNO88e6caoLwar4SvJuTG0RjlIYOGIl40/nbXu2
6citfo6V1TNADOUtanj8yFq6SwMtH0cE0r99y38YP7/WDMyb5M9R+hX7jiD8RMyD
4vfjCOvjVYLqWSGxkkRTI2Svi/nUdp48rTkw4UuEg2pt7Kd4jjzgJQ/zj7qJiBrX
f/eeSpeMEO3gzLLogj0rCXCxwFfsJoD74Zpq+o8MXmPY7mileP9WEBoRBYBiHC7t
MjrAg6NDJ7V1zLf6eMcgL7sRwiF+yV+Srk4PtH7HgyRfDXZEDF7c0qQBQgb5arQn
PcE+55HW4VsTq2yah8FC+mV9rsMz7T3nlICHFOmyHbrsYMfQmtYzXLmRpFBQX0kV
K9T5M5OLA1Yun5a7wgprBe5vMXaoNhTnA6vdmabZDUtQN2KWUnmUamXs9Y8ZsXcg
Ylq8Ixj3qpjuX6xyabMifH5ajuMjxSIh6NzFOHTv+kEmWuzpPH0DWi/Q5jFSb/O/
csZw+FXLsPR1JBHQ4LsrAue+83YSrSn86zP4h2yXtGQUn5/jDN0nLQ9lCwB/5j83
2W/YFjthFIaT2cT9r224hPBpkR/w15//RjCZPWMb6Vf95VcjjqKdIdwRgPkAhVAn
WXwN1jFVNr20F/0U4LrG2FM1711TyCd61uOe+U4mzHp3CJBr/ug63QqVchk7m+J4
hOkyaEWOyGyOtX3bqnlHE+2RsjHmA1KS0Uw+lJFdQIogatwbM0Er2fp8a37E9RZ/
vKjVE22b76KNd6jtfqAM0P2P97ApCFnQDb00bUL22nrPmOBr6Ne+c37EvTKPzFt+
XPTw0dxur4iqWfIoINlj2kiV4Hca+8+j8ye7DQzfSoXpJvj2DhQV6BvZC9MWu09J
LQkNihRZWk+9Rn8wb8m/rRZNsuZtxuZUMjVAajU21h3s8GQy/mkJBQicaUs+Wxn+
TSvl1Zvae6mA37EgDBOBS4+IaTCWVbsdVzqz7PvcMQzvFFlcLZ2W8sGNQ2M7gx0Y
k0v3ClAPD3ptMtrsOEhwF5cvy33Y00nKi3INxv7Ue3KwuJXecHwdVLrLjqlKJby5
wTKEHmvVFFzRQlpwD6XcAYLXgb+BTLdLeo1F0LDR5Vs/HpNAUFOS0ws1RWntDxUO
BPMfAjXvRQE7iJ2GcwSkVgvDmEdlfU3TNT1SnJjgcVyPVP7WjaGjYGvIfKx6O29l
mXMirkG4jBDSZXEUMNZn7JjIOf68rsGXyignMV/8amJTE2MF93Fcmi+4EesSgz4k
x9R0OCE4ndpEpEhOY6xKnXkl0TG5XZNNrlHcc8BsrR4dzSF7UBWeIKb5LGySsKM6
uUvViQ4jGTDI/ybG45vN4GGENYWTeRlkHgJWVWT5Cc1tr/zIUJnvEbHWi3LGJcVq
G8TLg7b582wWx5fZkIKzQR0QBQ26gTrgg5xvsauE6PAKaVLSAu/otGdCstLEl1wB
U3qp57bRp1lV3jP5vIf1GcxXve61dseFcimuivPzgFHBidrgYEsHWFNsZdqt0/Tw
G8mVWYcKyWXgVDE1IW7AzKdsLsL29UouMORxZM8qS0rqS1RovqMdtHrulBVH5Vv3
MOd4E6dvZ38ZjNQBfWC2IVN0qxbiuM6LoXvSgvOy+qyKSv/217YAKa6iLPmD6iFD
ILEgpBuS24yQM7SlDxyC6LRDs1NyGACJ6CVE5RfgbstJubal9PxxLfDW4aUVuRYG
bHiDsVgTgmpEmzw4wXKdyNl3YA3ovMcLDbBczgQLqBgfiXHBUMfc629m/Vb/YIo8
vyKGoRkqAf1uFWG0S8oqbU5YhJMeRuexjtyfHU5+DORHnbL2ubtC3k8Ta+tvJlQJ
Cm9yngGaegh6JQF+PLEFSkbbl2hNSGo6MhZI3RzlH8p5pjvWfd0MRcAmTy2pSWLa
D7V5+ejlUIiulbaDokRQdXlxST4vxznsJBObjB4K1w3eqR4kns72nWlGNG4KnQH8
4XwxiiN3NhYCOuohlqPYr9+W1g09BzD5vPElTAGpAZGtY+05KUzLIpXj79d4y/EM
xTXVqNz5lTamnVRMX00MQCWdo+1ZhKkurxJj5W44BGUOVKJuvaxWw4t503ck5kbv
+JKSpsF0Cl0lh8PyuK2BBDynguWes0ol4F15UjZU0seI38p35Gk6R0maVKcYhU+h
weT1/5YrOLawKi9Mym+7dkIggRNJ4Qzfcxu8xst0H8E3mH7uxJMExXhsl9/xutu/
6cehpNLjChaK5jUYTA3amlNz4QtqCA6T6GWEwngkwI4GshQ0V6uHh+D0MpREnNg7
s5b7ACAmxFVezwdx9LnUHsq9dD1cZDAkJjkfJ0pqX7TfBIpV5oVw6HmWg2VRMq8w
aao0lJ5cFdF98hRY2MkW0BrH6DEvg1vLwzfHEVH8i4XBwswBXvXmnnm2zuM0kR2J
agk82txBOTWnECL3L1pnxNWJa1yActjC+LXtL8vuUHoACMKx8twRrUfWqRKkRnPB
PoTesWLJGSYgeiqqNOe1bcZGzUJbPGuaSWHa+xSkrl78QXF2ijcYUV9gPjLTH7AE
tIimLSzbB2T76QeTvuFZPH/72YeokENEMDBw5dNIeFmIVKVZ+CNqnVPZQA93b1Ox
/qWVoroGkmF4mI3+edmLsfNiOY2ItDRYliBEXobV/KJYLI3XjF5z1xPf1NkxcOvn
hHZImzW22jWEghxMDW3DIClqe1onuo26zJsnjSLpfdYWRmHuq2Mr4Cn6XbvhdQaX
luzwAD9PhjviPR6tDHfo1nRA0TLh1OnpnGSMJL+Y0R2e0cwJv5xuDomqjl9WXngg
T6QqzNH4L9GCbrd5FfJlTtUXOcxtnEANTZ/TjtaBpRcYA2SmLt5Bx2e3raQab7ri
1JDk342NPfY3PS9CDCi0us/CdbgoJt4frKKyitycreL/3x81jE+gwqIRtbKtC1ST
CSHrdwSLskDSAFLS443s8d1Qgsy3qHBs/u7Vdnt71kGGryQIqy1rckTceiOpjSop
yUOrJKuzIw3hzYgdw7922RGPBPYGoT38x0t+dnuKat2L+zskoJhdwt2MfNBxaR/Y
fi2locoo6Q4T7tBb3kpqj5Eg9yeDY5jWWNhwt/EaBiDzJjvm8sD5gycDA4VKLbAZ
7EIIw0xeulpZgkOb+ZyhtPOqMnzNNyMupjukG04ujSicWYkI0bM35+1OKCxHi71w
isVa7gAiemLPva1n+7CEKBQ05kYU0eG13ZecMy2Yslcsoml0ghMZRpZzhGVUivWr
R/hx6PlGh2aIE8UZaZg/q6GxPs40bVrJgFjb2S2Bo4ag6T/kzDSgvU4YeZsW2fDB
BpbShWXc6USpgv6Op2s1JYGil69SOkFOojYwD/B/CYF20lwvcUhYmeH1j8+py0DF
3ke6w7T0fZrD4ef6ZdOv3KqgOAK7Stnmw8rEQD5TG29PI7t0hs07+4VjHpy+tz+T
B0LJiVjwEDRam1akeezRrcvk+iJM5yy3wXha4vHLpgJdjYHqG4zDeny42uJO0U5P
uiYye4zpV5hsaCCjkIdQ1VHBEtEr7N4f5cY7pyReD1DmMrXsHAMU0QMbmD/dllUS
zeR5dLWnbv1RMvIihfvW7Macx6ESAfgUPE1OfWFl1YEO6OPs35kMehMGAsfnSM9T
Syw7s3U3kobj5dx7CgFRRyWuFwcm6RVpMSW2EMRte8R8hhM8rYQAhvr0yqdI79ER
i4LmZQIIsKZA8kYmHxp5gm5AVvgFRXDtE+v+6uPtURQwLvNaCbkowKx0PA+UYvf4
uK2c1BjLJzIwgQ6OmjPXbL1Fjxg9RgEHuEahTafkKMTSInR+ofczqvIH5V8GbiUv
1bfYTlqkMTu/QmoLsVY13BZ4P/e8b4h66wQ68ezSkcdH2kXCOYbbpoJyqMI6faUH
UvUrsV9pQTZZNdyTIDowTqJE+shszP47xdh7xfYfIOZS6L8fRcqeUrYbaYsGTZxL
wnxlPRxJbgTmZjmAqR+gZWdA7AoUeawgH40jhLWUasl28Tj+Lh7sKuC6m+mZaH4Z
76+atmMXzExqKbuBbtQJMv3Fa03oXEC3h1NV8PX8+bTuJ/Mp1LKl1elTfmdX2WTD
nXtgB5jajEyoZq+Xp4LmHuDwODzSPU/3IDGKbwaHldNcC19O4juTKNNc6VEvJB7S
xc42ROwwaOY1DTasaynbcvumdtqZLKdju8NO4VZJWsfYLJMzazhBKs5wVLykehs9
oKKP+lEknAUmoRqYcDl9H1nDxJ4SnlSuc+g6sVJuhotquk0LwqqNUVW97XjteBdg
yq544k3cpTwRuzayblupW7/24eoEzTfbkYzUIRDjijiRqqLuC33ier3RPh6Y8DSF
93myLNS6CvumnM+tXeQ7rM8N+E9xPBch3x7V6Qh55opOP0hvTqWnZAjmeX2qZXmz
pcmoKsgT61lLD9ySh1lb+dwxZUEDFUSthFlpFP+aDgmTE2H4HR+sCieg5wjT1nzt
jNxCHViRICBiBkc4LeUKWsV3b+hG+HdqpDUQqm0MkC83BZVX+WqL86uIAif0FPuV
QtqrmeFU9400F7DWsryXGbsgBWpQvsowgo4pQUhxd4ZwMnmMjbqT7g6wGoJvhDCY
jKCby4ifdwuHfahY9JaAugNfC/WtsvzS+2cUw+1rHOeXY7sV9WIR8qe+dOJr8Yky
SfiT1IkEk9vnrx+GEtPIFnLw5eb5pt8UmT4OZLKJSR658zgNLNgVu82HVgqb0Yhe
rywcqTGrhSf1X8w0oGthQG16dJAtWoMlFggxpeJJi7ebQ1rgo1nQOQ5m89cX31xS
lK/EE0EcKCn9VcStm+aq4JwVEFIHyBOhPKP/1umkYhsNfkQwtAIWwWOV7b4eAWBA
UvYRZUx4iCQrCGBNNJ4YqZc5bPBj/4TNX4DfyI1K2jeiYIyr4bLn5elx2c7NQ2cb
lpb/OvzgQ47cFyu2zSqnU+CdjM5c7Np0P/ba0ru3z6BW/F7/xPrvgTp6SuGiRy1v
PLMVgPmBgbX0pXcechjLP6YT+s0F+f66TfXhb9M+W6thnfLaYJspYZIZPA4EAUyW
gGKgZryCTgtbKqisxKwMKNItRQLdnI6vYyrSxvOUyRLBw9a0fMrzaKE2MaGpYkH5
ih5KR1bCWRIthbu4jXYWldYhkY7O/XAzufXaDUXkaX8uUzR2L1Ze7kGu+SZyOEEy
kX0H7eL39AnjNuJfuhQSq8pc24FC6dhTSEmYL++ADYY2XtgjwJHICVLpfhGBHExl
XTjpUxM8cIgkqDQRyM82z14cEvUYZLI1P84/v4M5445tzncvQj8WgX7iGSnMbRdw
smA9kakxeUFe0wEI0zcYLfG+TckVbGbjzmufMYqfHlNttx79bVUKX/wy/fpGQ02O
AQQ7AINu2UWhMwYMr8bYb1d4jBowPihvXBFDosvX4egqdHIlmyGmYChoGIE3tjsA
zgRliJE08kaZkHWaRB0bFVVwfvGzitjO5o3ZbabZKlrOo8J1kvW7+tugwvH2qP15
QbwD4u9KKsAP5MdptOpQgqJkyd6SCA3GhcMmsuEia/lAR4050fjqGCtPBvXSA7R1
Xwb0sfKw5jiChf7EhdPmCdeLmpTWDapxYRUh8pRJDPNWOf96gkysmsHdSgH9NCJD
hfaV91ReA341QMG2Q0Sw6x84aEO5l69/gRs+YjDdwkUgcotG4TRKl0KYTspcwqE5
UjE2c1R0ZezrMy8ybV+EbkeHAzETG0oVHih3k9oVfeM84K9aRDnppXwPp2vwQwSi
J7oP52KfCt+w12lAqgIxMaURkwhnd9NSFJ30uMvsyXT0uztSdCUY4UeUzHTYGG1r
ug38WoTHiNPIsKLhWizIMn1L7g7c3NYjMKpaQF+B3kGntPqQw0EQ1XpvT7CzHwb6
X5EOf0wX81mVfH3XATs/k83NcGZ+W/AkKo3KwIeqp9Mr5XRjKVPHF52fRTdNbq0c
PLud6DztD5HdllojTJXgStq1sYO1XVI4oDj5FyFWSUF9K7tIkIrS9YyEe1euJOIH
q2kIGmVMiVCQCoOh8YalUg7hKOsxwTxVAHqLZOd1qsUKChu59tHkLmfo+09EX8rv
8I8sCjSQXuUKj7iFl5EuotVs9O5I2D5HhEwcRR/zG61Z8f7rY2Y6IV5NsYAUH260
6P9ZliJNybCz94VY9+r2A5ldYCExIFd2nLKcQ3Kvnmz3+wMgjv0bDMkLW8zL1eEG
ygKW1PWVxKytd6Fx3siVIceaYMTc9p436DtDBpggdV6+t5twwwbWC63+ofrxV6nt
DkRQZTeQDjuarpmQGZIs2HR6cx9LFOZJwNFIRRKRZxHWgwJ2yuyUYHW1CxqTnLiJ
qEZCQ7d6T1Ww35JFKCoKB48QX0G5S4bY4HDwjbDZ59uHI8MHbcACy2GEtQx6+gk7
XFVRph1/nbNhPC8z0kFXJp5h8FOEZqyOgx4usw3XLNetbzR+/OVSr5hR+dAWcdGh
gemoNjU+HWmPMOf7gHBnwmI4K58EOBXpboABOJhsZ3qg5faEaMGk1mYliAJ+YGoG
JJsdkyFNS+zmdurGma/Uu3wDLXcoJhrNQI65U3sF7JSMxQO623ITj2tSucVhdksb
8WTqUvivgb2Aob17ktwAaOa9k0w9k3R+zpgRPEBzYa0EYwwPU6vzHlgkWDCqPaPU
MXpPMzl7eNdSSZU9/gucTs86l+zwAVf060cy0nkaIUzdrIcWQ0omBmM+HpsWbHlI
Z1d3Ga0IK8sQasLFOO1NQUCNrjAZR01ygUp+UKzDHwlNKf6ZZn1wmw03bfbiJOR/
W2mYX0NUTfqOwQT8r8eNChmBMHBw9ox4GHAXA48+tHs6VHNp26JNY8XSACg4TDHB
xTYUA9UYfSFbKTlc/ttUHWVC4/fyEvt5Yw/oDRgddU2ESwfh39O7pHzvndguTenr
vFiHZashwHCjeiLoVGFocRCm1uLWzAg1vrcj4CMzugkuK6mgAbTLtc+jfdtVnTcU
X5ePtP4GyH8GhgD2v05kMTsx72Wyn5tKWCqpliRcU0IdETo45fchjo7vdhIZfvJn
Qe68bVf4Oyx0aRg3o9EbHwxJayH0prTQ4rV7y1TeB6xOdPuI69kmt06t5pPyUhFH
Odfq3Xd4DMqRIi558zzlSTRzmDwruILit/Y8biWxdsUgNwsGNIbrzE3O2RiDJAWX
/YLXCPK1LcBYshu9YO31C1HJoXDdI7lBEmJKKRjjBRqxvFfUq/wN2t13HsSO7b9B
KpHRWaSBZ7R656r3/CDZI06ssehTWiCdx5y8l7+WKwtTHcFM1K1bYzLXfz3/g4zT
E9jgOUTu6FivOKMyzHCv0uTb0nPSlHFTtqcjH/nbeKx0apxgBrzsk8HLz3ABPR3b
Gr3IYpBsxQA7MCQWzhwRttBQVxJh8/gVTmA4A2Etv6R7xda6ma2I+NUd8yXAxKgt
AA+31FEvJrRV1Li6goUuP3FGS/ANfZ55wl64gUSp+/mmY3K0I0LNUnaU14oHFigX
rkRFVFg/41AwweNoruPA18eUyu+HiAoicNsEDMUULjtCR8t9ZEOFqurkvAdrOW1M
5qypGESxW4U4ag1ThjxB7bm8/mAOjJSC3x/2BvgqyvstdP4/blvKyW+lkthZ9lru
lGSyYQfXulRxKmJPZ3fczSqQ7BKFE1jH4z0V3e7wOSK1sxI6urMa9x6f1QPg4MBh
9ZFzT+o1NOtWhYz6FGGIWzWxC8F+jQeAUue+lXN+DcobXVkma2gDn1ZXGg0mtSRn
2OpAMcRcUERcUQREAQ4svqtBpeSukObIT5Lxu0KjXkvnDHH1zbH6saLCPPahkwvR
ch/HZS62zYpDAyEH8gveR+Igkvdc+vY11czI16eyNJimAX787NIPntYBjTAcpdxW
/KF53BLJvy5MbLJEoIXR514GV/i+zbaGzs8ktsuy36EZ9aR2N5NWLziU/c8VO0o7
USSpCERP3KotiB9oZJATqlfAk0dgcaGgFUNYhvNQyOXawxG/ylNOFYHiZfUAQZii
vZxBqtRInY76IUMACUlzowFLJXddewzIgQNoh86VxNlM7I09AaZeuDNwDlXR2ey1
Ld++u+kUuodwQWtdYTT6zUXDV+5VrFTBMEXeDE2dUWz9lucM1uncRxxwWCu7DXbK
x1cwtfnvwEjP/4fZKmwKUvLUx/PN0g0842jVtkFqCrX0sSslykxER1/JDIHuday6
kkNEY8O3DLILBfklSw/zjD0KrkCQPbv24rxlpRhD+Ki2GH98KpkT7Ei2ccpiZIQC
d4T9TYqpFabzpuDi+YImSbsJ01zRJ1a1qTXQwMImqBNnZniwwaIhPk47N1yq/Ph6
ZthNXirSFPBLkY1xy0U2Zv4NyDOMIpi6Qj0bRsaSTTk8da40s7+NH44eCj3GMbQ6
QSY3tDMqILntdSYbP+6/QjqzeJGd90rq3Vq5bM7zO7hRF/0jG3zLjfttGHO/zi6G
O9O9VwKP7SVxYjGEHnlsXPeRrpG+aD9tEW1ZVJi8hDt1TutQyfVWwXkrvCS6tatO
RvCTxRP4BXfJifq8cGceHS+kQ0Y5EjsUGjCAwQa9zoWLMZ5Fr97ybXUkm1zrfW9j
ihmKETv6hZ5i//BzgswFWnaptq4cMh3m5ZBBrkb+OfMDH6/BNtjceg4694G1xTA3
QUXKZtR+pbDZEblpP+9wOl+S+U9AfF28dnN1xNiSO6YEnLLZEoRK+m+lOasA5iXR
paKH3F4m2p5USl53aClDh7rimMZvVH34yAE8bsZfVV/kQn4bL9B3ryXNCJBOalkC
9mvchQ3mlPoHZbOazLP9q/RZUHQuJWxSpcOyogNM3zkA5JiXYpzRFM8ds95R2/Gf
iqnxqvbn+8QD8kM8wuP14D99LUjgfZBttkZ1FSDEF6T/TfgcDD2eIuoq1fDSwTEC
eZsS5WzGQFrRNpSuML0O5UdKy0uNCadJomZyF5Y/h+DstRsWQA4OGVAG+W3F/q4G
73vpiaOL5Cs/7grTdcwx1Toyn8oVoEsbTaRD1zaDhuVWNKmliY4jV8Wz3XZmi6YQ
Aa9My6EeBpISBmkXl2gRCdSQYqphU64mixbm94ODo+oeVtGfPuYzJ09CypMKh7eE
i2PJWbFzWeNMy12QM0F0zxEWtCcF+5mPhfYnhk/QHQS+Pbz7ZPdLmKnTANJnlO9t
t7pCV01fxAeycsZNsfcvn0C4rzHECIegcx/xx+yrc7N/sjXNwyWKeOIVJy/qwgFE
6aJNKp4adur+HDfMAKVItVuWqvj5T79Pohpi7IfOj0GKdZon217djwn0JTxVihA4
jLZDgD5qogNh1rARgfWFcKH9BNgnSC/+djdjwws1owKY4LoSJVF8kL69ii9fbQev
mpiMVl6ySx3o8HtrgDmnfTRVXYuQ3irhTy+0ST7Ry6dIsRm2qiMwQ2j9hjsDT0Pk
sgRHNWdazeADOkAjOtnb5hZf1AY04QUNZeCASCtLZxHvGZ7tIXMwfQf/kfyyzaqj
AcLfGL+deIJXmnjsGv+htC1e/wEfcy8Iu7ZmKIOpYnQ1wBaJcdzAu0oiYQy4j/1L
emz818OK3c05bmZCDHAOR9TfrohlDuKzMAQlItQhC2l2KOjbaZpNb3eW6ml4qb6y
YUtOKKf9vWQttXHYDOqBSLTZroe5nlS9aEdf5BfmWvhJMT58Q0PNPDPvvcgEU3rT
6vufsrRuUlUw2b1eeg7qmr6w3oJP3ifntERbuFOqoMbC8nvjifzgxWJZ3spuVzKT
pWSxxr+rMOehxlHcSw6OR8WXI4JUlz+FkTTal4+mTxKsQQZkTd05h6dbkI/AR8Us
c2MREUOOkaK6Xoqb1bJMC362s4wpKd515HDfEWXfjAzZKl0GipG/ZTT+E+tTZELk
l2EyhwOc0Se1STzG8yZM1HkDosSYdXnFvFCsulCYcGjfSKH2ACsNVYmHwV5QcolC
ZO4T84uj9G6hkIGafrek8HdiRAWY2nyqN4q+AZLMpNQa9FzXRXlfvHJKaiRaci5A
ZnxVv/+BD0H6/t3H3HGLVcCxugeFKyRt3AxROXlkFvWSgPiQ1q/pzs4ACIWyBfnE
dNh5TTXN0S6BW2JB7w41g8Zusf/u5ojmlWYe9pH9HKHABfFwzh4YM1gNrNDBmv2W
wakbGU6eHMdB+jFU9THr0hg14pLetykHl23+BSNRLAhpAANEOdcF5+jEptNopthq
iPoMHr88caDpB4mOnGILN8DSd+acnogAZG79FPCGX5/ODLpki77HxarYSPQInqWE
WLB0WAvM4HzhwsoAinvT0NxACKTPMG9ipMDzxBIzLLadxMpVLhh82ejit4Ng3VaK
WuqzE9xNxkODcxQJ5NeNNNY0sOna4Xw+d6i5LgeygugcysVsHEOlziEvqo2PEiQP
R7ZWGlbgn+WBw+4GqmQzjjsTqNQTe81Bp95IPZCBJSE7s7Kb0AgChK+SB7/H8/bj
oTrZDyzTjlr7KVmhAz7OditgBG8bETugWxYlQLMR44k8tWj9YQRPnEOACm7//PQC
mFecI06KiG0razMxxM5I+YUHQjtaAttliQ/kuOFjUw7VA/X2mJqHq82YcGAuaPUk
WhrVqln2dkSSU5Qr4DYgfxEYJcuU193WZMvogwx4h5zLNmS3ekvmob/16f8kHqx2
vMjCbfPQ8KsxrWXNjSGi+BZvvMPgynDQDNMIK5hezAP8dMC1W3Rhk06siUPPaXGC
zU4adWrHCuU2G/SBATRJyhmgowETzIzhc4WmRdp96R6jdVCq52RgyemIPmrpnsVJ
55wCPrfj1IBE4ILmxpHttf1Pl5OuMvjTWFcLVSqHzTEzkN84uR//Yx3Rss/Q/7dA
x5OM015+TTDFvy8cDmx5trcO6c1z+C70Wh5/0RHgPpBsHIrUxYEflL62MIvRHsKo
d8mi3c+ogArdZttQonHTpOpGy4y558bEU9wwYwkwTNKxLgV1qHyCHYkEFQTQHVad
B23rJzZjWqOtadwP1o41Ijq5VCJiOEFtXmn5HUg56gddvwFsYZnZXfYffRnZvdmy
nnTXVdsavkXvmc5tyk7whECG8WBojbX+Hy95F9rL0MUTGns1SpkjV2h3iv4ha2bs
0b6ux1ugFBNJUYc/mUnfhfVd1aYIcqZ74Ow9BhieExh6CUBTN76c6NlY/0BRxwuE
BPXMdkMGEAXj1sDOZa+Lstx4SMc+7neFCJxQDer29Eq5lJIatELtQB083yYWAz6J
KLIzdo8YdL14acKdqCVrT0i/GsyinKttIP8VMdvJzGnXqTI8SYf1IvSHvgznXJ6c
rAXiPKujpnh/o/auN2Guv/+fcRlSyPZP9ZARPhOnjIx2x1LtJNaD7z3SO0mRVI4+
iG+fVwfWXE/BJ+xuoyaYPBuvK0avzPinhhpksLZ6zas4T9/tQsSYtK5DYJGtH1pw
TPzR7YVWzSYHnGRoTwt8sg1PodoMqMCMNUjRhls/XmDo0FHgrkzbNd5jYk+Bwgj9
o/N6ZG2rrU0siunVnBqRSF7AU3ZKco68U2boBpKjglUDJUJYZcwpnHKm8JJ+J0vX
WS2j24N3OJIKY9hw6G+5bpt1W0wxDl7tzovnR7wzDeczOeRWRDlJAfJBd1mAJZhK
YzCReqiqZ1K7W+ZehCV1ZgzKGOW77rTb/Rp/ATFKb0MJAeuV4Iu0aQ3rNLGcrNhV
AVQ5gyWOZ5RhvE6/zOq13n8Omp137vi1okw64rfMEIVrtOwRMXJHY7mnLlmEtdQf
8t3SfsVMVSepfKKSLCHO147uhx8ltZOpkCzO+52sT3AUB4Pi9Apnm95Lsok+O/w6
pHFIBW51uuF7krLWEHkV1iFFUk5T1fTrF20RUL70/dNXTyXk9HoPT6tzVHTIDyfG
x2/NrXz5n4fB7WwWbSteTyXTQF2ozGUT7/JOKFriP8fc1KGP4Bwzmf3fTI8wOe2h
bdSguig+utT6bS0/OmGMiOCDRII6pD1cQAmPfp/xlw3+6N+5OoM7d5gQNHyR6t0I
mdLcPWxAla5dvSRVM1lt13ZE6YXUqphaNbyZ8THIp8QMhe4BWJEcEOAIlROWgDc6
JCItrS6ZMefla7yquRKQUVoLe+kDYjPx0f7ZKCdfVJd/4f0dSyzFIQt2wnedDh69
TS+QxsSXq7gfWB5YCM5JfNgkvg2kZXxnG1YewAVRRe2t516Ytom8pyHG6Kt+D7iD
a3Bo/9tO+13HIultZCx+vd8Wf9mBPeDZ2B0LyMu32M4CnAnn+zKf4yU8rJf7vaIo
WSYa3j1VarkP949WFB338un7UmfsW1oSxLsKTjibgXD/WlxecqvEnS/Mb34W25EU
VyYMfljWms/52Spdurz1jdZAwhm32hR0ubH4hzfXhXEohhN04PsB4e+yB3USkg4g
RixxXMkvZEivTuRyGQ3b4yVXdQlUUAcU/yQoTLk67RMEPBv9K3ruT0Q8jsok09EI
LPseOQK4m0fBJzpbTR/Atv+dClxOMpGFLFx/jCFgP2G6tYZ2i8Yh7l/4rU8UhdNF
/EokhRxkQngr/QKSQ9q7eSePWTQuKpnMjTEoiO6z1smXCChDmd0oSYrOefLBDI2g
JGcnJxyia/bJ3+G5JIDBHzmq+lDceHeYy8kdpRB5fZY1+iz10y6lZ3So2QR1/ylE
tscgLBLkEhQ6fTzH+4M2mAsSaNFu2gwD4cRlnBO+CvmuCSpZtMn7eme87SLpTLAL
LGKo/zDpeU/4j+1G24tuORLdfmItQ9qWBcqyAv94k6oUQSuzlOq1g1FUQ8QT9EKn
5i9Yl/IF3HW1YgLsrf7q0EG9UYGZJSXcIMFdGFI+Uw+BwY4bXI1lt3LIBqq7lCIk
rRuGL5LDAodEfL02NdSj6u4Y8rQNvp6P5+DDJJWbaaf4hiLlaBA5oU3YUxm2fYmr
riQWL2fBWGWiE1ZYjhYsBqHURIhrYo/ATXCWc7PgZPVHQJOJvlF2iIGOYY1q7UTY
hxkzD6lc2/o5dhgQWkVvRZ+HIoC4NRalVMErJgA50q8j0coo+I9L+evk2yBUzqTP
XfmSN+cirZtH3hk4YUFy/cwlFEPKZgikKhqo5KHVbg8H8slVpEWxKYIFdH3mOojI
Nq7EMMR0zomzVrurzj6bJJa7hYzzyfpdgMp1HjIYgSw8msyTIvfKVMqXIeHCDxqH
6PDIcLwWl2rO+7cV2/GJzlgMxwiqQ0TowBsHIcMJS/F5OqJfa/bZPvglJfKwqydf
wnNdR6WgFa8C7MjrRHuASa1H4OuT4lqssAOEvDHj49uW4PahEK5GGADeCCa8t6DV
EinP2GZxXxXCiSR5tr3Mh2NAP5tLCLq9OSrrpVjo42FBYPQMvFSX8KPLcOG68wad
K3xhd8N7YBB6vZapl3119dJOKLfP8SOBsdZYCjgwE3QfNagOATnHnZMPk4OCbEB1
3WsgeJbB1q51byMXx9G5XXM4TyhonAHmAft0DlJrfHJWuH2RYVtZGJS2fTPiIwzD
PRc7kGanNZr5q+adP2jns0p0dEFpmDl/QpYeGQY0D7dLsG6+BwhsPl/8bSfGYbIn
DB7Jw0IkNqnAvra2fYQpTBzP4Q81tUkvaz/+gXmH+ondaGdXLxH8teqiVF9VbZjC
ysu9knVndEOFb9u8VGxx3nu9WeQ6qssJxUVXSlMTL4GQzTZv6JqslaaB63EM47yW
Mby8TbSg3IEiVqUNB5IaHvGFWAlbqSI3bl/I97CaFOPI0Lp7EfEFmCG7W2zC+mp1
DAefLm2KLS6svhCtRuveL7oqc4h4+jYoAuSwEzobuH5sm2kbDq1PpyKCA330oFp/
885vzCEsBPaZAFhPyajAJrzEGiNBQZn/555C6hKD5Fi5X575tZ9U1q8iDZzPRTEI
Qm/zJv/pJZm4SDn1lzBSX9ukGToytLbvoulx2uTUxE2poAsycGuZjrEAdXyutmko
KreD6tYqmvOVOqWTB48kvLf/q5uHSZe1VpCQ5EyBFBB3qwJannNdcVC60YHUer9X
S9Iiq+MPk2GDHvV8YMyeEW6AmVmd6iOrLMXRbQQVVAOpktnqEOCkMGPGXJUZ4otO
tY1MoeNG+r5gBnBzOid98Tn34LDNNbE/ohpLAkkzJ6etOLIibczlh7d3pUjsreVd
Po5RcJBgsbGSaQGeZh4lVO2NJRfmJReEtxWLmdJZXI4RKyLl7tdpqejviGtr9M9J
hepGMXzC2VZdCsHyjFNIXSWo/dAuCvinmFnTat062Rvxf16tT7/9ZCzGsocJlXtG
Ojx/E4JpZSjZEO9JwKnsAcTKf/opATuvuodapXL/6N9Af0Jqh2ojiHsBXL06OeX3
HLxx13s/LY89+EhT2St/Wq6TndQGQcvtq1RGIAhYu4cKDj7EUeoozKXP0FdVVZOL
HKvFddglKSHKnbdduy+TIVB7EwPLjgcwV/Ot+5wHl7r8juKe9aFjX15/XMZp2YA3
rF8tdszyndkXdnNTI3zdXUM23WeujaZk62X/cjAEcq4+rtom1ZOeNMxzhzd+Rb6j
Mx57jg389LAmTJriP1YTgPhjEzQeY1ffRh5RBQBwJn2UanZEpliZ/klLyTYVS2W6
vxSZcIRfq47YEI20YNz2zcnHt+IcFhI+39cJPiyDP/fSCAvnZ3CPTL7kxotdvQPK
aIBUR8SOxaeVtAzfT9JAXNpTszEUciiQebG3NdgpcU6FW3uH+HADzz3lRnZtGLx0
bQK+DUSSuvV3vFP7DP3iChyMfCC8W/PkgSjmjo1dHjqTKeT4Km7ozkpHdrZ5Q3ql
urIkeyFR1nuJTwXsitmnKOAz5hmGomh30fUJXOSN6EGd+Wtv8HVnuXTDTDsFyksc
XHtOXwz1cXzuX44mqMlzG4GdZy+Rw4+/DeKcgZuNf8cRa5z63+HvbBK/yBBQh3KZ
y/t1xTWsVyIS2g3ZIT1ZAio+/Mx+8Xyj04NlyiYBlmeN5y9pz/CBekZdF09wXhu0
wAt02QoMzqAKoHXI8kB2SQ4/5pU6JNcH8/oO6I8mOoXC1J3lrGLO3WpLKNP3bWhZ
6rYiZzoTog+axMMzcAm6DiakAWcVJnC+GWqikFKUX3Zk4XnPFsb7NkW92HiFetXA
WlaRGQAivVWvV2A9yI5qDYTJs3niV8qsC5vPyGhKmB372UtswYgPKlhu4CI61Bi5
VPzCADn/ijUGNymmP2O/9ApfN+nqKD+m5NHpP2Hh0tXlO8mGjU7WhSM1uqfyAtB9
HxsdDW5G3E2le3l8kGUDFYxLCFX6mOXFHmGEhJW71cHUb94akgDad1iRBDi6u1tc
rGdmneM+YIt67eP7cWD1t2zZsGVvM0Wa2jJWa2LtA/p7KzhAbjjXFkghlkRdXL0q
2O/i1De2D7hwT6V8a2fqBOomzoKH51xV5nJRpCvv0aEiW2lhMtE2WxIpCDtI1N4w
+Ob8l3x2gd4Pina8IkuKbD1scrxNILQtPOrNmCTRk574DHLv9UarlOI0VJVr6cmd
sMfUllFHJwD8ILtyf2pQBdifPg8FiVv8nIflykYveD50WlPxXgNmsmrNSeAqZrCz
i42SL/K7dVnkRjWZ7m9NO/kkfus57QRat06JZafREt7/A+M2DcYCIASbzl32cHd+
uobGQRSWt6ICYRSQDXXD83jKLtM2i3VIdpiGaKrqVDkv+DjXq3fxAkygk8t7jieh
QbGMwdDXp/yy8Yjnawd8E7az5xHjPnRCrOHTKcTmajn5qMeHXDhO4LsZNFDEIfFU
Vo52YMVCLxTXBbMHIYjOEGzlw3ObXn+48eDJEQ6cBojHigWOyxDwbdqBVMxcVzpH
JU9E26W2rwW0Ce57VxFDb7XWc+C3xKTNlt9mUt0jvMZL+5FbCMBOiSOFfGn5pyUW
BxHmiRi/v8v4Q5FD0y/mAFzfppdZyp+VtYo9rEHg5OL9YVWOssql51Yza/XehS1t
TW34ZLI6VnnqUGneZEhe0tXXeDA1YP8C0l/OGGWosfFkEsnaGcA9/zV+npygtZCC
9BAnXlhyHfHzQCs81o3wPfyQu1L0Iv00g9HBD+M9h6hhhKeqAXtp571EnnujOC42
NZvx64qcfvGkoBQGrGrHGFXTulThhyk6OlsyFXhDUUwPv8BMl9E33SEQrklfmLki
T1jP9alcgLwaIz/XnpPot23Pxdz3/PIfN2RjFckWWG1ltkNIAf2ed9ESkHZRG6hk
BBZMyM/oAmRlW4sG7OtgzpVzWjbBkKO02A3Z9YOSpea4LNRf5i5hRVNU5OUDKBSO
GXdCcDxTYS4V/Ijx3pWlW/PusXdq6JFi9YUbBFjg04IQvq50flXUJmmcXBTIB9EH
FDf/bcTaU+FI0HF6NSlDqxTNGMeGduOY8ih1CRRYPZUjpDIisTUjv5Em6QA36rOE
LSKStTJv+R9ljDRrvZ3JoAalNiiYot1rW7Ps7gt74S/Pty0XusuGnlozd6AEIGLc
nAilYBduaQ6w69c/iUny4vJtTlZlzSashbqPL7eg20Cdu/Qvz3Ucg+LwNlr0zNgA
AWCKoF4Ntv4M/yX+ediF85xmelxxaJWGN5rF8fKxR2DdreBW39MVc3uo6VeGNDKl
DDhNPmWgx0rXyNlboXWKc2R642tzDrDBZZHLBsanL3SVUZY6a/DitEsqdLXOnCJ0
tBA7Ivqw9jz0UMKomRTxMzLaVenVmRynt9n17EFu5a7wiUwOmX9NF3XdH2XupNbU
JNrAmijRx3u3famtsobC8BTGEa0dVwPspGQ3RWvUZz5doGuhP/qih0KOpgaf9qad
efaGI4HZfUxJ//6JxaxJyMFgKinXrnFDdO4iFDES0EcGKJVLfatrRDZkA4ytm8N7
xI2qeGgnziuQiQe3W988/Doyr1y3xQLFV5Oabwn5tEBD5SzHhSu013B0B00Cva/1
o4py5mCXbniZ7GxjqbvFxBthtTpWfJ1ZnU/kIHJUn+T8LOI8i0xzjjLcik+oyydr
mwYMIixDe5ltWF9ew8I28pF82nr0NX2XG+uKLCLxeVPSiy6vqv750jcqZJChNjGS
IgZIUOIQiCgPMaO1Z24T5+f5ZGjAQe0i7pXLJQGpEYK0aV32iC4Fpm+ZonVaalNV
WAZLLbjnWjNX4sGl1DSr1yywlFyYFyBYg5IvNaxil3ODlW7lhGqtLqiqLesbTafH
z/t3+gyn5tWUPeMuwpi2ItNawBQWw1wHYTpia5jwmrWjOl07MzZsAQJaI9KcPOLd
cPS1POS8smavnNe3FnnWOwsB0OLy6PNh83Zsv08AKDLjaBm8g0aqtheeBmYz/E1k
JKQaxnl4AEsU87S6G+Gh5SjoZmgIs/MQzH6/b30S+P34aOhkrWFg8N/9iXyovJGq
RzKq3bJA/DecWk/KksaObwVRR/8+YxNuMkmrtrBqPcauaQrLNxdTiazunLHiGpIL
kXsljqREOyXLFQjdGwQsvOZZrQF+fWTNdpWeg2B7VNb03AuOuj5/Kt/cdKwCTfO5
iEkq9d1Etfl26HP3pdvahbVZ7rHxtc+fVuYMfZl//Ocg/RFv4Gz5LoLdo301wHPz
AxHhBepnRIngSZcLyUYPQrnZa7XbdFvYQ9gjzYs3UwrePqlS/+MlmAv5ztMR2+tY
NfHFXvuMlhnX7gwX2WhOvCJ+jaW9Wiu0fbja8XKHwxXsyKNcrWOqHdsHfgkwL4Tq
VuLB3W5v76+IoMhzJ8I60b+Thh9Jgvo3VOfZ/MdzW0SecZkrVJ0OfZL7eVEIe/Ec
ypz9GetUXIMbQr0fqDi8bfQjBl6FzLqbw1MVom06vnaSHdT+OUl8GqZFX4JgixmA
1XljT0SLZBCYZ3IrJC+I/pkJWMX5OJir/92ibCSYzaIKH6cONwwjxDsDOtkFd1F8
FOS5bG6JxNxtS9QgK6kAe5hATHgOvpTp8IJ/rtTvGjY7M+VOa/U2WKBLGLbSF00t
rUaM0b86EvMlyoc7mvEm3jDhIjDExKyEjOcJMb16qYxT95oRlorTOXJWEyoJ/6vk
guzWcXm/kOLbEMQccIbvpteyJaQetJobPzHBdrU1KWuh6hFVnk2EaRX8egiUsq1j
mA29r7sVElgVSAZXp8i3Z5A7U/pJTZdIlGNhqv8t5jwILgrFAkuo0wVgwVXjmoWl
1yz9XhyByz0OD4jAWlLj/wLT9MTVNfH4bq6wDAb3rzdSd6hN5dyXwpcM4xoobhy7
rnxM06GOLPWktPPrDzqu5uXu+w0o/6FcWPl8b5DSgLjZd237znMgQUB/MXTkP+3h
e14Q4bZQ7WWkcUFAocRXzjtBo7tL5NlKBad+6qz6Qhi+caztg1Vrm4m+pDsDCcRj
a37yKCkG0ci/E95O4q9awR4B2h+5VnlfEMG03Ef8PUbUOZ0rvPX0B7/yt7AQpKdI
eymdrUtlt9W+dG6xX686RVHPId2aw1r22AI77AJh4WV3iMxmaijrKll9xZKCxzMO
4Mjjwb0I6LwhICRlFmTlP+Imo/0TF3877zqpc4Za/YLSha3Mb8qh3iiNEcalWjsO
4szAHd3iOHFP+IIxnX/uRskjQ0x+DrVoHXXJEWbu59nTZZNz6cH1GVEr2cpsVI8d
2nThOADtUVim1LgkhFRkitc/CKkEzoK4mFRm16o0HTEg+8RjGbVkMGaL305ZxBP2
xe+h1QO+ZLzvkQM5eT2jBMTme3Mb0LdWilM/1wAlxFkY+AKenJznfP+j0ZAnJY3U
eo1dXfGDWrLonFQ4laxQNOt95X8y33OnsLuzU/aiY2IH13yLEOWPKttj+icdU5f5
Wa7OjUmq7uxFz0vjMBiXzL7k2rjJ2qfce6WuR7zpA5yWa6WeII5w+E6kUrBcJ7fX
pn0Z3Z3npDTf/XwIJxR7NxtBAttibEsOWW8mSi5FDC2kd9HDlvuGfzSzDGJHOy2X
E3R81rl2qruKY6+HT/6ysnjvddI8Cv5pynp9dcX5tyePpm5chWXERhrcJ3R/LtE7
fEElsdtH08rsHrrUtq0Duukh8L2M5Yqc6mbS96gMUl5hq2K1Y6POSyVApWpIyODo
uPFymRTMMybWRFYc7bvgnOfIc4KO9YtsmUoUdJXaGG0oOibkwbKDW+BfLYWTEjZf
7Fct5L/hXMcT2Ix9HCWLf5/42nHGjd8gdC1jHZrtC0G4bnzrc4m8cPQ+Sef3Pstk
6uq8ro0UFe6uyDBSEP84I19cG7YKam84sbkgPSh0AdEtVhUT8m2Z0YaD6GLGYYGA
yqJT3qOpOpZiggHB8D5KXdAydTTB802qWcNPi8itmCX04Vjm4n6kEb7manaqtWQv
7RfgzrwRKjGbFSCj3NkQNOgFH2hYR+MSRrycf4SbEZNHW2w6tGGFbfWthZ5wwnFg
hQCQH8/Zs87UClK4CTr+p7lNz/OHeg8FHS4DnDsi2fIjZmGPYMkrXrmqtEFYTJeg
yl41iEIhxP1ZLVXDSduo8RebUosy6A6PRtsOpH8Wym05IyP8Y42pd6BbGIauzGQl
SRVopBwWwQQxoZxLN1goZlmrOJz7K7yvLOvhmZRGMb8QiAUns/z3YBRrl2XZATqa
Xbmu7RmK3IUrsoJy+IFHQ8yUe//HbtqsYaqQgZ3AzpP3A8lqlDFsmbhyDTDfm/r+
/tIXTlxLKUxHq4Abobq0ZEq3PRaJW15G9FJeImkJGp8peWTp1IUoI+1GfajRaWif
V2iAKHZHxrz/DFMzg8PAP+5VvJcrTJ8UvSIxIL+Lf7iw9m56Xc3IRB61uFIRuppR
4/Nlm2COGwYmr8EoM6u6o9UwM+d6UtN8FTKCs/SMy5Dbb2D4cMKuSz4tj3BJBu/k
UzzrRQCuZZdE0XKQcNDolwNowa64/zQAjnp8ra82veTxm3Mb/CGc8rxbrxuQStxF
a2+Cx2/7gTNYkRMLeyKJ8BoZxksPBWHXdOOxrtgQbTRh6u6aespE8IODNTlsV0qt
ZLsfgdCnUF/blxcr9xTdLz+xydxTBcfaPlBOKnzPj5fX0ZOlDUQtM0+v70TEe8WP
7jOR1UWS3pUXVBFlsvk5dWuAua3GiVDF7SJfX6j1i852AwKBzfC5beievmeq2tc4
i+LUuhxyEeqna8nxRHn1UpGuZokiQZrW12cOmJuBQSkyvyMmxh4JMgcd5jyn7fub
CRHYN1xDBNExSR8yhatZvfjL1mrZBhvNGrT2WPEwStH7X2xzcuR3RGhybPMZO5RX
NyKKI6OLir5Gfsj9m89U5YpLUYro5hbYdntcX99qVjmclPotChr0aJGruht8lACR
Ex4KyLwFltanzhiGpRoP3BjI76yV3d8De8dGeHgYK7uhYJXyVA2437nqRRXt0wP/
/rJtt6puY4SiI36Hej/Nzv/+ETn9O2brzRXPGiHAfgTOdv6lxTsCmFpSe9aM2OWX
ZmrScsQkIVm9v6GMlgs1LNDsVl/H7FPHS7oqECJal+C9hCttdJn1qf8QjjZPE8Mp
+C49E2O5PYkPjI5CiGgWZ94n3ew6aeF2SWdijMyu8I/U+VbaZLq4JbsdM053UFQM
V+J7ekG5hCUZjX4EI2oKwvk2h8SprFGrGxZkZkQ0NqNw4gW/wAf0Jo95caW5nHDw
0KkHVEfrE7G1lefyhqckQyHvGs9YxcDZ5mizkbyV090SByDN0NWjPSy5iI/5hMfj
w4cQASYj5TIH/lGXLgRrUwau7okswbPm8F1g85NvXw1Mip7yJa3CsOZIjWtOJoNj
G1+fKflXl9wNbWYIAzjDOy+km10CDxqRl1o03IcY7ZTA6R+wY5/fe+HAg8iAUMVV
XC40WIFQrQwPmPBLSsK9ao9OLNXGIiVfrqmEMSnuDmYz1H+MLuvSy9RqyRz/fM4h
QCD+hYb6VYENc1JkJlLkS2mi9S5Fl3R1xDdqgdPcCjqUaIYiO8qeC1keQOeM6+Fk
ygBmgThd/tb6v9+dAKNZED+qDrgrN4sXKXq3wH2GlTcxJqkPTMCumrp0FyTa/tCF
+WHgeIoUFUS2VVNahqWji6bRLF6yjx+/nOsRUtgTYVvI3iSZ//uyFWPSFijIjnbn
dtUSUyTN10pO+1a7TOtlYjFN6dl0KkMWfbk/QfrNC0nJILHVFpWBO7PY8+obDYUW
JTLtj7pTBq8QTnDwhMueeoFQcEYtid3KgmTILA3gEN+Fa9rG+ELHa8UjV7hraBQt
GXbCUVdmApOoIG97AKF9mUuJpcK7hDFOMd3GqO2BWjbVbHP4HGU8DYLVs9JlFoJU
OKlWRnE2TmrfDG2thuRmDDIqb+LT9xBknpiWQ7HihFWEL7XuBy7AwN6MfBTNlrDQ
BBOsIP9P35HQclL+M1dQEy4ZLJ8nR6EHkLI0dCbXCO9X/CI4bMiZdFEwEZ1EXhPC
27rEEt4WM1v64PJujy4xznZN0pVX+A/IYLpdh1pZo2DSTkhsQDdFCwZXfeOuTZUs
fintykewlUOwNFVqY4kWG4pQwplYIbsyjx4PZyussrh9UQhayupYci+2OMRCBQFT
f4LVl17uVcukQ3iqf8NguWItbZTqJM6jcpXIiEfu7OngUrPtHLPVxeyaMCglHDh5
THzty7Ee9mOPzRJdydwaNvvxz/9fQrB7GXJgexH40m4WQS1dXxogCeu1JsXC2FJF
jLnQsX4u54lHKdNE3UBXdlCYJV56GOiU1gHUsUjlvY2MSx1kB/kCwGVeN3zyc05s
xJnMbFIrET/BcgQlIA4Rd1cbFggt3QhY/dKSJ3CjjVoRz74DCXT7jF4IUZj42/eU
pcNKpagqZ4cICIp1XPXxYGQIj7fPFCJFd1OigKFiAewNbcErXC7zOL+BQ6sE2TNe
bYTjr+9S8OPqsORG6dAg7jdRGD9Rb28tnsP5TimAQ17SvGoBDVID0q9pMD/FM9cS
A9VDembuYX16m9EaetUbVm3Am++WF+70KNQka/ks5gUZ50ZTLdtZezYmQHiyOK7J
YLgeaAU20DAZzokpLMk7++dByfkbrJV+5+8SHCb4c+FJ82HpH6CMjothuM2i464r
4v1KGzcBZmC+TDD1HjbFVPYcbXb7YS1ibMDeC3Ac1mTjUamlFK3YR83d3ZxI0qAG
9PfGKC7PibVh8W2pgZLJNmASNgfIe+B8rI8E6svja2pYj5fsIJf/ICUZgHPPbFDv
3cjI0E84zE0UFEf70xFPp9sXav9U1mNbIuz5MnKQ3a40j6QMRAkDZP+j2QJVIXIU
qSH+lmtlzFBEQEFYPcwayDjtGg1lDShFhFRAA1ThegyeumCbe1ffZaX2YvW7+SxQ
I2NT837nxayWM/n9KmgaUcD8LkBoqxUoOScpjVOvl3IjcM5EDKlPUkWiFiF9K69L
q2geoHEtvdqvgP5UT018yZvuADmevt0B9bWWGaSdjZ83QCF7QcGva7fMX/QK3vT0
1k6HvHHl+ITSQzBZSaRlB5fkEjcRGJRkEpHYRqJsmCw2K9YOehHzxMOC+glco7jN
Iaos9KXAhWA6Dc20rB+M/RvlqDUD5tXj4UOquTISWXyPTuu0Z4yYIk2eLLWXuGjb
sPc1opRHxeMcLuIWtsn8m5DIebbX5Fe91kzgZjGVhDx+r4FdVITc1oo3muBFOGPV
emxvGONKpEqPZl0xIA1WJf+wQa4JXvDzjq7vicJ15y/uSPqUHSWkZjUTHjHanxq8
eh+RDrIKj0grFID5+BzeN2V/XayjyAunBnCdt47iRJEPnsBqTtcXcDOIPq/kvX91
o5R5oSU+IiTsDIei43mbAtFfktbEaeunPVW4+pBeAlri+1ud2TMfN6o1Z9gzeH4d
rQncEf7Sxg/SlkERuHBpPGd/0cQVT3oUyifDGcTt+sAhfn6svr26AAWMOsvmKToo
jDB7rlqx5Wg8m6oKdz//UUQ084WvO5PwK+bJEH5+09V+I9Jt2iaGt9PSLZb+FOSJ
OUwoM5J0NiZnGL1HkRX9GfffOoKNwA8+VGBcI1aRNbfT0lkDuIfDQe3C387AiR5z
D9eGVtA72/j7TBdMhHCDzzBRC/FnY/3v5yzx4Cw1Nh66gAmradJvUdkIuWiHxfmK
D8ZM/r/xvu/6JtTbLv320D8ED46Tywr+snjY+vZxQHOtha/t+T3J44VIzpwNhQHo
onaRz/6bGo0uzTy7Ww7zea8Nhu39ljGrt2FqWpNHEbJVJ4k2NX/qyYwHn0Fv4SJk
33KtOHM2ipJd7cNE6Lg33WThZjZpIlNn3+rH2lzz9JCBrVauS+j0Uze7w/8deJNn
fWzU+0TzJtHfbNxsKYb0NxOWgciWMhnEzIRuGfqfgq5xGNVOlvmrQdivTckVtnb2
JjZEr4FXoUpHvcRWCpJLDdIr7UJLlWcArBotXXhgOVx179KM+3eB8KZiRFA0iROk
R7Hy0PF9vL9V19+jYQU3RmSB3z2QeU24mZ/znHCHLncfFln0hFJKLu7HD0KO/Jga
IRBYPzEu1Y00t1Ru002+aDyBxgTQsq7RHqlyEBP52N07ZZqOTp4j6eoGkdXZJuJe
VvHym1jGAr05sqtO2uEq1UTgROXYfwfziqZtkyHB+1JftxiaRJzA278GSFwKDIxo
Pod0b+VKsFavz3a5M2K+TSqAm2+B8K7gT4oUfDJRV7qLG8K70OjK6grAPc5Oj7gQ
BmdH8QOz54SX+taC/ttCFZFi5eRxObPY44vtdt/OKbssdaOjp3XhyhdrL5nFJJuG
VS7PQVUCt/6slQuUvko2cuKS3sV4N2HBIn9261mFYO/YXFbXcp6AzNGhORwyCYET
rqYq2rgbSRBJhId75xEK+NyqIGNbIdn0Y+FqIQD4qCM9O6FMS8/E1yArLTFmOM/r
8iX1B2C7o5zqxmzbawRkxbsELcCNf+9q/WkIEC9IO2xpZSqkc7MT2qXK7YDDoWut
e+jE/hy+hG6GqHBOYktdqczTRngi0gAAKd0IwsHzS7LIPyMcdApGTcq9dBsKWOiu
d8nGBa4HWwBsbET0O9F9XdolgWt7rN2gJoytj3wpE+udfD6s5iP5xlF3O9AH/IJs
LOC3/VqB6q4jOp/dm+gG7Jdpk3qyTG8oWtILzYTkV+mA5ehikV2fuc/AhgjNAxnq
b8E0KSoKILH0By/fWHdGqGOxbKuZxq4NZQDL5PllzLL949+fYTwFTxjhKlqruTW3
T+wI/TNlCgxQAzjYRt/2ewv00ykM5U35zwS3E16rJ41pCOOFIDJ02E6kFfKgPvdq
Mcl5uqnT6mWZMiY5lCPZl9RaGh2mxqdP3fTaia06ncsLcotK+MUg8a3NAfdTSRNJ
2LZmgM6fVO44OuHr7Ua8vzcELbZdZDAZJut7QKNi73avipTZzSXuk6OBPhxMt2+P
JA35yRUv4nvwRr1HMTlM6RufhDoH3dWeWUQNID3LFyZOs5E3gh7pD0MehgbmJkdl
/zaSo7ONvpi3PfIfj1kZzZdpdS7XrtGcJK1yhKprdeUv1aPTOJU64IPHs20TDNVl
kqfHF8+KEwlr8kjzOyLBgFfyVrhmsBTQquygGgHby0DcCKjUlGlKMdAPqlIO7Dju
d4zr57QUR7cWYu58xWBl5AlYChV298hxKoqnLqRvs5HCpyhBfc0HHrEzc8rIFW48
PbdePQ9P75vsulfF9BkRQuxBoOQx2aeehbqwuj0fGhdxgQFSbKb0qckvfnQhDEKo
rWfvKkJuaO5ViNWaM9P+UzxuCw5OC2QoJ7PxuirIWnIJp9ERmSn37vO2OsHoY0Cd
2vbMxJH2MHu8ABEe0pMv8ibutf2QVo4miiUr6NiloJugqjg+Fdak+Lfp8FKIs3/D
yV/8kQ4sih69GqXqnSP40U8ZoczZbX0ibvpJ87iq6OYYrce8vVDS93NvH4Nvp46z
3npqF0KCsFIpfFiKOs0EW6e+0+JisWZb+r4LNXyOEafkWhd2IzUdRlCmF+vpaD4q
3w258b7HXkP//Ldhx5CH2UcGrOB1Cfwu2owoxA2ksEFPPuZDFh/4ec5+WAcz0/P8
EN96MX/6mxRaXbNZTiwkrfGICxBNveVlUAh2rDzkFN2dUe9e2hm2v/wEowHyKIrG
8/Bur/zF0K4r9en4plDzgFjq4gD6kl+ghP09JLY0X3Dg1Az4drMHU8+99Eipg/m1
UBFh+BmT/47D0AbLUxoVg24QdAprhVjIl+O5vyYmC1zT6mXFmGhulFHFNZy7ZYi9
xZYZIGnU+IYOFVqyXd0cjLc//dYZT+YGK5LUbrJnRmpgmvvNEhBsugAQ56RsAnE5
CKxGkAyCcvMW61Yqhe0/l77ZKDO6wmHRAqdah7LBuJH0pXXWEZ3RdAIQxcqfv+yo
NYJ/dnqHVFiXHCOjTbG0KnxZnEXrdT0vdq8wV9QiUquTU6X+i/pZ3r+GGWWHyEXt
mfG4VTzDXBfPOA3EvfIi+/qLBME3uYyPOGNgkisg6UjsuewiOrkmdJVyOvYm0VVf
StM6aP72WSvpVt0BstH+692ilgsED2NBqQu+hRvRDvCLqjMVT+ZvdZp6VMTqlTov
kde456hD9UMWjP1rlhpkMBqMpwAbEyzND/CCkfXsvaOkHC5chtNBLmxW6fLm3djq
0MGnCcbT2zw7bknDA7ODK9k3388dK4aLzO39+SE2ylBP5c1q81Qnc3tTGLSznGk/
j6oKQNVCSZ8z8sYzoU3fIazMEHe+DGnBcNJNN6PMu2j2R4GU1Liwwn4sw4t5fHo4
HOH2L7g6/7u97ncMwAOfYGq4zcGXhtypAw/kHkd8Tg4hmSEQYkLrEmLMSFyKQ+sV
o3ubM6zWB2oy16p5WRiH9FW89elAkGBG5HB0+rJq6dmGyETKH+KU9kK/pNLUQvY9
2+tvWf3BuVuxRIaONyo5d5BTt5dXQwaCY1rQmHAVJEf32xaG0SugLbNzIVstNkDd
i7EjjRepLk0SsDfDPnfbg92+2k2nefu7TpGUtzVF+iPJNvjZm3ySwChEz2oO4srD
m2YWjgAGOQzRWAWST0D1OYO+PVfIWrWmC2Dn95eKbuOT82WScrom+q8HRBXFgWL2
z+UlZu0nKdwVHOm9bQaOjOVvz7lFibNEGxn7GSU7S5/5VlJtKPPCmL8h9RGe8Q3O
V0M5qCddt4A1+4QNcyaEPZya3GMO5mRrQIUHLz8KJ976O6nemsWPwpzMYSvzdr6A
9IS1yMnLPZylSyV5ro1KpeWvAzOuYgqL5qJ4SYIfwK0I5qZmTnF5d81hkrBDAGMm
5mfaa0tGDoP9F9haPWSaiLt6MczyhZfBs26kKLti7i+TF+5b/XDPTeXG3EEza0HE
6cfxVoCeGmm/zaRMojGRJz4tKK7gS1gkkbvYHLraii1nHu6RdXwaxqJUq81Xbva4
31JKJ9zuzxFODd6T0+fnZ6O30SLnkUDTAhLb9wZwp/7RFJy7alG9MmApMY2gNMbp
5lxYhdO8Icw651Nit504m/hpsMvsSb1RgyCtUVB1S4nOLWzATHLKYr8ZdDKlJ8Y+
sr/4F/VMIcPIWKq7QqqKctB/DEtVqFgNtuKGmCmG3WF5L0RKWJm14zTiLlUBTkZ6
VgDpywZFqjrByXRl41ffR8PncXn09hARANJacAruGNmQos42KTKWoQWj0D3Gonhv
5YXer0CxHKOOTuTZSPoFAH79AWrnbhMHZ2tMeM2uBflqaKhz8s+7jqdCf+A/EmyP
4mIMEf9Xv4GASv4KJpnNjqDstff7e3sAmv2cW4D9Jt98USXrBv3njs57uxx+nLjr
SsgEHyauBTjbBmQib8JNKMIepDQ/NEFIO8PxEXFLZBxgbiM15r/oqJIkxjs0yT2+
G8m1dhAWuE2o5+lyQmOykMIq+CUEKjXV4SmGrCpPugt7B7WwcwCTqvK5quItU9Yo
4mkUUN8mMi0MGwUX9VYschdet0QkHH3DsHOxfysTPlRxtOV06n0NRpYOdghCBTfz
J5dMwIpi5y3GaIpv0/haHyGrt84XV0JNjNhosu/K1PoL+Z9tuA41nOuMd4m2cB1c
L4C/L7C2hJyFAC+1hM7b2NEQ67GgY8LaRS1Exfxxg7PDIRKZoudWD2oqDccGn3cT
NOcK8FJBLzXA4FYYuwjr1Ht7pHm7h3XSI4kI+xlJuURiy7z9O0r5HY6BiJsKnAYN
Naqh71XdE9jf80s2udszsrf6lp/Eb8DIJEacsCXSEd+g9HVokNM0PvQEsNkIYUwn
mPdyog1lTShM1nkvhWiZh1oSCfCQHjeRgszP+hI5rlzskg9K/6Z4SdVSuqbbY77o
aG17FQ28VmPVyGAKBBwXaA4nEnqislHbuzSLpQyPVkQdIMeimBwCymxWE43zN6zT
W3BN8Fc+FuvCeq0wMWc9dtjjzde0H0BPJOU/tRxJnGG2Pu9i0jYIWYDGj1J0Xhwd
IZbFcx7fAUhRQwrAny+xS2zhElkLKEH/Yl5QQZjbl7v7jDFlbTD4gyRq03BN8Avz
C/hIdmOAS+DJ963wDJFpitg+IOpdnm1jWvM0FgtX489Mt9A4RfdIcise9XbBvZbB
Me+oEJLiCWn6wTLeX68ClMZEC3gXvOfJXwJAbU4S6HJaQmoli90zNZimIGwTta3R
biuHohz8PZJUATdk3NrcUdLNSEWM6+L/3lwIsLGabj9ZR0ynjW3euyW02sQRjE71
9OM3TtE4MOGqw7aq+vs6Dol5u0ZxD3qiQyitCSFUzj8Csi6gFRADj8aaItZpTUDB
TAtYXimTCszP+Yw56VgSsDgNOH0JbdlsbrR+v3Tk1iMasDUdW9K1dZkdKMpxbW9J
oXlvYhaNsPCUXniD9gnNwj1141vsfzGWQj3qn4ufLFF38iHXl/y2xAzK6wiY+pIN
tvGJEeuOtL7QFIzd821tna7S2xIW+skw2zT+OdoRtGSusrMptSjUStxPPxsi1/3q
9luDTkH2E69WjC5PgtvWesyxnHAkmjqLrWvruen8OVPeHDdE57S+E2eHyayd6kAW
6jnzijdvXVRjI7yVT7noJVavdH2jemZefR/e7CRFqn+FM855n9hycjoxbE+Q8LoB
AEQIH5kyiSS/DvrOkFIfauluB9rxxJRH5kKmKfR2/ktDRe0FbDigU9DJaZF7rqoq
ChKMCBiisgAAesso2ROs6QoxPI4VcQrhYmGrnqVHB6FMdOWO0rwddGMK9x0TeYVT
8+TlHJRhNl2DvUqmWA7f/GNo5nd/Ivh+QFgYbQhDiVR4zbT44kgiH/x8mFpyEIYu
8ooiMCs15j1GqL7WDBgXHpFB0gJvkYLsokERC510ad/PPgNb4DaJzs4ZO+66UuJD
y0GGSkndD8lHVAZF0DEoX9IUbpXLPoCXhWfE/R8fJADhyCdvA+WfgC1TvMyFQOrD
mDIaL+4F15ZvmwWBfoq8tJunJv3QcnSa9lwJXXZT7jiYVjqZVKQ5nARYnhBsvgAS
OJhpPVv+sPsXmNtglC4vFQa9m8aCiOlwZgKmv80VeD+1TnPPqh7vuRaWg3RnLbOU
qNyIOAE832yeje9HLqvnqo6RMlAIlYh/StkX93lu824wB7W9q+lYcROMY2xZkuVs
I1DuvCONOhZVAfSOxleWgWgIVoQbKPgSd5bcbUrf39hF91b11oC2Z5h9GBbVBsye
auoEX0IrK4vtv2IWOht67KWjJGyEqetJDp8p7dD3QkR/X4kvIYUZ2ptHfjrubrwt
grmErguR8OdxAEfiWkGwA2TsT5RKrSazOgbNfTszjv83uN/xuxLAGMAImiOPOFt7
/uVzHuoFigkIp/WoOKWFkh24kjQ75eS/6pXSCJouKjZbZgu6t2X2dXys0OuDxTE0
F2JsqhT1OqgwN/Q4UBLsbBFMmeoHcr8m5nrog0E6nb+oUmYGVOamrBI2Hhxy7Il/
NFJFajLqE3BluW528FFHwHIGLqwVAuGq1RMP0ubxBgowrE/Obo2OEKvJlFsuZJHq
pupfuAxx1Cw+nGl2sNRMzS/TvPyjZ4CT8/AaPEgY0gY=
`protect END_PROTECTED

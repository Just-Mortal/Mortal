`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6oE7Vlp/c6z/CZZ1oSOjW5D1uvfy1a5hbJ+tnycjrtLCPZZeIMY66utJLhvboG+
87F9ryDD2gfHTnFnxo+oXFkzQZQvv+B8XOSDYmhRwdLaTjjjUkKQVMnpXTfEskDd
Uxzs6pOLBMonjbXW/bP6nDeLmekfxVfymWYesbfee1FxJxFO1mFOqFMTz7mqJsG1
LaKX0dYZPWeQfZ7cmcqBRaEUjhDrA+9GTFyF3qoKX6VNTXxUTpZZrwNWHsQq2grM
u8slA63yP8q10YNUci/ufQ8ium7iX4vJcZOIieXjbjuI7IQFgGk8IDIchN+o0A4f
wZsZhc0bW0IzF9hFjeciM/i8aJDbVMBnm+k65j2Rq7zXu2eNWI6O28cN79UgQp6Q
Ni/z6Vurxgs9t30lXgxxKH6zlmOvV4PqvaGIY+IPF0F2V6c9qSEgZAOArmQ6S/FK
4VJ/49SPO2hp/JTO6OVBZuiQxOkKLFQaz2Cc/8VcTP5U8RyKViMlgUeiNEvPGeRD
HDW7rTAOZsoLXz9b+GPy2wChWnDwXrsx0fV6dLOjGgF9qKR4n7LuhKuPk6MyLDNx
l6RqsCnNeoQzYI9zqzdpR1LOCFVWZ6m+Pw52CA6XtJerR0yz77vNf4sYtsL8DoS3
w6lEvaD/M5UB0/TdMypxiDp3wN2fcVkWr7Tq1HiM+wKWTfrs7j1nF7QeKo5VPK8Z
2Rk1L+re+aHfsWPLNir9BZZsXDbmmZ4voRR3fXiCEoWN+YEUf6MM8Q3MpK37zD+8
nZlJd8h8QR5/UhYrYZOLO9+HdsACt6pBcHiGUA0qA4Zgpr+mEjRv4nmy+et/cj0P
YlWzr/msxWhjOhlPoUb0VyolewiBlC6GQHEICpP/k1DbuIDbP4JejC9zeMvwFTb0
cWZqOuS+5NiOdz5rvyOqDALpuOL0jRh3Uir0uZAc23PmNcrW5E+WJmIEcl5NZJ60
JMjK3nABO3lsziyoKqDSjI0m4L8mR6HGNIGivT89HCfhW2N/oD+8Of7HG5WIR8AK
VR3Xe71aS9OYG/ImMKtDLb2SAHCve6x+lHhKjOhy6S/P5tyvJiOsoB0gBGrtj5ri
iiFroADsmbsHxpth4wf28kLe8j4z0cofVpKRIXH28iW1dfzQdS10XSWkHxFixF6k
+oeOONjUMyhuMbfJDax5IsbJf9uCvrNavJaCD6+pehqBO6IOLgT6SitAorrHmUJ6
fo7yJMjsDRUwmJ3m1wfpznnh96k2W+sxUt/T7PhAH6tK//fmwpxNVhmW2tA3Dk8E
HmPpeHQbkpGElKZYRihhNgJE8RY6D6RmrdTEDNQhBI/uCNI0pbB/nYEYSYDolPC9
YPN/tmK8ohPVc8nr0BsrV2b8DkFQ2gIKqywKIYEJyc+0M+Ih3UH4kv46GRxqDn63
D/+TWPzV+d5rIVf3PBVCqkiQr1240Zo9tJKgMdjIR4V1iekFNKtHnbFZbGpVi3TU
`protect END_PROTECTED

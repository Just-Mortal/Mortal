`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rjMj5Ob+Ob8oBdVu/bwTUaVlLD3X4CK1SjKBdF9JDL1T+3B1YtzQy7tcrz361IXs
f0btx4alqrlwjOfsmB862KrqKDIM134WWe28sKX2z2hFGI5aofjWqVt832GYOzig
ZLampAWfHCqAaxYaeQhmhjDQD9zA6pBvQdy6s8t9OVOndLOIXFF5ysk+5Q5Jx9GG
Kv8rGRns5gT5yLgBTGYEVKXG5BCEhdHFBT67CmC+y9EsDaoFZt3bWWR0cfCfMPiL
U6Cb2P4GKAMQr2IBWdMYC6WjwolnJxybzaRN5LlpBXULsS8HX2Pnxk29wJAQtfP3
AkQDEFrRHKaxl0RBdW+cErf603z4+Z1AWcXvYG1uwr3dnG4AoLfJS2qDApiVbSC0
GgVBr6EdNmwUhOxI6i4yQefk3YqEY2PsbI81AAQXkDkyT2T1VHo3R+zoPuMcPryI
bPfCTK9izcEcKfn3FeHwUXIHb1s/fpi2m1Kk3BjC8z4n5uqn7UTixz5jtoaTlDRl
5Ruyp3wFZcofpthi6IjkRnS9EecV6ZFlare2g+ae3Xtzx883tD7qq44ZntZPpvXt
DxhZr2L9KoMnBcAHLuzMBZu8IeRESoUD1jN8oDEkx19qhCKld0s/DcMlm6BM+C4b
Sk/d9MajY2KA0D1KJDaS0tArBwyONwoQ8xGApGVraPN6O2t6j0KdkEGeebaRvkyU
x1hF3UIBJCLpYll6rY5O8EaJnqw0ZBD6VMrYC4X1utI=
`protect END_PROTECTED

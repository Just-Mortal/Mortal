`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1NyZQslcKzisi1O2EsycBSDgQLD9VQBIP87PNx43fMqjhKNq+RGAk/wSwTxTC2vX
QDZeiZ2HjaI+6gRSQZq/AbnjcXUlm5Uq2BgpPYyONBL+Bw1CBR+FMVud7CRRWfeN
G+ZG0RWob/BLg3z5La6lc/0nGLKjZDbNPAHXmlCjo/jOk0lbUD+w/lh3eVfBBhKf
UneGgEHwAeqG8D9YqlOOX7YOSaps9PnOZsDkyodTHu/c2GR0uBcyIQfhmrCHe/Ba
/4UCEzBe2B0ntu9IjdgFpBfY/59cgid7ESjYYNMQ6h3jRlPIye72XXyStLsx6C2o
zsHgWOCQH+RkVgkClfztrD3yJXBtcBkHYnSfZgqZHT3nfFuVOclkOxEZM5zdQXlU
IwfChDBoJVjv5g+IXllyAnvgSDnn2ohbdtJ4AwlAW/D74BRT+zUNrvp3t1Ci+PZS
R5hWuLW1haxSBWScWyi/TA8KLJ6JFvvQed2dCC6LnKgycAo3ILG9IWMNDuAsCi4z
0YfMvaPWj3kkzk9/kEYWpRmrqdf8N43M7JfnGKUV0Kgr++hB68////1q1DTu+lyF
VDQwaU0dHL1k0WOPhKIDF1W0i2tOrJeQTTrqY5yjZmNSRm4fPtm5LwhXqdoO7JVj
dMjg47hhXiU4DTqxYveIeLFuJ9hU6oWlpktw+LYdJKJ7E4n/nM/E/+RqpxpzCYvN
ZN5ppNXRVY1rX/vDKVISzQDBRgNANkrkFNq1kR4cSsONhPJeg8p+vzhfNcBQOW0L
W6+HfpjQs8GUBRSINttNFH6T6muSGAWnlJGbnM4m9aB5cZTF6furEIqCIT8fiSWB
WkdYjWdok9O57M91R533S8d+uPjDr2AG0mO2i+tufNpNWy/r7L9Hf0uVHexRqLTg
6Zw7QPLW6JVzTnm94XvlZJFf/AkulDaxxmICH4g9Buyg9lEbFpo1nUQTnVqU4BUb
u6klfMKqLtBoMUIV7iO726hTNUTqdB/7/uz94S0Jq7GfmTc/wIvHTRAffIpHBobQ
VB507Vu07kOdP0D4Kez6Y9o3AdiNj8fjULmdwstmsFAoyESsPsrBrzohoI99pfH0
2mLLCImk7NojFlUN3zdUWEw0nfQxgx3pY5tLlq9/VMcodrymqqUpb8kgkEOApM5K
NoFtME+DI6hDWZsdTDxIuCQJK8Wyu7lWG5Z7zAU3BbMEoCO/bxrttTf37wJff3it
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJVwxXCpoJmJtWqepf7GQuZADf1hIfhPZsuRBpWzmbNRl9Ywd+UC5IiXT8qhcdAy
xAG81VqEuoW7LoLPITaaVbdmJHRV9MGlYk7d9Ss5KwM0jykR7j6cQkDdMjxjUeqD
SjuDOn8aAu8DNX6tbPkA9Xjs7nlintx2X6BNLqBe1JSPBsjMzJroc+hxl8jtM6Ub
MclIqo62T7bb8FZ9dS0LlyMkSXBsKCFtrR1DIIFeg2QBdRuXRUBhuWC+/HprUL0L
Adu4WxyPJgw99D5iywYVqw==
`protect END_PROTECTED

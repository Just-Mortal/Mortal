`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/UlfhLfAXvuXT6xlSHBXgqirdjKSWKyBfXB3QqIazs2OU8N3Y5z95fRNfyS86qG
HUluLGvOoWK1kQ6PtElOALGmDNBHRNSeqoMAiYW225k1TcBJOgTldr4HKxSBBKgl
PASQfGL6XiYr3uyic+nCmkVCd/VTcCsVt5M4odYaEPjIp4jnUzb/lVgElQq9jbn3
x/1/h/Tbp5BjnrdSVuQso/e48cju561J1HQCrc32A4cHrAXqexMl5CGi8hr4WbHt
RhEvHSv2itRuTZtOK143Lle9GBSedqTquwzGs1ct6PAV8g4dSeRxejod13WXND4t
AKTHAOa9tjKuJ0CLERxy6gVt47W+tOWy0tqoHfxt5pk7KDZx3jl85Bbg0lREnBXS
i6QuWXI3nf+eaD+pGQKlljujxa+isomOz/MQ5vnIKRhLNij29RrPudxYk3j1bZrF
QpF9L0PW0Z8tM/MbbitvJLsgIX2IJxIYowz05yBKYgCPBSQrtLEX3kgmAcUDEipA
OroShyNC9hXRMJXs407+PncgK8/Nwl2Mf/ikieEX0vKSVLqBB3yyFMHgFu/p5sUQ
lBWQHL9U+nwidbogUm3EZ3KjrSzoy0JO+PzN7cbBhNjaNR+n11Lz1zX7C4qP3dMh
/c1Wqxwnj0578rzpz5MMJ/AmqozxVbr7uexAmFFEa1pB43LU2VEIEFjXWPNFa5Lb
wM8YLilABr7mYHNinR+hGNpCw5IEDcuoxmUSdkpeiPt8LG1QnwXW0m8SPy+giacl
3GOkDTiIcq5rAMqUjJDgdScMxDIovzvJIm5d6QzRt/UCoXyIKCD3s/htVePQeMui
ibOgS3lrAHL4k7vD2q9GXNMn1iiEGozdelhimATeivoQSOA/iIp5pnze7dHOwtV7
2TgHMs/CDZ+CqpA4sfseIxUXCs9k3ZY8sk0TYGNuNbAucleV//Bs5gZQ2j3sTjlZ
OKujFqqK6kY5gNU5a1QojBDnJrHYmz8o79wbrG9vtb3EHUysggip3KN7G1rzpGXW
+86QA27cOIurvx5ZQkAA+ZN78tH3z7JhQlNwCLjNB6bqOs+7OKwoW1of4xksVCrW
sgEOZSjhxvuIkoqZO72/2lypjOUaUOEenbc21YC0oOcSJ68ih4/ySihRX1EKaj/g
bEKdYEucc3nlz7pJD5M3LsJrv3BTKax1cGdV9B/hHGZUTx5Gtuv/IizBSqsVswTz
5tHwNK0EraHzSCpFU9/mI9+IrwzHZMuEua0t7It8hYVG+mwdgsxzavwDf2bb0UBv
wHHlYl10BUaqoAumOq/uY6wqsqKmRgIEq+pY5w6FU8rYj7+jzSSngNK1dHDtWKDC
xcfYJtsaYORxZ8y/yl8hOrs1Z6JNxew2MCkKeZFBloYpgksmJnQcW6DYAnoB2N1T
5jJ/Xs8A3sCjeOq1rvS3WWBzR6R/MG2WXWa0ZkQxHIVj/r4Yot4jh2D+zbjzLqyS
5TJjJNlnwKgsRrAmVtLTbeq5SIGGf+r15NS1YoNUb9LpDJLCohpptPLte3FtGBO2
Xk2GogGoc8voZCc9wPf+1HRqCGqNWh9+1E8eez67C1kY2CDVDgsDSbQuGGgkGtJ/
NtsD8UbsdjHlUYjCwEnFXakjxf9t5n0N1Vihhbso6Ot2qVKMF9PEpfXHaJUOvIvy
ri+ZWwJnqE5cwEeIHXqVwuioqCILjJXB85srFguzySJvqz+bXC/7P7KcNmrUAFrX
6sD96mZ0Yns5bflD6JO8/Q==
`protect END_PROTECTED

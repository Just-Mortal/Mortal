`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqZv4fEp50X7M6pJLqXzKh0ezgC2NOvp2sEfLsekgp/khJuNmCkTLpvOXXOs2hDw
xz7gOhTRuHGIjQSgnmFJIqsqoGfAYCgLif/iry25V8rczanmm+ZVHDM1ZCcntT3f
T37X5i+1+TCqjNN1VfUjqyJpsnzcwoi57/7OV58iSQB6AaeugwYqm8/Qcz69AF6z
v3oujCsImXofn/lG5V6ObIRQOB2N8AEFsFjmSzm8fV4fH+bjtizLxPW7QcxqEmn9
TrNBdmOejXEPn5pJZGgSH03buRndbSisnv8imxfdwMGCIsQ1fVc1l5NEZ8PGDs7k
UEV6QE1dozTBYTO8XRHt5Tw+NpjS0qfmo4OpLYXIzoE/yE5NaFTRzCsJvaABTEpK
oOARejsSa8QKXyPkn3+c+BQefGpO9N8lD4Lp+6VkKn6Fl6ilPgZoReZyHeruSAaq
V/KNqLvO4RjwfDI4jc1Yty92rtbow9Dz1g/sSq+aB1WPfoBXuSxpSXaQvMPAW4tH
Fl+y4rfMTVo5roYKUeFeocZpvCpY/KWHac7HHqx3s2CMXttkE9LuXnubyaLaRdtq
Evwso4XAYZKqu5CqhDj/9TVMV52RK2xNo905dtRoydIrSjVpAkeNJDiSC6KjLCBF
GKuCBVWxcMQkjH1OZAe57j2mvVqNK+3sCaEvGkmHaBFgQcaq9zQJgptQxi7gmE8U
vB7QaQ5sqrJRaimQhF6JrZeuZRmaQe8ZTlOW9B472PjsdF0u75YOvrwD+i2hfQ8H
IeMhE9IFsoSAie1bxtE93g==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RsiCo50Y5D2SyFrkRvOc5RbqjBITuPzcp9tT6ixeMFeUbgCsp/3tJK3zSnXzW1ws
nkywDDv81oR9jgl03EIO/zHFVc7/JobK7sDcbG1LNRqDASbmTa0LgoU08y4tnl7+
fFf/FjXFoEIHMyg3kF5sg9o4zbsAhTnb8iEwyY/XGq/TvIJW1cCDukCzaFxSSUer
ZjNrkQVbHRofEfMlGDlQ9+7MlKbJQNMqN/y5AADatqIQgJ30Ejb9zNv7c4R15Ahn
gXFRX95gFyrunKGSAQNXuK07JzJoc9Os3G5xiTCk/G8w4WReeURKbrezy5Af3q+o
JOaFDY0KVD6UsuQlhr+iVRc4CoNNxMB/r/iaqiCgwgy8JY6eddTNjHgwJ1+V7ZOV
oSTn7V0zilDxttpDTeLMgEbkxjZS98RgMl/cWzAlI2LduP+P4jeJOQYZ9xwxY6pX
28yNcyxyvHIKz16hykakJ0flZtpinn7hQKkabggo40VC2vH/bEVQnWf6+63AzvxM
ZkwATYu0Ds5NHZ4o9sonnCYAaymT5lMJb58lNAPD5i0vKpwuVI136I0LavTblNI5
UXWHeZVhyDL2RWeP23HE0tLtQ9/FsUu3ox7p143rARlUVaH16zF/sqsbx9Jk88tR
qTAi1gGDrlLpbStnG18vW7uQ34ZjCezMEAAoTJQxwszm8K5Yzd+/5xCSXVej82vg
n5wCLSGMXdfMYqxMz6tAAuCgh5QSbB6vT33XVixpI7E5HGdWNH1w80k25wmFiB5l
STyUUH0VFVFv6XgS6rFJnTacqIYMs5B802/lOU1voYqT7lYL0Y8lhjbWq7MQUMp1
mjt6odjwOTuGiN96fARmVtzM26ZlqLFejyc+c/7xesF2qUoa9xnMCMEg3/XKiJTH
RXuXKKINz1jLzaikAh8s76YN+bnSOXmq5JpjLt4gb24oUhcX/dEd8H5CV2r6pcSd
TTkfLR7vokwuw7DJShWJi/F8VlUZBzbTkj+Mwx/231I5UgcMalkoye5GiTMoYalF
7IhgZ0nJ4QNfEIoHLhC1s+umjTepaUuttQ7uvgKdf7BN/lFWviTye0FWcQ+CJaL6
GhFHULM/JcMeoEjPskIF9G7RU0smGtZCT6hBG/8rxlvCpnJckDdeSrw7kCkfG7Eu
XRhWSNhhh0Bk2BucQku7CX5ECjvNB+wK+X0XlcBA0NIGcOkUzD7neB1GlJgKbUrD
95D1qQgpmMW4quhVsLvA11N/pSBm0x7PRpp2E1KSrjXcixcgdfxx/5T6To7A+NSr
tgIXp5orpta3vn+ezId/zAxm3j+kx7KoUx9LNTXUOesGL5bJD0qYygJrOlitgS+N
2RX8EN92dwIEPO82MvPwWrkh2aSwbPALQtJznCR4yiaG4ApYlJ2ens/+6PD1exgi
YPH3wHWf/F4pB8rtsF0faqqi0VgPLhyaZcUFAgOjjiQVfhgK9sx/8VrP2vQm7NfP
zjUWf1tZ4qGWgjnnQ/5G0dMVcZC6mSpIlSvCNpU+Lw7naJh0z0BWtLqZ9T4NeOjY
8YNq1w+FvUUymmiy4heC/qIiUeCovQL2qTIRntd+gn7riHgu+rWBXprwEoC7uso2
6UQED6qOqqENBuRUypmPxmorZ0DBhuKsHC3DcKQtAwVJdbVauauJNuyiBBvc4FwI
meLCkN7p0Fv/JKljRo2PojyowX3ZGpjgMKqC/hItWMwwpcId/KCNdudTWPgUbclS
fETQDtdZ8D5zHgrtNfK/t4dyMh3BmqhDE8blG8/WOF+Zb+HsE1jc72inDSy3PB5R
c1OYLIjf7DeBHmpu64A1/3eYu1AgWULJvkPwfPfd5SkeE5BQN9gZTsfm9op7gj56
LE+6H8nsXtIi2Uwpd5cOro40HRV6PQBin3zHfUke+MMRVx2PJSkv5wdPw6E+FyI1
JFJAG6gpljIhFVY8vBza9GUzoiH0+TteWnICUbN2ROhYDoZhu1brzehYrN2HM31t
5hYacrApqWL+bR52M5LK50oVAg7BmtwIBxcpM1XvXArXijJl2XCqmmv6DmfoMKcK
beHei7DDsHRCLo0ruE5ZTJZpSMHdeSIoLRxN8GyX46+z4pPYxyDmIO1xB8AGW6gD
G7r8stijrwVLS0rqiPzWxb5y+rSPm836Urw6OaVm+WBxnQ0P/9YJE0LxxhNURg2w
+XLjVUA+MHJugMMXZOy6qOHsBefTa4/hUn/s1nBnkoMrWGGzV8dSRZMxAWFmyhLN
JHbR52PEMthvXw/Re4LHlQIlG0LOdB90l/BH1xgPm6dh8+7Ij7NWUPhhsLSDixnA
R4ZLXadxDjNSO3q22VeB6vuKIypJtYrfe81wBRw7/x2TcSlYnvz5ulfvnrf91Cig
IcXHwOhRgpVqiridnO6QNpjN/0PIKpN1Qdl4aS9BXIDHOpvwZsk2CXvw2RSfMwqJ
nN5546N01dLw0gHzPg/vfwuygdcteXrDwYofrl2SU2coenRZDW6SZ2uWL2zSPfhJ
Pr4vYp1swdlwEkAj0RDhq1/G7rCmypnW/zYc4JFcFA9LQoI2ptknH8gD5jzxnMU1
3Rke1CIsbTGKraLImljqsBLQJQi0y92+nPyGdXA7juhln/6ICd7lGIWuhjbLVy3Z
Id++gZpX2kraq1sAoFJ3uXd3esfVrbwgd8GUrUMS5gXmkUtgbJwrfd7cRK7uXFz3
h6ldNUYWFr0CKdKcejKvtbFDKvJyGfFlLnmnfRlnrb4zIFRgVN59yEJ0DZhOpLsJ
FCoVPdi63TURGuLV8SIxOSvKN3cRnq82es3LLOWQDDq0s0D989H7iMz+Kr+c2Q20
KRvKzAoLRpiLBtjkoUSLBARlmU2f5jwz27rJ8wO5rgWgyt5/VSRNYPEa1ErMfBG3
7Jj50EPB8S35CE0t3/vQcxyafxTvP/skW6PPqx4t6DMyS+d9hrmt1ylQeejk5I/i
PuxGptK2vc6/u7qR83nwFRQapFbHWZtDGRgeYiTCg4sx35lmc6aLS76In9F6O3RC
Mu0DvxG93uKLIjWCIWru1qsNC4QznBaT6Vzr10kC/BjoNzpUcXKcFjEplvnXew8r
0G4i4KgBGgNyNlTAXoJSYTuBtJ0QnOIo1LRIj3aHkWY/m+usf/Oun0niw4IZurNb
7ImO9OhCbS0vM58/yHBPggGjzdchuwgzWHS1CJzOqXtOUljIp+fevQmC99UwB/Xo
v5/SUdgLXr9C+TYxlkJSMOTsN7jWF1w83ClCAZoBJMkL87JFiINYwWQWAvrM3g/r
A5U4vZ+7f6Pri63kNfIrOxQLwdCnlKlZZnBACaWB2VkQUx1YBoyB8UQDSVuwD+Nk
MHA10w87NF00ZdJqPGw4Ryg6Fislu03bEQzusgF+UF5el1W0UfjulfI06ro0ORZr
0m/Btrq9ewvwbZsXSfSIybv9sKw9TQPpflFIshPvxC/LAHQQfOtXDtA0MBucuTEd
VNl6gX5HfZGISwGHqVEOjwlSzZOdliMRMpovRfH8XFOpERKyhZHYm8lr/1OKRxRy
D04W1bhxpsK/ftZvlOSVWBM4+FSpd5jnwHwYV9qJHD3E+VQmnqw0Y53OY8s+xWPu
2nRYO69EOhxKjQzxU8Hpx9jBCWNjqE+qolVKShhevIjW4FSS8/73ow8t/oQNnhMu
Ku2DKe3waGo32czS+pJgzmBCVIqD49T+YL1/ogMjWOlzJcRzm5oEqtbqeB7dBMa/
ZWCkK5ZapbdMgcNvL6xSbEqNwQ33ZWdL6VICxEO2D73JKnQLTQbXArXLV7iqYAkp
Yeo82BQvVjgNdBofevOL812MhC4b1LEovvwGCjCE9lZTc2cfdy3P6SEPt2fvKab1
wggk2bcMNJMu+0RsRuSp/GuL/VIqzHgieJyP9u+p62bBcCzkKaQeQO9AUdRQPESK
0ULzs0on5GhuePeBBxeOQD0MV+X4SJwE33TMK5GTk+1nOIDH5rmXMsIpTLIvQ0ae
1fnJe09skWyINXhGPIe94nDa/0FIZytSyv/AS/I6noFJNgiVRi9vAtPfMjM35cWj
VAYSvlUVUmesuNLQy387C/9LcYFLCQhiHWSHagIf3eQy4xMf9U2VQGJg7lJTyH4T
GyxvkZ+HfqzfEFCRuZ2eByiZmwXxnJTfNryXCtqoROA7dSc5EtsRE/8MrKDm7qJU
iuHub00D8zZ+Tk2RpXP/4n9Bms7XVCgfWh1qz8bT1uCCX20kghXWAh4X10VrQPW9
5SK8UfyRHzftQLsjo8T8hfwwRijZPmIwCKmdiGvUmfp5zWtKKDVhCh4DMnJJnUlZ
jaPFxa9D8GujbTQg3fMJ50DPy5NSsWxBCnR/KRD+Wr/S6xvPZ/lP8XhH6hf1VO0u
UNn8SZTAWqyFbYsvLuim1FHffmFwR+kofT9XyDgzWXfG4H+Rml5HIzIqg+TuFEzF
UlxWK36NoVbYCG63TGegXge/ORSU8MQNXPvE1XCf7atsMNsTBqLBbN8Ch7KQPsrJ
m8lLrzxBPNqwirZkbyWE+UR3x/0FTmBP+ZKvhueqQVyGyj9WgNAaOx/u9Y+BoNL3
Wsk882zbkugTtN1lhn4R4+9MlFlziq+HKVzhqEA7FQBu3c69Jzguoh45kcsILpxZ
K/00OPoI70ivL5HvxjPJ66PlybFqB946mzIs1Vz/DOFytBPsbOaZISl1EGkzHIJF
WDZcudzsndtRramkTy70nqJuqjMA9GQuV3B0f8nM1XB42laijeFIZAPx9gGCfOQr
mA5GD3lSaUml/nB6Yvm358TIwdPH9ecGOTpeGmumoNDpAUQJQqcs+bAr1yN9DaAK
b1FXyNvypwJ6IuhUNvbGmSdO1d5pvwFm/XVa1FPfNx7slh294p8l4VWTsMuqk57G
qkCOSjTGCHHsoFtfTibWcA7eSCF2p9orCS0TQthMfT1YgiLOijKOTgkMkQdQbIQl
Cv5MNYofz+yucIY2BTEhu1fsIhWBaV4CmrpdOasRgzlMwxnu5OIkX/j1NaQjgPuq
bMf2/VGviVVI5iHDiUV0UvcSYKAYiNpDU71CzvhYlPMpfRF0t7Ck698XFMBoL8Qv
`protect END_PROTECTED

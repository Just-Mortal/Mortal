`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r1aK2bFfgpYl2Q7GiIEI5Vu4fRvDxOWEfkzr40sE7rcN0Tu9IcnK6qwFPuua9lp4
cxigBdCmDJQWV19AP0gYyHdh3CBKjPB+/EFqDcM+DwYDBN1tC61HqQ26+lWL63mX
XohePpwswUjWesGYMH3v1Dkvo7QPZZTV0DHDxQNljB/xJSTicF+pqitiAf/51OBy
TlAS9z6a1Gc7zPSfyd6Ji6AUCX0YyKR5W4gRKegk03w0CVXuZxFAwvOacsY1wKFZ
gDRxHBMtdRXLNNdGWVdC9w5YGkYo6w/SLEIHzs/X9t4p9zn3bVM3bU5n/i6wzydD
nJQ7n9CnJfGdN0Wwdn61Wpt+QMOTmEBYqprsEUay6SstC7Ih2Ly+58RuA+kFpIsO
aIlJ2wjOAaUpw/eBi8YkDmWKlId52YNfpQ5lU9b3Lrtw7taQ5ZKsnukwpZ7/3+XW
SPXQptT6eMF+4PXARwezvCeM+YzVchLcRijVWoWef39bvwtTJM+jyxd68A/KUROd
roYh7dNHlgGTGJgEOy3KE0aTXtsOZ8rvCquT6i8lYIA1jcAkDw0+kQ7ywQiHwsHO
QrNFlfi7SFpRlK0pO+QyhIrQsjNCEiUsMMHuAdL+lo2KgO92dNa9J3uA5J3KZSUX
C4yaKeHEf/pwD7X8Xz/nCKZzGZccIEFnLg66h+GmINNaOr80UJYeFFRiuqXiNN93
863EErqKQi0zWKO/oT0cEVnWBzuK9grApTN22VDpyb0utWsX8k3/4uwz77v7gYcS
67VkBhktVRjomNz9oF58AYsLZZYG1Wk7ixtKGVnveVH6Xt8lDF7cHn0Xz8Snedhl
ynXz9in79FZKVsobUEaNGtcLqYd7VL76IwDDvJBOvhnqcimnS5vMxBUAsY0ZfABI
/F+IYu84OMXhYcKA4teMGdWIomOPXnlc6L+MBuO4ScbQPqF41/9XeDD04Z1uzNRN
1xKR5KuFWLCkOFQWfVsl41CheAfNAc9cGis3ekUKTjQNiSt7e886SRSSVzBeou3w
UqjR5KvsdtoWBj+P3vvmFQ0lCaSxM0D7EMsIyCs9GxIV+OphMk9TZ94Jxm5JhqzG
yeb8a6vP/hKwNYa5KOx2olVO3QoXMzinGqKnYlc5W0lRH2a9uQuIG+jdDusx4raq
+KUuivc35MInst2QXBQhlTKPSdLtiLCt/JJbCSlaJyi87xgUKjmJyT2bi/AyNU0j
HSD/SUAUHSrRfP+WpIfmJjCRubgKBp3+d/r95RcGSKwFmH/87WPcQHolDecQZ3Gv
ho2qMKqa1l9CHdEIfevjTOU85fzgzUzvIvKL0zZrwWqnZD893ft9OrGCNZnAjUgJ
TvB5nF4Ysu9mv2fvmuKK73XLv/pvk8bRp6puqKRBJA3TPbMSj9VPkiBI0aBLfbSw
tY37HTbM18yRGkNF02vIzPMTipiLOdoS77z77+6Pp9Euvfx8NF5pTHSm28JuyUtH
bVwXyEMM+gPm3eBUDVfkMndzSykMTrKCuTIQqpCqPyWs01ROd/J8Z+CkX2xbsKhd
bMI8C5fYQM4zZKenzVs6wNo3ed7OIxXNDIMP4dIRterVqb87tGEU1bwSi3jOMC+z
Yj9aXqIGNMPbgJ2Vq3vVj7YlTDOKK5QkYhCd5cX2eVQZHce+lsKhOl2uuVkl+85x
Uq76jDKvZzDg/qCOLRgRjkxzg2/mmMdx87jEyEX3ayWv3CT0wYfThrAUN4k2TAfA
jazRSVvKwvwlte/Yriu+ET+8KGfteODW8RMa9lXXAUU6SphSt6kl0t280XCVjONS
HKzv0YYzmV5zVW8gZXug2OHbWqY6OI1FSmDhTbUVyXwDXyBkT0PPt6vDd5iVn9n5
p7nuXAxj3V+4GYua6kfVn6RIYWVFNZT/oIwQcU0tmv4Fh+IRXxjJ3UXZMvS85hfw
YeQUWr8lp9RTJxoJMEOOqp4/rZezIMSbLDxjHWp3jkRNoBowdIcvV3rTE7zzV8tj
C354p/56Z5yntihwoky1fNquY4DbDcw0eB9TQMKNrykR0EfLHuERg20F4iggneZe
HZEpIvUbRciL5EuuTgaysbOjPPDfZhClKGopxXJiAgsYR7+4/tEDA3k0BoacY/tV
zC/mbgebO2UyOlbSDQzVp+jcdU0em82lVP/GYdfXYIYGeVKqYxlYe7e65UOiAWOR
PoTK+3m/BgVmIyU+cliWpbM4+1mbpf2aIk6V9Ri7mE27WyXUPDOBdp42ANMP6Lmc
6p+zksTBamBDe45t1QQWlhJzc27LRTZCnkFkBEbogbKsxhLHwe94Wv43MLh+g36b
1gDHHW86P3cUCaK3B1X+MJ0z6Du1nvipkNeZS4MKzJ2XmsR3Kc6+oW9VzaS4VP8U
Gf4u1fXgoV4kFXQnfuO2AAmTpTaiwl0t1QCuNYRy0mIFQqLOI2WI4G11kP/uMdKc
JI7w6BNu/ypXVXhfWx5Nt7ue0S6paoybk3yA4WY3/XDuniXbTuRoaKQ9ACvfheSW
0KdqX5jllFzCfNJ1erRQliCTaOTKA0vD8o1pdtt+wc7bRgb/Lz5pKU7XEieTDi7C
OyztHiZGCWYs/T0+heAvVRp7sHB4+3bc+zKBppankbI3WlilVHqN3nHyLRM2E6P0
SjB/QC0Uu6H+hVIluUBoJSAS21193o2I/pUhiqZCkbmqdAjssuXsr8C58wHrSZBI
ormqsb5rSqFUSKfDSI3S1T8cCMPWpx7W4soKeg4VLXmya1ehW68veWZUkocdZCBD
F7XWrgPSTxKYqDR5W0CH66m+sZ17yMVKvQy/a/OuJtLnjX+CfNUYCx6LWTEk9exl
Q8XjKFfXCnqmQz8syuAGkrS4wKxCrz3W+MYWDdIv5B/66pnHurjTKwFTqvjVwW75
4S5wix7kfkwdqjklL89il0JQRcYkmz8+eQuAzFvwfKZitzAdRoGBKqa/I7ZdVeST
7A/3HMEchV37dcmLfbCdG7WJ/5YOOu8bzY0xNtiZGUd7s9sbEXqJVmA6t4fBV2Bs
1+FjgAtwxtpakQg5WrBYoct1MliwWScnDtI253NCjr2dafPAp9bUYuDFhqqknxl9
d3ZLtzS0fPaTafp7y4b7avEJVJ+ZnXJ+ia1zGc9Ilp+JxaTG65MjowLXsRUn+koZ
o/WleDtBZrIVbffbHseR+T5msmKQvZPMg78Lw2qqYNHxsTFL4aN1UYxS98bALlkc
JjEoWCnV5z4loDH2FNqvNYPX3NdpOcmfTEehJ4Go7chS6LlaIZjzd6EYeBgRqFI2
VItBGPns0dVxVMxhZW2nrH0vq72wcnmRe5hYWR6oQ22o/CPldhHJjZfQrJYeBUvi
CTaA5jKzK9hU2/3TJp1me9fB0P9OkX6tcERGmuy+X5wMnAn1AfZ1xb23xTwsJB9J
iB8KJExg5ZVVkp+Fi1iBoPq9rgr265vFVyQYZoW6L6bG5p+eKGA3w8ohugQHodCe
sHwRvw+StyFMbDUwJJHgXjJiRMEWyme+3T6GUlRs/OGWZRmwYDw/Ag91SCv7wC5H
L1i7EnfqFlOx1t6cjhjrroH9+mL+ReVNVWNZJLMzS1N0QWfIy9W5ALwHmy4P0gyW
wpkZaBxVL+PTAUewL7pB8ECQM+aQrqEzB9R7GJDfv2JPU7gzizgEyfsJx7Vfkcov
CXfGI+8Oqmv+LPhV96THJ8HJ5al+0ARb3EaKKSPeiqsq2FV5K6IboWv2+8RNokYR
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QNeaK+CVWtQsUA+OAUpwyjPiT/7QOCg3HdMc7KwlbpPsHjyKIHxtQ9LMgCGcZqd
CJpfzx+pWcylNYnxpaCDQTdbZ1NNuIPFZx26pOPWzmEfl6LjaPSLwo0m4Rg01TqQ
xfXA9jpAE+IemIS+EZ25/87zYnXEuGs/CAaEM+NEeNA+BAcIC732LVu+U0q/2hDj
poJu+gxN4W9y4wIEk7h050MYKCAW/tnVpHQ18PSM2LPo7mro/A+XLbOFJavJoR6P
h9O3NU0/xw9T8B9ZbLFq4aNmym+0bpnEAd1UfwwDtKMlRaBd1sdr6Kv7jpQmlgVo
agbA0Ll12yBON4xibZRn2M6vFIIHYGNcD1CDeKs5TZfORHNkvT/Qsg23RNkyUtnz
nHlnldpGAzX+vpiV4ARKOGF+H6K1+Ez5coGeYUg0LT5LNLQUdCqfrLUa9kFmwqXV
y3ssSAXQo0eJD6Rjz/wlQS6kyo8mvDkJ5S1ulk4YTOUucMSs0MtDgIsANmXvS9L2
WWTMtvZ/G1mgU0Pj//RkxRof+FWSEoi8RDq0yeIxi+4+i2LtBFRUITvhDGsR2+iv
8sE/UyDLGdY233t3IztNS9W7T8z1nOaS692ZBA6HyNKPHsguThgvkY4I4kialN4D
Onz328yHWVs9OkEQUNA2Sqd3tnc7wyOA9AUzrxVjC/8EvAJ2NLAD6OjTQJggMoef
MrPc9d8i3+lmzw4TdufufLv1YNTbdn7W2aCC9clnQCnmSloVdJYANYyyorI7LQ7m
lj9Gu3+kvDx8iZemrixiCqlegEuB2tJxPE4PAzAPHLJzv+ntnPXA65qhI4MympZF
9Qy/DXDnqGwhLRonFAXNbqvTcgFmUujJbjYi9mGGO9l/Y/vgggYo/Hv/HNz0Tqwv
ihXYbofq8FlCijillBmQZhk3+UWZRPFY071vQSKqHWc6w+4MNYBMm9a4kEg/erAr
TGwrQl9HwN46zTePCproE3bC3nW1ixxmw5GdIJXelpIwpXQ63N90qpV9rPPD1uOE
lkw+w7BapdEl6m81MTTxOCEfiX3sIQ8TDTP8XGKakmchHlRLNLCTUqQQs/8m2vG1
LgO1ePYQosKEeZuJiFHwiBMRYbO6dIClTPm+EigEDNQYa6GpjyIkNP0kVURNTYH/
+9ZHwbsAGni1E9x/oLVlU5PdWO/OX2PJPCAlmryLysBCir6giqbDJMIStzllPNsh
4bb+xQe7hInGp+PdWbsgjV82VzAAaOpOSLte4ySdA7Ud98iiDfbZLMJeYPRJENt+
d+9nkugAtWuLP35lEJ/nNO6IdklHiBwP7WGDjCvdDh7gBy57MffyE+PZT/nsBnj8
rsLHixWzcVhMiTa7XpL653Q3YhQrSNvNE0Z1rDjEv0+/LBb8fHImNq4WYY0k20p4
8X3/o+Y66x9hfWZt1XmC5FhAtpF9RqIahjRIdBAO/2XZbg0yFVNCWttgWVYr4AFQ
aNPr0IhHYKT/umlovAbfAjOE1FbVVSDZEw/R8vpf2FFNAKsSlRnE/NEWBEsQsYSr
ol1S/eveqF3soZ0yYd5Nf0HWwQDqjRiVH6sdHea+p411V/NgcVHUKTiXsPGhaiTn
Y6X6LEwbgFRULQlRt4dguukSGycu3T5k8KpQvQl22REwOFGrZ8NoSmnDhXRs+C8W
NeMaR7jVSoomIBQWxIKwuXxxGQAE+deVz7daz40XdDfc8UQKZilkhsXS1+msQ7F0
B3QJ5viYEVlMMNGTYxyZe4sf4m2GmSGcJixggAs0xGThRkrMl5Ovt+yWAa5ZOOK9
Q/Ix5QpAeNbYNxvPLo7XzcqdKB6ACJmt32w8w67ocel+sN5f2r/u6xOYp7jS+43G
swLMi7GnafOwpM4p7jEnMXsoCwo0QkNpwKEBboWVKM0rhkaCekAPZvjRpIudXInA
B15ZquTNvg51cwAI4oq2LCE1grKSlpI7DQytvFO5ns5Rr3ElfeU0UaFAW0KWODpI
bQZJwUIORoDwBhc990SxqzElda0mhDbmA6aFx33i0icfBz+Zw7OXSx2jgQK/vR/v
e51PuQc7U4N9xDxMdPGhPbEvAVQBoQjXroagwFdHkY2zfWJ5W6EfEv7swWKW5mJA
Sbui1IxgNiqk7HMcJhvy2YKOhJnYR8wkqyhBiZ1Nsqlc13LLzabL+epsQXZPU/oo
Mnsf+oZkh380itySHr3d5GRw0NgnDFAXaH8qWjoBPusymT0GWg7AH9QOXr4KmJ4d
tLNQ/CfkOFIuQuZaL89j1soGk/OOwk1KkXiQs8813q1KjfTce0LN/sUPu1NZrXSm
Oap7Rlg+SYdv7gCaHdufb1zSV9jxICQ/TgedFe7XtuD0qr5JnvKymZ8NHZ31f7JM
P7CmfVuwu4MjseF8fdr2KKTYZKWIr0LfBHCoz/gR/+pR435rjukM3xtbS822FJ9B
W8K/Zg2StNc1yB2CnoBnkJemrUB2dwi1K9ubgF7zZgoaquaYeMNwv83mLVBupPb/
gq8/Vw1BFaqvme/+M1bWT6CrYG95JoYrX19kKJ/kNbIqs25SdBKYDyAp+pCvY5pC
qt+xKRpycmM1PfWgalieDm1cYtATQgEWWyNNHUUNSC4BPj8PsL+M6+q15KxvCWRY
FJ7JZjrQl0H5H6V+a+AvMEgVOITVxU+FyCmmjMNcGDuaqFkPbohft/sqHZ5Lv5V7
goD7uyXSKmds6dkzUltIr7PsPaqltO0OIKqj9XkxO4lRvqYwAPz5KRwMRhkAZxbo
glYmblpX5jCUU1MgK05+h3q1b2F3D9wsE7OVfDcDZOwiimv3CE+oQf5ym7EUg5yZ
WbhvE3MZhhEL33rTSGE1YLorU6SoEgzgHFBnSoFSRFliWObFZDrrXhD1VGIfsN0k
mPyTjE7pQc8uuZQhRiVvMVczTCtsMYNfSVwaSzhrWe9HsIbW4xa4IZX42PFWBfK3
ETKJmIvgHmJ/WSzFktx/zetjfPrQ9kVYd3vE04m+9B5x3YbeYGI65gGEbKZjFL2G
oVSKgykuaSD8Qiw6dD2t9UmBoUtt0oLn3PDQt0PDh0eXIO8B8kfTYw/q7wXtbP34
YSE9dhZGB99ru6KBgvJqo5ssVCzNwcKGI8/v4BY1gtiVO8w8wgB8Qfs2HoCeghQW
giLhpHMD07VRD/HVlogEbEiuf3v2Od4KlQYqDHZSvDADBVGAXtDvI5R8+ZcyFTWv
hHwz6AjX+VbmV4tToQtiwfKGjd4Ut3yXcbuF6R1L/vZBS2TL1jRa78gJKH6/D84k
cI1nHZ5hkbAupNMmkWc7wJWlhaOxGD2MCTufresMXAk6plJtnXGZ/Ph0NqE99f5i
I7MUya3f6ilQkNfYI2MBGWMUqFvgyXttagmj/mBFnx3u9fjCnIVWQzb7+Zi92LuD
URWYxa3OvVtCBqUIPv5rrU3LtqotQw6HRetdtMZQWKfd7U+y6h89rbdzhT1plZRM
uso7+mIUlwPjsy6DtWyVUpAeKgFV7YTrIrawJlAReu2OuKOkjZzc36KVPBGckfgs
tuB1b/x8m5EQupNBfz4xZ7u8SAiPDR8aG6apxAol8ZIy+D6jTECgsbKOW8luj0Xo
IxJL/DSikEe9PWXDgKHVc0hKGiS8fLvWZ1EPv3/Knt+eOl/DtY+Nuq4LGxpkIv9P
bJpHO/4bWUmhzStbVOIItUtqIjWRddcbkiPRG6L2W8p0M2NqAxgXGGc5RtTeJK52
99g/yCJRjLDcekLoczOVllCnRMW4D1jGGhUhrcNwFucPcZXspumhGEyqzDoyiv4J
MyBO3MENVPqwaRtajvWiGkBxFCbuARoP9OPCSuzVIzGYjlMrC1Jvm7WGLtiBAh+c
ZjlDH9695qxuS2hJBs8hfi4lDKwlOMfJSkKXcQa+WGERmWRJFleq4LloUlu6Mcr4
DcIKV28AfxyP36V7a1PUWHY5H9dR5JR1N5OothL5CpxBUTbSBm8AvD959F5RNlLV
RWH3RLdHND35322nxwGggY4irVQpn+2oUECIJhmOFa28v7kFhdNh1JnGaBE/Z9g9
YPiNLoTL0wgt73ivtkqhmOq/nzxhBUw76yprPd9BgsHu3vf5ErrzRC3NseSY4EZA
ISqnNY+F8qyF5vSfga5pIvw0iSfPVb1loHunukMLtpIyHvQZY6V26HLwfio+toe8
/eIWaXyaj8bDBkxeJiFp9R/fVJL3mZRIJPC3+MBP+jdruQQWe7U4uR1MGaD3x9fg
K/tBpQG6KUcMbmh2ZXGHU8dz0sWrTkJMj/JRESzeIA83Q1DlesOsxWRGSAUJ2fkP
anBdLGJwQAOrqg6lhz+05tKuH+YUUaNMVmYSWtuC8qVfDmRTpxuLeERufOG8UQsf
/umhZZFdIjE4DzitHzfd4umLm4axOwp9GXZeJAdFqZyQcdFBKHYENr9OkE2g/6xQ
A+LKmKbRvIJcDrVLG65jAbr6y4WSie2hx/g5X8bZfrlkKR11liM6SsZq1sxS77fM
PWiDY5DFr7Q9up1TZSazqmnULLy89+JVF5k4hnwQ9c5jYbe0WEZwsJxMlh1rgJ2q
+qkzXZHWL9CDfSlIFo8E5xx16O/99wZ7BiLNJZTwrdi93YEPuChsX3pwTVgRI7fC
IiP1PXdGF9mgtXBIMzq2fuxJpeteZLKEvUrDHZ4EAuFl/gbxntzB3Cxk1jz4skEq
NW0hl/S3RlTp0YZ4fJThn8qoQ5wmtzAymOZQdLy+fi9Q3luuLSHMhb+DIVld5fL4
+LsG5mSqGO7tx/LbAgfDEcGIRhdm1ssnTYr4D17I+pCXMDrQtkRkOADEWHV4d8m0
6DKj0dmWTXrb0hDiMoWEicQGL1ouIWVVAfktaQ4LsN98y47LxF/HpI0vOjzNKxqz
gfbdOlWq0qrp75pf5dfqtBQXx7TsjfGrBWFkNUUiUjOTidOCOGP0zh5FFW5cm8g2
BsNmp7ttt0y5XrOTtYUbC7MXCIFAYxNyLvbb7Ps9WPa9cUh+hZE5zV9ZC5rVhf7B
X4NKgeJzsXD70tKD7Ga/7THxeqnHKn9nd2Pw1PquU5g4phdrrRkZ+ZXkRL5FdiqF
r8TmVyngeOUh0GxsLwgJtuvaUUmipWbZBan1+FtkwAQAixyqh0QL8P6DBQn9Iis2
rPTYIMB+e9U2Bfs61x209dmEzzSsPE69adQrLfAfTR3VuI3RfzZLAf7w0fDGz92d
NPBBMMNYSDlES5i34jyMWc7mu44MW7ZB+A2UU+edx7BExcVLoFnb1qDNRLgzIlEH
wg78K58JFewZwm+gyjtlBADjdHA7kCap+wLtn6TNPQY8C5UQR/F8L6VH/pdUWVOK
yD4mu1CVqr91n+Ph7hH3jjC1MqrQjjYM/g4CSl+j0kKVVOAVCxxQQyNB6qscVBIJ
/PrtXNnwbywrfCfk30qxPQxze1l8PlkiMzMb9Ykl8jZoo9Vflcfs0OTIbHuvS7r2
oLbNl/6zqyfB1PqMMsHpip02wZfGjVTG+nlTnerAXy9fuK76YSE6wlu+4Tdy+qGl
xmnmcHcdxs8xTR9zIG2hNv439R9X46DgKNygJwltRACLdHVOgTPEbWb0kOYmqd3o
19o98iyIaOOCWP0M9DdkrIAB/Zd5lLREh6SPIJfvn0JznL5CnlzyvhSOtxHsCvHg
SNLFfFiIG69f3PgaMsOOMExtoDZ8d/cW8fOkMKEq9VboIfTcidXp5L6KVdo3QIkp
cfWUxtYlyQB/kppDcNSMiY32qQglSMVg0/yMxw+GBMD7D1HdXfSOcKMQX4E5yst5
lbNc6QWS5FxmZfjiddrCgiR3s+lnjGiSo5JpkYvEWpRAcDKzuwxhFnXtrhwcsIxF
B7XEH2jyKUxLmMN6tNtkUV5KGZ/tiNHXS7qoL1u7SATKWnZ9ErxhJ7qo8FGDdi2r
dlgr2I3b+Yo4kz5OexJW994Tt0OnJJlaU0H0ytKw+5e2jx19WdmWX58R99vxTkcT
NO3OGwCk5Z+2KmMbv1fOfFs/WCMdB+qFx7I0ZPdkniacqz38HcKct9kPGVPrE/ml
gz2b7oA4NUnX+vdw9ZN2r//sJhFelAof/+xITn1dbWcrcJZuZWhbmw0Y36vWxtf1
bhyxIN4vjiSxXHSKW9DhPy4b5RcSVoN3624Dghar3DtkkbPFoyiqE6c2w45tUjbD
yZ3aUfYiiQ8FVrHiMVUd8su865cBne9Xr2AKLSKzXEkFzj2VFJR/+uR/vjaqUT7J
mQPxBEu6x0vwsgKmSnR5ouah40dw4rPN8RNX2305EJSqkq+2t8JZjGHQyyXL084x
G+E+1TDTjjCBQ0eKqEUTV6am+vlfzyaIm7WfnBLAnOJuI0OCJ9ORExnE9H8vONuy
2IxPOhy0pttsIZhcg01cqnqYOLhuissN0bDb5ESnMUKtUZOGWucklW+W5G72mlyH
sugirdLj2jH5hzAqVqef6roU6jN3DXZS/YNrm5ckRZ433FBdvhi1mHLvL7V24aaR
VNU+7QQAsujf6ZIBRH6PSE7UjGAziXsaXMsEGDNWJLoW/CmIrldSKF54VS3XFsQW
R+jtOEGcnF2ST0l3CZP3ck3q7MDkjih5IUEwKLZ2kIimtAGiGG5iKjsjgTH/msSu
EJjIbMnTZVHbcTuEDrFPFfOPw4w7uuIN1UiQZV69KiBm3XEeacVX9lVyYab44cfA
gljVKzmurlwDXxkQ1xI6AeLenmAjZyJnDdH0NzEPE4fcT2aXgA5lYuHfbijCs1eO
g0jsEUYFzuRLpGRQ5xvbOYTDs3/9rNmf34uVedBdYI4LfN/BVlwwgwxE+ZN/1VN5
wclmhRlKEx8wcHF7Pa9DMg2he6KwPQx7AAChhdg/XOx+ZoL/ZXyurDfnH0wSdXK0
7kUS63QoESnCtYW7Zjj+TXwzvoCaffkGVBSlnxg1TWZk/KK2icc3ay7s7iVYU/k/
50Qtru2+5uL+roP5fXPhNqt+j2IgVJYSoQzSYFB7QBG0R5CuMZLy+A09btXr3RLY
pim9XeFW/hprE+k+hBNdjVpyC5EO7w0OBbYZNP9buv85oNUJISnnjZazUbyYpDV7
PjYlERw/j4hfQhzht+M7ZKRPIdPK2oQ8utN8mtfcdgrLIJnTMC128dmHuRnnZJh1
3NArZSL+T+Wo9Ur1yubloQFQuSMoBA3WHPKZAEB2aL7wive8XD2AVjgINczbViyx
1hiEq1j+kTRPta+ZUy89UKKjNLrP602AdAc3y14MqiM7C4/ZMHy+woGDxlv8KBAs
l79r9Fk+OcSCTjFTHo+00XztJ7Yrrtquounn41wWfPWelV+WwYVw86J38oDNQlrk
hNEOpbhzODJFUIEw/QXJdJIW1NOFA7eAWXggIyP7JWUl4UXF6gavTYhh/UiOyG7Z
xdUsK67YL1XmyH91JSADeXOEcwoCVzmccM7ubugj3XsXg0bAgqNvWc+mSkRy1dwC
V3dZcPqV1CW5h7BP2Nndtn62HpwWB1g8U/XMIG+nX9W2U+F4maB1aYZF91UZmkgq
c4HXHnviQzPMvJKvyOR9DMacZxRmgoDSGJJTjdknqodsUm/Uu5A9vWJLhSLw7bYi
AMJb0MinOT1JQo3w7y0H68DkUKS87mrF0D4uzYeDXkJxrq3yIYadJlUlRCMZ71kP
6iijNE+9i4EkoSmTj7MeXI//M41vNJPPbQ7CneyFcGyDVb6InsBsFOB4NxoVCwvF
5W2yfHfFDl2swgz0XVUW3dvfvWEWS6nmx0IMFjSqcJhMy6Hi/TSi2B3VYps3nzci
aphQt893106wz3wlwo68rBs0ny6jFFygP8KmkhgZMBYXsVzAReeoY7tLZL27gG6O
/Hq1Urke9qzHM6QmJSCXQ+5rSFEHxlOKQ4X07zHd5kbQvqVR1m8W+TozhiBERwsP
H7rz0kc7ryJk2DaZvBmYZa9y0qGtrdLSo3URKpDQ+NxsaVGVTUM4vNYSQsmufBXG
5hccPfCK4LVMxkVlKOwlUn/DN/qUqVFR9FP+SFyI+vAqRG+i9jqgdn6FXPGyGeB/
YLlSDWtMEncFIQG+Q24+Xi9RhSklJVAPPqaM43OZAf5gVSXX9GXp+eeHZMH0kbgF
LdSOWTwmo+tqr5ueZ+N5dnmUz/VQBeINkgUPlwAYll5hpJfeVO5OtEVWu3dDRep8
XXGMMdQnUf0l2T4OgKOvqKJiWbT/pf78VOV8tdqR6nqpZ6+ep5YGlkWUHXiAp7n/
G7ir03VeAczZhycX8r8N0ornvw5loKizIDFiGaMnamJagjQV9/YwR9vtB0et0Q/x
5hbixQHSeCrn1FxB5ldBqfuPKgx09RSkdNwnjYHsbLDp9lyx5ukbngpob+pODHhb
b8vxco9xXI3clc6JlwhbQlooUrpvX070R7BznFQ9QXtM1wV/kjKJXho96qIP9CLW
QEXRet/d5pVhL3NTzx2Us/IUEVleQgUemaIqeVbKiwRwYzVCj2/8MtcKNgXrqjnU
cjk7VuRufRUzyU5++qCqZrUC/A+S7atBymwiH8xnah9pXBhMTels9FEuP4w7gBBb
lLFc3OrpR0ZlLB7yXPu4Rb84aMmRYx/6Tfo9BWlKegwuaYhdK8pt9mm/vOR3l80Z
QdyoM9fWwXngzSkwWnD0npi7ZGPCEchDY0sAx4OqO6/HMqaqrhGtpTGtn1TDCfh0
ecvmn1qrMrSm/1ZGbAq36v51Em+rP+EejTvvrhWn/HqBy8BFii1py9JXhqkyAYum
itEiI2om43Sj0LoCqok3ft2FZHgnINZT4FqqIElb2bsIXJoeUvxIVEd+kFxaOkK0
1dyPK4IZBog82eRZW7jxcXXNS01Bfjd2fBdHcyevu+H9dprb1jgQUn/QaKMYqdWO
gW7aPEl2OSPXzPcMBHMC32imVO7fvYdi0Nkgfe5RqOGAG0CqCtlDrOCsHUQaytNi
2blKRVDzhrYby6y9NjYJefyPhVWstNlKP6d/rDfAwyk7XApX887xf2jI1P3+9H5D
KMsf42f0+1xxI1i2HkhVLMtbrjNLvyUOQ5kSwVmpIN8p4YuaqUbuLn5rqV4y9Kb6
KEeTBZebEqk+QBOR4VwL2lpQ46XcVjZCkkFrGFuszPgX0oXRAL+qHdoJAzwd2Adn
Scihk3S0A9AsHSCSqAMxcT7f2pDtqzQdlUiKKw0nXMMkUPqaF4eG1g4plO4fHWI8
DpnpuBau3aMDSrPR760ZYITaR9poTgyhdDofH6Hx/7An0maxnYFjlPQJaqUESeI/
n6pjUYqN6zeCllEp0KZ4atqBRKYRYuJOFRiMRqXeMWWSkNYDePKxdfjKTSEu5TPF
U2lmYbEGenNVk+BNd9gvprN1/6VchBqyBeXk3acTPLC1qo6QZEiHFUNmbcemMb2T
UCHPn02iVMefA++VeGJd8/mxml+9QgO3o+wcQiriknBwszyUqqG1M4bRNG5IHRBz
jSpX+JH7Mube+mq4NOTmYZeBe32IVVO0GyEI9YYdht3CF1gPXtouQXgzT8J+7xNV
+D8Kj85maFinM8np8DZ58CTrQ9+xWZuJjX+bwqBYPrLrnpePbnh8mq01vvBna/gF
jKR/ZsfRK4u/UR5x5w66ck3oxXMfBtpwK1QC1vl1ZX22MMnm+XsqX64HVWZ/Ki/M
jrSzpcm0eUANQcTY7VcZh894TybBKwh/PU9fR+r/LsHGlRX35wh5fJFFUAPWRakl
Tj9rib4nPs74fhDj6AoLRQMqZODvogekEs3S8G3ScEi/02bPeO0UsqRBzJY489nq
/1jDT0UqrCCCg3HG7GH3e54pkAB/1GBj1URNyhhwsdMCiQTiuCIGqRNKlThi7BkX
WCB7+Y2qo4bttv/6jiDBAaZXUpBWqrt6WT4AyNhzQXC7D5VkjUYcNThcAl5btXL4
Z7XCvxWbUWajycG0AkBDx5RpTUy+eHqQeCva+1kIT95QvnOVkeZnlWdKRkmUUQlK
Xyzjl24qIzBKakDFxdB44uAZOaKQRf4eyB6HzJQPLZOGAdgV4GuwBryCkHMgPG5U
De9qbs+42OPFZtVpCFQnGAMCpeu7w5SiwO6WRzTa4GgZggPR8FhLzPLzl18a1WtU
yg4LQI0nalES+Yd5KrqEG+orX7o9gLmgVAcKXKaWzqFO8FjlA7lUnyhmvVw3U0Dd
xc793UV2gtsHfsC3TZMUaUELm8r4ztJsUpPVGSs2HqHxqAA3ebZaH1PZC1qopk3P
5uul8oUW7dAHbodUsYfM5Ze8jPsykfIyKKxN2KstenX7RmCO9gapD25PstQxYGId
iGSIH3Zk4TivBG41/1z5sriJ2meE0x/9T5SGmICGGT1FkUbCqS5WDsykJfV4fr5o
2W8cFsOnRW9XTFCyxRDlu+TTL2dHUmOpRlKFFtiRH7hcWiRgr+06mcg1QNYCP5hG
3JsoGuG+a/3lu9gJsYUYZ5cb01B8mS6CRxgLui3M7/TIzXIJtpyn5SQRCetIAyTo
GIQbQa5ffyDqICwwFQ7+ZHd5xYNDMFWYdUzF9/1PLhYdPSAhMbvlmm9v6lNKLZts
/wl6fJ3gKQsq+J2gUbWWBc4VYFTETrtHZiH+icPKbsNJOJMCnN4VJBuVwiKqngN1
CMlDbgy9ZZszWWZKst/1aNGbCEltL/iVirvRAgbrix6ptu7DPNFLK0AuUkWI7/gc
i1F50DhQ8XDa5R10WlAIRq/JZA2TLhxzdOLLDYTIbkTUNKr+0UBzztzlmONxeAch
oXoHGrmRSdNRe2hD/xeZRiGPFzeqhTC7RQOWDPk88GxcQGChmZYjVH8qTbY6BG79
y6P2VIZP1AnzMKnUDTYti2iOb0JmMC/eYsypUKKb8q6AjKZQyZp9WVcVDY4Ad4KT
wCRLmyfKa82bek4fjhEFRG86ycMkug3O3pejeJHfmK67GNBxiVjOuypO+PZlqDUq
nRKj2nRNVd9iXI53ok/GTVoxav4ilwZBxMRjRD6Gc+lHMFxmUaftes338QqWYNh5
hHpsWu/cdV9Lg4WCMGQS6hJeSBZFabDU/9av1fkHDChOZblgi7614602WnXgQj7Z
HC1VgZEjp+GKbZ6Rcu7lzdr7XatO08mAcF93btiXBynWjh+x9zqowb4MaHXZn6zF
Adg732OyuIKP0CWGc9honiQhm2nGm6UJP47yJH9PoYqmr+PeunOaCr1LO+tdMTlH
il1VIHXUq+ZDafdTdcoTNe4iwV9UFTtcNl5bCidezjau4vwnXK5DnjimnO7+deCV
vGR2L+z+KGtBDjtY9XAwy0wBtXP8ZASyzte1LZB97L9V8iYkYEeLmbgiRAPcw2vK
2kIhRB3egBHVAlVDAzq3oSA9o7tKjzBDBX1TIk6IjAD1btd2zYkaeTWkOm6YxoQl
znyBGHeboWCaXI0JvoRoWh/0vGClm/+0EJNQdIeBAePas23Tb77yDI/jYuwbCZz0
doTIQaB9AFK47bJVj3HbAaAL6srUetJKJSwGuJ3ybwFheNu0ZBZg9am95vWIGYCF
hVw0o/C+St1PqQ4RK5VYRq2duTDyGRge+csv7kX4WKYs1o5d5HqgV7ITZLVRjKSt
OMzVsAGm31DSD+VX9abcF03IEUBgQZWbVGlWWV5vKd4rlyL9Gjn7RqAzNqACdOKA
A9z3rYwguwy78Uyt7M2xEIO/Z0SXc923Kbs9BuTOgW3ohh2EL1sztMbqwMdILBFQ
ErqleS0/DtMDqZ+yGHRaI8dpNCnaG6/SpJ3Nh4QylyFEblYiV2rxjp5ULYmsM674
q15//YENMn661dBiFu8vn85GdrCMJw84RXJ0wD4JX2r8kqWUjn0DuVmfIIfEWFtq
KcneXLWIvwxFxjz3NWn0JFkZmQVTWLBoMRaRYHcPVJI3WH4UokajzXaqxTb5ZbgH
LxwEbZqY+5HbWdHa4/0o+HfmFMOuJsl4blpa2Ao03gEr0OFfgfZ4Kkjnnv3EgwhL
3HATky3WuUDav2Zh0NrvNzs7VpUZd81fiE+WohBZ2SseLtD2RTQKujQKSNx0Zd2Y
pqgtyD25BlslqvF2ikDSfKBsJCrhCLe8YlxPI17F539LskHFo1Gkka6K06eQSwlD
aU/Sf96/ScaWFNTOpNaf8Q+0wrNtZaWEbE6wr0ptydgDy1kyJHlwY1t0b6V5jrwo
n8gCIPgwWkYUgz4p+e2VRVtbMKcnHzeiJAmKQa4gOSOq/cT/OT+QuaXo1QXdgAgT
7xm2/ioPPtGUrpMRkln/I+51BuxbI8LkCD6q+RXzj8lOSHd9OKuIiqMfpQ153zUm
HFmmThNAiOfwE920xxWkV7T5UV5Ngolmq/Op+Bey3NdesjsN7H3EH2ZC7PprVYHy
QU7l1c4EartrswueuSrKvXIfPTVE0c2qo5s9yKzyzeocUaPNAZ/b337xnlh3s4s2
tc880m4lkHB7hJFjl8mlskz64rf0cJNUf/TIibmspeepTTkZeKyPr4m20N3Xku9M
2YAqcMpKr1BMSgUj3JMP5FjY0ar2BbqntahM6epUPFPq3x/qW1rGG2Sq4vSz8Z7c
kcShw3vqFQibClVaIq4U3VqIgCClWqOp5UImYp3HDRL/+ZQlto8H+An1HbOLIEDQ
Ozp7Kwif/5/tbef7Jgl+1HEfuzlDjGZmNY2n3BFZ9dQa+R6FJK/7hlv5I4xlFzON
I5mkgcINsTjJNf2o9sQax7eSzIZZUD3N+hwaaI/WDnPqtCtc7AoFVFfLkL5Xz3pp
DESACOib4NIHNTeJpMB2EaKLAk0yGeRPa02DXPha4JJaFDgGkxac0nX7PqP0Os6Y
+ZvHyOrm4PQQnfogvyeZ+LMKgCP562FTlXzAG3GY0YbjVPqdZFA6DCdi2yA3PsU5
btbWXb8Be6sz3E7ZD8qb0AuFKHwh0DfEFpabrHODmnmskMaC1/H2VPhTwCMNboRR
UslwOD+CHrS6QMIUHjoDZ/L4Q5m5GAbUuHdxblaE1Bb9M09rRofdtsMG+YcrQ43/
r+Y1bCrby8fnX0KHhAb/bH4A7dT20lrNgacb/ouMUZfVj6Tdvb06f/S1qKB6W4UD
pQSFEbKg3hyiw0ASbK6MbhO8xF5ACu6qZoVNpQq/qaFBS4qYFIE9NvwUY6KDap2u
pVXylTXYR+Kwzc8RxOOVrTJ9EL68AtT+zKGIPiY2Y+/4fbVDinpMyE1Jx7tLkyv2
udaOcrc7UC8/9myBXllgt2DBBOutsR1d3fM1+UjReH12T1R0h1BEh/kJ4MGLaZUm
0boj2DZAqow4oM1A3dl/Vn1Vktavz5mdMU5sdrU3F/faClO/ROitytoiXkuQSabz
XkFb2y+gLLajBm7YxBdBs4jTe3SAu6YPp5/cq7xo7QTCGM1IF1YfSVKOxfXziJM2
fRizb/L0F26qPbbvCYV6vKI7yXiDIN5mZqLhBoZNzh8J63CPLVgA0PC4kw+u9Fyy
INU8XxPjzZZY0pwKi/FcjcJSj14l6yQk2cV5Rb1NtFBUZxMOQ9zAW9lUDWDv9MiA
Wvz6mavDhL/rMYUPy4YyqJaBpAA7YmYiaPV3vf7QRDTNFlDWGpIkhza2VD8jO2L0
rkRwvujeAseD+nQgS9J8EVxSEy5lhWzAz2gGo4Y8948n2TZ+cFsZfJXkd5cfu5GJ
4FcdFm94OUJHjoTPSCJ+Rj5xZFtBXHAhHFrVseddTldRlcXHY2rQFQ12yihSP6KQ
fpfPdOxakBwMEfPoRW/2EVPIRa7eCoVHO84JXndhBhK8piIiTPMuiLAORbpxznl3
GemNuTustp9BXq2+KgMj1wfGzCeP49+FDAgb927OvSoCI0VHxItZTBDoUMDMpw/5
HyzK1qz2aiUrCZi8I8EDilXpAjfBr5xy/0+kSaJ0T12Qyu8NoVCV3sDPLcFrfxzH
8OM94aaDNN6tdloqnt1/wtfTHvUVbchrtxfJZsjzemZbpCV5CWVDd9lLKNjQONiA
L0n/jzIBCXwXmHq2avkJbJXfUK87qE2GuCqNXcFMUTDKcaBsWq2qbbGubCWD/1tp
fg+UvPDh99rsuq0MYva+acDpdnMrNcEUqYI7vgvEbozKhnAgWFRZrn8cslpiu5Xp
+ojZafXipx//yo/8UXC4mduXLaJGTvuPJLpMzj/eo6p3VorpS9/STj9VBl6/B7HV
7TcPIivMxqEuAiUVKvXMtiCeKuedfCuZk1yvyi+tlT35gTVUR3diZWJQbDz01rIG
eR1ghZkM1cCk3BOueOM3X8XDR/rKlXU7puHlOC0g2OMAC87eaz/5jUxDJnIE1Vys
110L73uXXPt25zboRYzFYfYh6Kw4h69UkaRmKRMz8Kjvc+2eTRiIjPByjzyHzuvd
m51IrMVAaWVwNNdc0aZwtUlxOaK3EfaMhbZGCfic1leKSjx3l981q+1lMQHhT45g
CjGZVH+GNolboTFTyzkzk6ucO2hr3YsdXUQ/ogYKza/7PNL1qFIVfxuQZhWDH45V
I3cWQKz5hkJKfoloMc5DfN2iT9XO9xU1VSt44irKVaBZPl2hrTe6K8Id1h/kf6UP
62+PoeoOsZhHriOfs1Jjg754G4XrffUDVaWQl9iRBpZcqxWJ4O0jOmo6msWoRTKb
9vvA4WkMO2YpeM/8X9AV1O30yImMlNjZoZj/TEhdnGDKW6NNQHaBSOZzoKWLvlgo
W61lTB1pXbsTEpueiMakNIBqlbgR1dbIdWKdu3qgacfy+uJTlSy/VFDAtvuVGirF
8kgKMD7p95shqcFHaxtpDqBGJ3+M6MScZT00YZxPnMLQ84NQ3CIY88adMtqhxgHv
pURmpfacv0eTIqd0nGO4UarEETU5N318eF74g3GlVMkRHn8PQQS0mRLDpCZEfCd6
BehEh7RAVHMSLJ/5zuIJ1OWbYEgNYR8fzA5mp/LzKByLkN0vNhvfAqvN5YJGAkKy
MSnKzZ9iVKNwHGJByu82rflb8a9roDeX7oQnwvGVpd5olvNcWG98cjjA/sT3fSay
3MwzB1r3ZmngbujNl44suXLO5eD6aMafUEXBY32z5ivF1VytwKf8WvIVtIfcihYh
dBZwTH4o+7dI3TqhMAheX3yTTdlpcTFObds7U7v06ANRPe7zNzdbQPrgvcfhGCDQ
YdqKwVqBDqPgnkBj0gNTFkOOcGGnE2AwbXvTLb1opLiQKeBxtlPvbqJ2LHyZeTYC
m9e7YpEGPoEC+C3NQqWzxJbJFvOEPDUB4sZgu8M1hhg66QlN7hiQSfXz+xYL5ily
g4R9h7zEkM1hT/OLoxmasMF23clSlNkEPSSp3qV6W8ThTopgACEaqSu214BNjJyQ
AHCNv+VkeCvYgCxgumLKQXMK4nOLXv3VhEYqY9ZFoyQxPpfA+8Orx9QTBu/ZOVCe
+QH5zBtcimqwH3gwkbjFJJxs+WlGbXL5sqff69g+m8uUET/u+bACfhSVCFahLw57
gCjBFqQsp82DtgKOInw9jHf6Nf2XvHH4W5IpLn+NqHFk+m0opPKeanrcuHUe6vKw
YRMAEaXx0ZTTgM8/sxkod7A4G0bZAMbG10odLoz4jelFXrSJuZukIlOUW2HcWVaT
O3c9zuM9itxwnJVOzE8bqup/UYasd7LcqBD1yamQsW6URLxXMHJyAR/7jgw6e7Pf
LATb6tVwfvdQlrlYoxLI08gyNOTjXP9KgJvBUt7yfkFiXekSthHiiH7J3gYrgFOg
FdSE38cZ7FdKb6Lf8YWziE/lEVH3/IQE4GP00gxAc90t9Ep2foD+MLDit5nQhrHc
PLzcOQOwYIDW/gQMJGDZRV7ptP2aZSa78IVUOAAffCShiWZnvKNYEYKuCBpKRVGy
xeZ3OSKQYQJbpd/3JLvjLIb4Do++BEsQJVQIBXx3gzVkfyCJCvTmH7xj5C0TcSGH
pYmFWeBEpaPXVdIoEfWlJP8a3PH0ZYD+oqvsLWcHRKvzBNKtTA3o5bBP9QJZfCpQ
JQXUkWObdkkKRre0T4Drgnb714NDkE6SSoRLBLHgPyts8GRfg8BlkQ+j1KRBWkuZ
jLKbS5JvNTc9dzxVMzDb7iv7ibzKxxnb6ELb/GqJTuQNhrlayAk4GjQocNQSz8wv
hSx8JUq7YiHZwVQZKJmRrK3+2vw46CmmYgcUas926VaDbleBQhUXYyCyA1ELED8T
RhlGv5LaJLULmYjjVPYI/Sr42wewywAsjtB5vmwN8ekoNIFHZZvb6AiMhjynyvQo
zuU3nCcvwCS0MBztwGrtC8SJoa141UPKF/bAr4vbNsPyXr75AU1X9mRFNHCX1rqm
KKAnwni9BIr9T+NlXzbKpVXoaO0k361FQSJzoZQca/mI+tmitFbEZ9Zzn2SnNsZr
lwKGd/SfQ3WuAMpf2CTtisRdGcy032jq1qZ3ty0j2DDr6oCE+ro38+RHfzv5Cc79
kwQYeUQx5ukehj3RPn4NsxOJPXZxEXqYMqY2NZNTD0TvtOLSSCefun7a7o0hhBW3
s0zVghKWCBHQCajsPM8wKDVQyV0nf0k8y5gXz9+w8Uk0LeUFeLujZbF57scGXeRD
Ekk70YgUL9KRB+EEqyX/StRybHIM5hNz8nE3n5hnFSyupg9gy451/R9QwbTFYlfy
d9jABNYl2/RS4uyTzPy3cDLiV0pdFrcb9aRZDRpOOfsgHRZIVObZc36vrIJWKy7B
NMbQg5DILpi3g0SGkgegSjNKc5F4N5nICt6ebHZ+RO8x6OoejT8ksi6riZPbNRt6
AOglhaTeXqq7jiytEMkJMaBu1Frn9ZDr0Ryah0zzsTUm9GCLlNnbgZrEersJL6xb
U+r4De5TXRh/YQOj1/qWHQqUcI0N7rTaUG5TH/Rpmx/Ye/EKPRgb6DqWbK6vtJ6S
6Dyvcra9JpSsImExe+kZaGNa2z/4BgLocZbkUm7cTZgGBLPBsvy6ZTL7NmNBa0X2
A8afqtefLrJtyizSVVsaECoTLoKRRoUuobLPu6eI2b23e/AxqWTo3JA8816sYJc9
DbgtLeC0q0aiz8UM85zoH+Iat5XdLSUcwNmFWDHEBd9jLRqP66YMkvggGA9WLByl
cVMvaxJjwKiKFxuJXU9sKiYT030M1wF+74d+AXb8QW2AsyBFAw6ylU3/+TokNKEv
tQgtfYIOXgQCoD83SOHWKcstFu0WjhSOeyvnV6rFvM8sD0XPl7a59KxbzHhfLgKl
ge0lgaZofq+puFYWgpQuDgn7YYc+NE1LfAk5QToJfnFl5d3icMVUsIRWAtM859xG
WSnfGoQFuQJg4iyaRludIYdOgoyiifRuToPeStWRgrpDrIUxXxyStKvu9AowDj/l
wt0w7ugABoocWCuNIJSCiTrSDJb1z7dg7UgNjLYdO4qBjhMQx/BCvgguzk5wwGul
LvxfY0M4yAhGXufR5ZsqEsVa/ts34sFxQ9vFT9euX5XcZAmCMsPwRQD79k2azRDk
neBkfy+N4x67/7/h4uX/7UWiTZWUxikU4mJNclQ0yPKXFKvWO9VN8Jme1/qTI1GV
mV5Hw0ymV67RRMTUmKU20CViaJaZE3OEJT7ssNHuOhXJpVTV2nufk7hcl4Lk0EuS
g6jdJ9+v3/yuxOySOgWHxhYm1dkSOSQc3f1koIAi0Bmfm1hqlKbd4rbpEknyTSVP
b+fvjw2wkMyidlrCpz/CsLgECQCX4cBNsmG5wZ4U+0cv1SIEbRHSEXh9XzkIKXrp
RW3QbsPZTSKuN7xPgyuNVkOOVDXxLZnPhffy+IVq5i8QifxanUTyzJ//29gp609J
qytmZay1REDJ04PdXe+wUeSzW6AXkZIxghowBIBMdBiENK/wJBghobarPj5wvGgZ
zqOrEnrV/qWnDw9yRr0yxH0jGeDv+UWW2Hx2VUn4gJo2hWV3szxM6GR0ZlqBLFfv
552Pk9agV3P1CnwfedCfzpcg0+Krk5loao2yZNjhn27y93L7P18TzgnOU6geyHaZ
uWIWW5zNyNcfvnEnAHx9zdj15fdMp1oePKm80uMv5Gt4yr7xXhVHVRCyMenGTRfe
d6VWCmqZbqjQGopwE7S2O7oVSHRjuCFiCj/dGCS0rYGuT9P8uKDkfzvGxsfSWtc/
tSSBMl9/VJBSFnQlMxjQJU1AVUg9PFMJqZ3xfapr6DtIVCfywGGzQMEqclNfg9ri
5vh3US/23NA6Ao6lvjM99TGtOdLK2QGQ2ZsXPBArGSjrmwtUuGcACKyULHqgHvyK
SAJKiYBX4DktDJesW5lLJvdW7R3Hw53d18oWSuET32zZ0bXzuqCuT4VVc4wajVzc
HYNSYrUdLapYgaISp/1u9wEn4kAyoRVx2lOI1O7tcnHKJEFiYWLaBovC8JPeBFkf
qBjc+ZNT0Un7RcYcQ4cD8I5iTJFEiGnYztbqeNCrnJ1KiZ9Uu8+YQrBLCbSzK5HI
vFnjU7/OQuw5zZGLiHu7O3oBYxaW/GFK9bhe+CxAyQGL2Mt0Z950UaN+Pdu2xI77
VJiPlUbrHBxBe4AwFJ8v1i0QkvWsVtDtRy7XyKZC5pN/UDhq3O9b7SDp+FHBq9kS
4ZTRSW8t7PtGDEQiy4xnWBjVLLUo+KYX5b/K2nvOgps8bEvFiABM8ulI6jhegiUW
hHH5+cXgv/GHL4FvEm+3Hx0ll3RP690X3BphrwjEIjYBZX2D/+XRdFK9E5JfFq27
6CFQ7Cwm+2MpaTSmJBp3uhrJYDbfN1Sf8aEL5mEw0np88j7RD1Jws/KFvgZ55Oco
PRr1k4YiU4Q19Xf0YA2OhaCa98C9vhqHHYLb91XH4f4qffa1v/tBCUA34sPkF8IM
IhxV02HdkcSGivLm4CwMHpqfXcNUgJob5PGmiJ2QhzuKcCcVu9LZi4djkOShsRsp
ppsGP8nd3EiUIXdkG8cuBo1AIjRUojGASil77kOcM3EgYzUFpF64pZqaze18c0+m
yO+h0gYNm+npzlKOdEAc5F4hwWjOVdKIX7nrd3b4w9zeDIuX9aAn5sNAniwNpUd1
UcaejynAawc8No8qjybwcfFKs1vOyCZpowCB9o5WYNu+abYiGqtpT/KycZS678X3
z4jnQMv6BsuEXKQ8Tq35NfTbtoUuRsqmQovJFnU5wMARwgPoLsvdxri1vT9Blu/D
bSA431M27YhK3Hyk2M9ulePTmVdy2ImR3HF1DlI4t8ZJyYBt4UtvRvGJn6ho0rXT
nJQaGI+psgVzKRYgNOypanB8tCCDh0zcfUBEZS2lYrMAjbR4tkwyExjIBxMgJOBq
CHrTfV0/WnvNRKarX5ABBprsraAbLSJhWQM9httffgzen8P6MydZN2ejh8AYydNh
Yb9tNfhQTYPE91Fvn704wtOFnqP95a0RSoAI7O1YDI9Xvczq+5J+kn2G4Vkm7Oht
/W+uBgiYui6GmSBt2OaMyJK/U1hYq2tx9mQpOfqOwz3zVjMFtm9j/bgHSqzeb2bb
50g7FesKxzry5Vn/9g/5VSdYKsyhcD5/7VrKpp7I1CrKmfaJipikF+rWLpJNpP1T
f2FLS6QXp12tPy3SSGFhLw/icw6u5EHS965ZVoCwJw84AaJuoaCjVIaTTILz5vJq
jCk20Qfy59d5FOIYAmE8lh2C/kj/H+jqpjtznlG0/TRtNsjOpz8ODwCGcmCTJMep
BXTB1nvsxdsJiRm/cUTBK9wVU+SPeceXXhTZWRVNEvyeXeZCTUV6CU6vQp60e7Mj
3768t31hQQeqts2CH+aoalVplWJTneSMAms83hmDMe7czzq097aPgPDLXY7k4VKo
nTSBNyGO9lspbroerElsQNxIRA+fOyp/bfg1pT8kSxnXhE45PQbsjtTfBHkxcMM/
XzNo+pU/ka2DQggO6YM9CtkNr61cZ+JAzDVnsOu3bTvlEH5VegDP0J001HVY/0tn
u3yPFvv78a2+wa9DDahmsIyRfZP8Px8HX9NVzmBkIJLA3sDjXGpI233VGIwZltfy
mMYUw1shDHmFrL5m290y5VmNcomK32v3xYyX74OpXYhipx5s2gSMDFA6rUFlcJYM
yyGnMTWVH4jdq9jQcB8XXBOpaPShcraEu64lwD7qEB+5EN2K50pToVdg/AbGMZmj
ahJdBEJ/2FxVdi1lkVmIDLKdCyqkIF8wjTyc4Jp7+QlLZfq/22s8bBWjJ8aicsz1
4h6AcGMz6HR0PEsXjX9jWCehqZbJlLNSGn9zHMTs2BYwjn1TUS9xCnbipZCVde5i
p99RdWjMUVa6z0pYfmUEjb6X4mu5UQbDnKQQGvE+VROLaNOcgrzO/ifZhvwatEkd
yK9ZeONKGBX9zCTnI56mol+kkXDkFFzrtIH04x1wlTSwVny8fERN1U838dksnwkM
36DixqNqzuZp85vWaUsDvLDjl6TKC/uy04y3o6vf9FYR55iozwDFU2iC65JdtYGu
2LAddA/Nvpxd6pI5rprEw+asZ8XZ3Z1HbTTwL2A8NuMLXiT/CxD9Vtd9wP3/WLfe
wDE/n+JDR26+7Rw1euTEu1or6otvUrTU92Uxcmxbo/giFWm+vvnkglmGzgAVfcln
WxGIaw1mlB1+Hwi/VIU3+2fE6uNwzyN9oIRDYKxx2R2wTLhUX3BLyzwwwuJLblwf
+jY3tVA/AAhsKaDLBv8kjtnm2q4IfmYDnlqhYJQnU0j70dhD8BwYqK5+eQtqavRx
RqbnwCPF1kKqG+SryD1dOUr23NyceeuYJ5WA00pjepeTgRxfP92lLegytm8LG/1+
KOS6Qv4niOlGTD1jEdPSpGAnaiHQfGf1ASiiJgnx2wlSbBgBt9wGq78f4ex2gAOo
e2Vf6C2uxrR24KaZzY3G+qmePkVqFDjpqBvifWpVSD5AySqij6kHklFftUIgJw3B
XZhhWFQPtnin3B2pyWtM1KeTg+eFY64BtqL7Xs/P49C9HO0KhmOhYoYCOKyJRyn4
gYcpGG1oLjZjFKF2M8TjCbXutloYIJOM9zU4sRnv0EynPdzZYpNCCUA7wx0NG9sF
BY5OdiUwLOLar37/TZ5l18UW9Htq1GSlXhbmm+JDv5ZE0o9x4rVvr7sIp1x2mF9l
fZDB/K2lm0RCqbj11MD9MMj4nKb2RJSizX/ySwWOK+8zijEkO8FGl6Pesmtepl/Z
zXai3+2hBQjGJBzXlcsC5xzxhkSvBBwM+UM0e3D1fwPyGvIjiu6IwyzPnhoZAP0q
deBpiOTGUARzKEV5b80OkCLAZqcFu9Zteh3cVv39TnKOEg0QJmDRt5tFL5cVN9r6
cv8RGptYiaI8MwuJBvUXj40+0QZarizeDckX/FGTQN+F43pFXsQtILDGpbONqKJn
z/HeWzSwYN/8x8dgibB6ou2Bke2HSs36F4P7wZxWMAO2mt5nFPoNTRGg/yTiPGI0
tZ+49BdaJT7J12crWFzHxam6ce9A11/WBMF2/6ouzlU=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqqjUPKdVSxdSXDPTlF7QDy6hFM+tHSiOzO5eXXcprF4dO0RuNHQDAQpa8tpmaVm
W+lNQmergqUthTcmnqCW41W2TxgXQ3p2sliBvqr1INnMkWw2Ptb7c625KaGRk/5/
RSM2/cuuEKI9afCbVlqLMWaUy0cSJ47dPIy2CHov9dTw3PqnALx6S/CCJpQcmwRu
yWYKMNMQSEUP+l2bHaPpXyodSZty3z/8Vdl0EkEvtaV49kfApv6SUdajODmkd8r6
u/aOIRPeVWwdsO+lqdLHZks2sZmmYc55i5SHBwJi5BYrYU4wh4b7LDhITY2O6l2+
h313UBrxtqHXNVlO1RboW+kbFj1r9DZgGf8tjtbrAAmYbEDc8FCHEpMPfXH186dU
gKgjYSVJvWVB6D+NWrutBS23S1Sm/j0JeleQ+LJZKHUCRHLYr3TZBJSHjD4WwkDc
sn/E9KksibVW3sWljjEnazf6YQjAnN56EsUnYFJsoKXwnCUZ+WLEg+uJay8+XIHI
OgXAQUBQ/oqOet959tTJMKZGPMjDg0l/GpVneLYTGslzsZdoSHjQ6Lp4TvhZ7/kT
/3SRgGMpjR2JDhU+hghMAKTKeJY4IW+NcqavxCbk+xBTqulxCy/GuNQrul2ykp6i
+1dWmve7+dESbA+wrxxsU5b+DTdaFNUNCcN/QUYEzwCwTCFWAlJ/6LiSLHHMSkKq
+LMWlKCkDNFZjrsKBBOs3wXoKjmQIUVy0nAfe4NrrSsbvCZ3QtV8OdTFPwcJU3yn
LkfNBr1AN8L69cFQEPGc7ihipUA23qrspB6AZ5gJhcwixm/n3kbBN8bzRDuxGay/
FKukcoNfMcN0BiiKYy8HiaeddYuX010SoQtxjir68sZEQPNFdNAHjvTt32TAT9YL
ETDK+u6GrqoXjgbYUpsxSgXRw1WEwZXwUUkcYI9GxzehI9MEK9Y3ggyiYezY1LTb
+oTv71HG6f6nChm3A9Wlhkf8h7asr6LwoXdIY14qoN0X0V9V5sG3eHn75Dxz1KBt
SPbZfNfOt5A7xAZ1FqE6wfbC22ng0REdUZz/Vw8rliGiSqK/S3kHC7qL95pv7/d8
SwbjLlPqfBAWXZm9rpTz4wL1r2VQ1xK6emRRaz7OAj+ofwlfNVWpmjkmBxZGKG66
IuPJHiqwFpsZujK1/p1vVVv65PnsrzeeucoWlEIdNmVjRSstMNOoF2kAlDC82Cqn
m/2MdAxfHoMw6PkVIv0koUkrEQDUMMTGzYTtcOCXWkBbfUPhbD8ycyhXNR0WlOFC
iARxa+Unb3XHHiQSRBZxuXaMhccaOIzpWkuKaHBiaaXuHYTR2c69OQG66tRRBnqW
lrzMlPXuCP6uh+rstjnDBmVwViemJ14pV8hPE0uoOqt0Nfix/YA2yhu5ns1Ezz3z
w63w7up+zGQ3x3b9GM7kIC0+pUHXkKkn2giM3JrhY7FVlsQHDNB4atkCNPPcuYVK
tdV3t6A6eyKhcbv91BDfX9JWHizsU8mPCWzGd0NhOvOntezYaOgIxVYU8RyBGxhC
3pdELOyS6eryDKp5NS9yyNh26pVxhIv55Z9L2IwqoMK87LuTRdwYkd6R/xghpgWn
9FIGfY1z89JZG/RMz42jSeU3X5flrRIUrHq43wRJ5yZ4pj+4uWfW3v+vV5yLwLOU
Ulz6TzYBW2x0FPRUDZB//iZ37tP2b6zdjw6fBbxF7P6wb10IAAPBemEDvrvbqxuM
`protect END_PROTECTED

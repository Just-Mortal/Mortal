`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3DgHLI7YbA7s6uV2nqLsS17JevUXE7X0G5ZBi1lvbSCXJIn3KgdfYxFVx+CHipp
t1FM++H/3oE9E25T6lgcpDNODqdzevxEUSCj3vOet0KqqGx6YR2XRGEGkxfKlbyv
mKip9zbAyMoS0u4kXACpH1Cpcoh5rOH2S7VThKPMAiaw7MHwL/Q9s5zbTjPI+VZv
kTqLkwxpJ3g0drYjQeU/TfMlqLF18s37OZRUBKYlaVG+np/tLHob/DgV8be1/b1R
w4vX4hKii4XZDT3yIWEfNlv/3eT/0sP7ARN8auU9TN91jYMSY6qIo7oAA5e9VOnX
9TngZHnVQgqbDFfkuOTPmG24K3NIJhFeLVrUP6wnt3S40Dsz3HhxLjR6fHEAWJtD
OVgsYGqyzl8cOZDTjd7lFlzg92fU36UWoHDTrnwn56NZPt8gkOfntKLXmQfVWaS4
TFyiszDKLLL9fKUmUPBqzW5Xwxz2z3YK+wgDNKpS7lGS3UeEA6IGhbSkHCEqafS1
9bkKjtW+vGZM/1fzmAPonqurQimDPLfOagq+JdTQRJQRFYS3biqtVUfG+1zvFnr7
WW66NinW4fcTxfJ0upH/1RocP2vCGILimD24JWsjIYhWeuwLz1TgTKH/IKAl5j2E
XjKvAGn+yhiWoiZhgZZ76ZxtAG/LlpmAcuJXEZfmo+t/unuMX/GHiTJ7VhmpqYh+
S1U7kyGmZPlwp4tmhwpd6bWGxUiGks8HfU7ftcEYqPT4oGuE3oda8QMOe1XeS6j+
KbDkY4SswqdFNEKSzkjuExVe04rls58F33oZwP4l5+hLJc977ITkdIBkNoHD25wa
KZnkF8inzcvZgu1e02ADbsKw8W4kl6HyJiBdoA86f8qV1JgF1reGAKlnWBXubPFM
Yfr4M020KJ8bdYkphTTRu49s9gTyjgKqHvmqrpJlwQOB99ThUa5w1gluF4d+XicQ
Jy3k6fMnbl8ZcejuErS6zygdxg3ZgYpdoCPMswKNNWEf6wsg1JiGY7KQ3xurc0IZ
72w3tAX4trBHnon9ceW3pRwnkTunOMuOqerb2bNpVFEjK8rQWddaInasA5c2ebhz
9vaUUvzEXI3XNVdqbK91MakJwrBL3eSKfVRQ4mkBeef0tXZiBMdGwB7PE4KFsKG/
459C78T3NMhzx8Wr+RnsI3L599R5HAxuWdytzplHXduB47bnT6R+/TJKJrXNmYdK
v1FZma5CZ7CEVFjpls06BGGGE94hEUhRd9BcR4/E3C5VlMjdcnVTxWzY7SLGSfXN
ClsAKCKnSgXRts7Z5nOuZICDLCmcrJzHWYU8PAmzEd2cyh1adRWWP4sVNyBOZfx2
B9Nle81lMfSxzlYbtWLKzaxvUzJzDcy3uq1LYHiM8N/MJ+vxY18wXOJMSJfDERzh
A6YkThBLMOYzbQPRQhwp+tXGKRbn6LSYWyGn3Jk4jv4/l1n3awQJT106L89A3BZ0
0OF/O/xvK2kh25XGQJi8XBFoPXA2m1UP1Ofy9OyMfuZ8wmRNz2J6gwYQfeaP1Zkg
Mw13dSyVrEUzB3FqgevVIfAmPH0GMnnbDLBCicZIXcVr8GgZgPQuPkQu0g/Emg2g
0dKn2vsCc1Cgy4BTNxGnYSpyErqOIGQdTNLvIpbLDiucy7Y8H3A5UdcnJs83to8f
bvJToGI3517o89CcAAzcuA1sjOnmHdDrWqvt3OZ3O4E7JBrQfP61Sl2xbdLg4fei
YHWcDvEBZtZSAUOSMkex4a980D8bl+NQZESvTqT9OZsozn8BwDsXFAKe2JEL+1eg
5i0cXYWrDYBN+dSmeUtBd/W5wuC7qOM8Ub/9OevC4quOtFIe6O5MIphfg2CI2xNk
58YNCIQ1zc7Eip9nunQ0NBAsTGyBrwirmpS0FMCDOlH0ZrEqWJz1gQo48Fi9BAnx
wHRJT1wplgcBdwOsMweB8mUsih+wEUal+ADkRPkZuiBcOdMcTiWAvc3KwXcBDZQS
qFD+6ZANNRTHvgt/5B8zq/cNCpyL3vF5lRcOE3o7q9daI02jdb3jX8t9HgXLregC
2Ak3pH+LfM0KuabKD8YsFXWKzyL3SJAAwO79cbKlna4BFTo8OyL+TdIux+2duU9h
xR/P1MhKpHW0CJqaYBBYYnKHWJvt+1CZ+O5z4fmlpVuv10v3PkOWJNng35QPZXDv
8M+mC7KO+SGNE1EkRlP+jgEyJ5jHblZe7rsZwEexAM8vT3de6lohyViZi2ZRH+Sk
23ua5/avsPDENiKi9MYDpGf60iwPzpr5PLtL9PB9A1W+qJB+WlVYlGvpzjMZYyDw
D+U6SpO1Ur1NwZHavMHQr7DDVE7U6A+UE2O7aJiXYizH+9CucpqwitIR+2PAhY5K
3d4COV/Icd2n7I2685vOPhL1o1agcLdsvU15XnMzvZ0T/o9KUjx6Tz3CnKbWbbjb
srJ64qjtdaPrufJm9yXzO5Wk8lou3GQqdjo3XAHedyeKIVc4vYvzsIZR0N3F4xHp
8t+/0hOlF4Tv7uWS5ebm3lvVsE1ToiPJKK9Rkao3B/OSq8UXJsFZOkObLLe///em
VEdgiWhNRSloch10UpF8MDfJkeDsgjI9HJRPc+rxaW1hrikyXL074xO52mDJLT5l
Akr/GHaXzpgguf582eUyDQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
56r02VlTRJbpIpDt7Zsa2m4NHedHFIftBM0ZPFZU59TvN5N8GXPPHwlCGkzgB0lu
t/qTe3yQ6FSehC2tNx3C8l07K4xl3ysgv6By2ha3Q8jEeY5S8TN663TQ9EJVpdhS
xEP8xF0RHaJ5LpuW3vD6b34xDcjYRQi+WwDgibXb9MFKqNkjAqCh9QwbPS/Qp7EU
vEYGWea0GL65fgxQd+1V8HMulLSHqcpSH0wxOdx0bbsSGt7B+B/h5SHhwZi7zaVr
FdRmDT8Z1rcKte6h0v3d5eZ+6AC/qsCFKglT7U5Bpydx5CD3/GFX3fuPT+dlFGdv
rbEPftD0D0NvD1lXqN1EfXNDh7WaG1wsH0BqgGZ3nG0q96JzbT8R4o3/Y+G6baK/
v2i9FCu34XE642IkTENoLuC6RKWkMOJz69Rgav9V/dvX5OUhE/5q1lEto5frfvrh
XnYverGyZ9yR/UHdCVgFjVZOZxjGqwK9a7n4uKY60HCk82hA+BH2qzcDz1PDx3bD
mlvFPBBcTwGMVj2SRHr/XsebmbL4K7Er+kJK8x9yhO1Q04NJ88sgpT1fj55P1u3x
d1SrjHh7qFGSDZjPLzJFzLRLNh5hvlQjuCXgCrrhZqAg4+hpHvN0361axWw+fSbU
Tnn7jPVKbk5mbnIOPTfN88uJIcSJc0F1XTMHVnf5J0U7P/nHxUI/RUVRsm3gYeWa
me3uwEXXPekC8jqiyE/tDFonMKHHiY746pBh8S9nS8md/UDX7gWjxJvq6btip+PL
eoxIJIpqJCje9XtC+QfQTO/EfB7dDp1kCRuGw5Cb2sCRoFHS4liElzbaVkTAOWU6
3LTldFC/vmhec7oDLwdy5nandqMr8iILouSgH7gMDdO50FCmJ6pCUer88RO26XrW
mfFW4CWxJD3kZhZ4MfWUL1jIj10py+P4y5kFn9i+lP0avH0CR7j3g8V2ax3uC5TA
5w6dluanFAQHkxIRx26I2nVA7m228jrGeRY3odGWIg/1Ek/x7IUo38X+n10Xrc7G
3hFW8+PCYZmEhYUNYgldtqvjnhY9wHxS7fQ2EFIyKymUAjzOvwVReEz2oN4Vi7H/
zhl6xLwKuWAn3rE+Qbq3DIyLCWAzm3J+qiEWecMdCUXsZrZTNP7oQpbp5N/vd3OY
eeC1SRPmckePQ38kB79VBOMgM7nXf5oaj8sAxY2bEm7nsTY+MpgtXAjbxpFlZJiB
oGCLXZuuDUepvSHK0+e29buIr1h8YBHsvPGVnxbvXmINYtYfwp5WDmOyykD5GIi4
UUgR5YEMRqGmnOQuk+QCIcK4Bvj6eQSHK1b0mJRJ9CF8CqwDJovQB5vJ9J1fqUml
Ye3JSNsuNkxlMk7SBXBe0QEF/baWDfl4rKBBeEwS5ee85ibXESqqQcM7iHQccwhR
ef6rvP5aTSudthfm3Shw5AW9CJYkpcaO+G2YqmI/47yoT6L8B677OcvWNZm0Fj2b
wRppg9asI9UwidsV5sxouXdzUtymsm4HZvvatCVjzDkKnGh0DvK37328Gdh+ksHc
vrRDO/dxQs1R576+q0SEHBxrt2HwNRnV3t/SiLQpHxe3yPZHjtPCIZpNio2Db98/
E+SXd52kDR1eux2O9Z7BVvIMmJD2GsZg/hqi2OqrZq/0/n1V52BC3gXHocvrSVzE
zb4YTxXHvW+LKRRBBKNzieus1A4ROUaaQ4LLBTZ6NDeIKv9y7AXVnfzYxEdJK+tC
zPD/O0gzR0DazYSyrOHsI1RmYQH1sHyiT4oLUVF4PbuRQQB07hRqJrrX+SEDFRw6
FEeuK6K55X02557snrqx1OPO4ircgDF80jlP3Xy7nIUaS5xQByWARQBgUcLqVjvq
yBypE6UyAs4HYoVrJfn0EdpRYl1k7b0UEKudQ6pXTGaTL5Xk+Gp38wNy01XsTidp
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oxy+LYBajV4Ys47lVEkJoGJBpj9hshN8QYtAmLfJNXlZVxvGxOfVzG9yYcCgMKaS
Gvp7ZeAoz+W3qO8ZlzBOGFx1zfz1h3nqhmYgfQVPT7pNYILj3OwnJi0MMFPK5I+H
2f8zRSC5Mt/OnvVVbuqHh4bEA2azZMDU1i/sJY8QXPsaD1U2r/db9OcHr2tiQgf7
6hqpjbrq8jHnqgIAk8KWhmFqaXeFHsMsKjl3mU0uhUAcV5gc3OF/b0u6d7MQb6yl
01E+qnQJ7w4uH5M2pEIJMuJ9VKlsaDtCSNpPHYQPlXkl/+Fj7XiiFEJ2IwyB9h0M
OuHz1mJgYIWGvC6Ic1/bDPftnqx3t0sMbasKyuIa+VuJ5uFJmnzr1rxA4BCgFoVc
NE5Eh/uuOtCgLY0HeFNcR7+tm9vObT0RiQpnvW6MmGUudLSScnXxaKWtGCe8KZ3h
oTnmyWnY6fvGT87xMYlYpv/u7PqCeBUjrzO18zb+GoPi79zEAxoMJKuULFJNox+P
4aBLfjSdSjwvMlHHtKrl3ApyaqVUGRDbYkUlxYy09ENE0dku4M5efqH7VYLdz2y7
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
awycjnhVGvh66CEJwHeYhwji3JpwWYqkWlhICsgg6K0iozaFzq8I9HoHwB5lcdqB
hR31EqLIxHWB2XtzGQ3zo3sH3ZgT4Xo0rv5dLSwMGzMOcNrrJt9zo04H8dVeDCX0
CCVnM96J+uYpOrAft8BUhofcTPZR4ezeeLTCK2cKpPo20pP6ox8VhbCaq/uLP1Jp
iMUIZxklv/RcSxaQRaXW4x/PDf05l4ejCXE+uzHrTb76vergtR4joTyGt0V2Fg72
G70E6CQKGmWkR1vfyHSre70vaKdjAbhgGZKXhhh3Bvsy3pLvQj1DsXaexS4AkEH6
HJ5s+mKmgC/1YLRzKkrO7IeGZk3gEVAdKz64Cpfln/le9R7MjsxSqKEmYoaKvT9r
kbD2jUMKTYdl2jRLfhLZDYxnwyE48BSsPGH7l780vhzCVaA9RYLX90nAxcqip9QR
CDHUoqt/y3jQ9R0Y+z44L1+Fl9PTZRg4GIKKx9WXVAtjN8t6Ce0r8gDMjgmr1E9c
gzef9wRmQyiYb7FSdqoY3mCRsfqINUwl07JXwkswjBR5ZMlVBzQXzwsyxAQ6wHfW
eVEPo4a9YFpIZXTzYQ43tB4og5WEFrxB+idZi7Ec4O2tOhg+JDQYRs59pQSvMScL
aIyFzncGKYx1uzL2RUGf3xdzznuQVs/vzSa2IS3Qn1wSxrRO32b7fTJqJy70fcaw
ZBeG1/I12+rOX6I3BNq7U6jvL97wZSrIX5fOskxvZbN8nR/VXOsWG6wh/TeJznKC
5UsQy0Sh0Sv57K4KJXRwKUF7v40ntG/HRb3OekifpEDGFr2JsWfXGC0RCUGGUCb/
ZIM86K1iwxglQRO9Y96bQY5Nv0a1R22oudJk8gXYY0Z0o7w13ubry/0i6/lZ99+A
fWInBBUs02rSt3W9tBByDRXWK9na6Tb3w1W7FC0Zfai1i7NfpniFJTWc7jtLwXP6
0eMs0sTKRY/r+IX0h/d9OEqsVnj1nvwLp+HGuCTbLLGsMjDt0N9vkBfsPONX0mjK
jBy1Qg+d1FQXhQmGMZEXfSR3Hw+3DedwS7uDAcWm8CkR4TAcKd9HY8QTVQd4/b2f
OknHJaogZLA0+XsXBCSBLJX91YxA86ZnhpMXAFzuQjII/U5qoN7pL7aBRZDDpc8Y
Kaqc8mNYEDcBEME6OdZm8ktEKlQf5EqJjC44SF4cx8/T2CFl6XpApu7+hk7tQK2L
4Qnmd+w++IlEAwvnJjmjC4aLk6yBETaG67bxQ5PeNE/km+qv0NFame2114NjQr8C
JsvXTC4MQtR9poD5exIsKXW0gUjjf8PC6Vpx9P/oT4xfoDZ69db/3v3XwGVF5rgd
apC4nriDCQlMT/5pOxVtgcE0DZ4bIJc3OrBMk1fO4uqavHcl6wsltCEYdLO8SpUh
dIsFHPxv572q3KwjJgb7f7U9hkcGFmZZNB58USYGcHZBL5kwtkRthI6x5UKUvB+A
LUITWsK4UGG/bcKNYQm0C4lSUnHThyI3Hd5SXMv/PvgtJ7oemOAEcLKTTvqS3u8Q
zpSvRGr1YsyyEnpQJd0IARG4PxYDJN/pSbnrx5eb84a7Q3AAvzdvFZ0S1HeweDm+
0frtLwK8/6l1JSXUorF4nFwWZlm9gfeUsTXUxfzSc9PC26OBPBIH9QlS2wrdp7kN
0tLeLA9r+105ugc41BwGdfw/s4SHz920DL8kAixgA5CWOiQigZ8g9NYEnfaPYp/3
sHRK0XWtVIP8CLkUhFUGe67yPXgbGQApU+kJtoIz2eP7CtwnXZ+PLKmvxngbUtZG
Fj1/H46q0h3RSe0Lmwn/RQs4OZNq0iaRRNiEEMl+ek0HqdAkrFpDslayXHNNf5Rx
/pdGCCSIyzhx6VylPjUrWNhFj7O5SZxJKSNqqwFmXPyDnCCE+1KuaKrWB6zKONEJ
OIL2Nbbnj6BThPPn0Kyl+M3cRhYdiS8UlNI9nK5npvcWEmgFhrpYggurhsS7r+EX
qXE4/F9VzPc2CVgS3Clt06SrUXdjYXclYw0S5ZSqSAknouOIvaYgxQTAC1nRrnPN
SJYrPeggT74Ist3/c/9f78HekVBR6HB59bNYjJ45ofVGRvBi1U9aK82uSHvEMdnx
WwzjkEj1kLyxC7Sh0q2Kw6vD1CP1YelPcJ9HraKa+3Vq3+K9eF4v/knNc2LYp0y/
25VYY/byLeNSleiHi+obrWmlQ6L1WY/d93m9Z3kmuGUpiJF3upQ7BHwyI71NatvZ
bdI5dAUKnetH2eDMqvR0OT1xIA3PoFIOEXWUMb2hmws97PO+uHha0IKg+ZeU0eYo
iUBRq7BWnhVM7pPbdTlw5lZAT0YY5FHyiIFbHBkh7CmURi59CN0DfVBCgbz1+Kv7
gsuwU1lSe+q2F5Mh4zYTSkE5A9Ace7/dT0nK/I0BCYykGnyv1hHUi7fICfMcmiJu
gGV1czekr77ajgdaRxFFpuuFJBC1hyicV6UCRGXGPaLkhQyafh/ByuaZPkSATbr4
fmu7ohrcuVy+u3ro459bsywT6nOoms4lAoFNYrv4CjCVbymQRK5bYgFMGXcfEzaE
U7FbzL9ZSe5+LBSK0UXV5+e+tIp+Efwx2zCY2WYiqsHykUFfK/XxLqWkoIdoxNvC
Umq+hGjVNj2VUxEu/ndvBCKRhhxmTxNkGkZm7OD6MDe7Wa0+q6QfevZsoaJcAN5/
R8T10sYDXtYfeYGwYjSmemCd5dvF0f3kVCXZoVkoAXx2GrPhf05POqnBRjIu8xn3
D17ldGpdrkyg6VZIC9t5PuwBOLv3S192HBFdnjx6zEW7y6sedNunlUDvKVrotzKb
BbXB8GGSAakpd9SZO54/ELpE46NgdqO4i74ylAncj1IIOoHqU6oxcp9aEWt/+7sf
DsC6zcd+u7/KnrXJ6N1y5trJMMQ6dr48XHDeO860srh2dKSF12L5VSkPk7hiACRG
B0XY6Bfs+g37NMVL696Y5G0xqvmY/3GytHe6n9gxyDZpnrLDSioxXQWYWQ3U+Y5S
gYw52FwTdU/zcjBg7wqztZ+swtHa7hgYJB/W1UAAjnSDmVQ/MctHj0kzpyGp0wEH
rg0oXy2iyU7vIkuAQwzsyo1dwpLSk/PEkXI/+OF3qTPH5KnrpUZqlVZWEbaMuyn8
GogRZEmep1Gu+ZVtYcM686l/dLIzhdnTecc0AVqzLsf6Wi0P3j3J2fRF3BYmEB8M
Ylt/lDg7UBHWB0OOlHKiwcw8lrTc+GTIC6tsKKbz16uPmWIEHuw2pKCAOSo4MPb1
VBOB/UONrhEoR44guzUycJvAM2LYYUB6vJuWXrtdFB1PGhyzFkyEDbfCqU2xT3Ci
vxVBJVrO5sJ74AVLBPG6HIQgLkmg4/s6MlYddDUfTXQ2KUzFzKVZDe0VlJF1+Twj
U9+ff6OgjVYKFamgumyb+UdhmQIry3w/jb9LsrjaqhyAPyV281GM+4JUUGIfFZRh
HVloKcAMk396x/3x1Y0AdCVdDNCpr/MSM9amFlzRTODhHpyKvShqAyeZqoU6/8nQ
SWBo8mVMmuYtF5va2g3hP06tjAz8N0ENleWKKMbJZM66vG5arP7UB2FYB3gNK7b3
ouXYpt8qZz3Gscc7dNa5jqtbgsl/jQyNAqiGh1V+AlY6b47bwpE/RzdwDO+o5TfP
ACu7bHEqllxXZ8wLiwYHpYh3OrZoPf7nPFEa8/mullTpdaob/5Pyvb4laSj1bHFZ
FBMp7/KMINqsOcOaHGQ7ppvPrcguhtCoYZ/ykoUGWrfz8W6b3o4UkkDW7b3HSSho
Zs2RJiyTnWDFbc3iH4VChuzquQDxHZL5MEdWaa6JW2e50GqvEyGQXijWbG9ORfIx
5V/feZvN1CvqUdfXLDEoL3sk1fI9t7gYOUZmd0cWtffE34bq0zuhiNvqcGWGguEj
1mWjXB4YOzC12UNVb4VjctFpmvCv3dp5GfdrN/SMfQA+sekvXCsfsLOaOsdyTxlG
tttbOVEAtPfkiFs/tfYBvYne3GhPr5LOHI6doMMkbS2GpsrQxOQP1O92fhC8mGYE
dPaDZZ+JpCJqzAE8sKSfduhyW3te9gfzVEW71L4TZwIaoswd/xzXBGLQhe8/Wdwg
ddeKNvgWBo/hY7vo4UUzqkkWX/YBiFDVVCPGcja6zgObgE2MAjJuzf/OZ3ACuhZI
mdwh0zJN37gUavXPUe1Zoq1b7h6TfHbApSnGwmDEQyQRa+6u2F4vyzWTkRHhpTQv
CvHA87GbWr5r/sYoafQNovXIm19q0h73+ZSJVbpBffz56UAlYontOOlni/YVBRn6
YLIhlDUhWp1a5kZ3pIF+Kzk06wSWzxcPC3DLNmUhdaPYZYcnEfgaUZwU1CqkcP4L
0vEaPfMQ1MTzpDmEVi0NWoePe2PFGqcLN+rltb3bMzq63kZ0K11B8bv6nK6WKqI/
YAl/SGdX2jk8QM2W7rTY27i7X0kAaauvoxZ3Sd86u72++tQOuv5Jh5Qaq/iWbwiz
AX2cpCYa8E7GLdxU2GLvX4ss8y6/BVr/tTpoLKuXx3OBtRPo/zQAUHK3vtAjI52k
ZBdDwIY5RNkI5wb6y/z0QB4/8F8486r0E7JqZ29goi6BUsvpTt7+BmfvQLBDQbmB
9RpY4esmqORW7hWwJ4YLuNgc5jJ1QhYqnaMonDXOgcCaxtzMaWcgWa4vTAN/EMte
KX9peuRVLdat6UzDeXzHk3MdLQk/tqzX/wZwNhdC3/O6G2WlHI0CG07GrEqM3loE
iAtbXEZah0nz5s1Al3iGLahADH2sP7qS+uyBAUrtIyn0hdLGk8TcxvFHNuiHw+Fe
3ze6ST5IrqjLKCeIoWhaSI55ITQlLj0LQRDIoQ+eZko7XOrRMOO2O0RRhhSBCzHY
AM8hdFWBVuD8uJ0TgNrz8EqUqPrLaQdujcZHz0EazVbmfdINDuPqpMWr5gme3968
DIADouYpAHhauboNnFJbpf3ZR8cTWMMXLyyVOjAEt8N9FtE+mf/FaJipeg5ig4Dt
sB5lWAc27jN/qZmZkQC0N7p2Nd3Kfsi3fwFesvhAbRTaWd/GvvNINUsiHkN6RusF
XUhlue9bIR+yvYibGc3/KNjTvIurdxK4/OAIL1EgHAQLZuBaoXixhx78oG8oXs1y
T/FApNW3E8w6p3P/Rv6Xqt2LCw6NYubJFbqolhxr7ZINqeqWwBxRfuAoxPQWPMMk
mD29aDA0IUVz47b0h0StaRkZTAtVz1P8SX0N+a71xKEoGypXnocxMoHt71rempQ9
vEnUfIjULddOP0VDgW7d4DTvVCqGzt24bIC++ySQdaIep9951RlpYID6zBjICnWA
L+GYVDEuZk/ig2VuHXDQ9x6Z7sug52912mJBlTsRZcThrwNyeCaMy8rvwPxECGw+
MUQTXnMpOE666Mo6EWyPdBpFQe1+lMAeLcGe4WrDm69Mh4Y04mqmKP/DGrhfp4V5
QOYcQmjuoN7CVrPoWGUM/buCTnuumFfYea18EJ8MqopkxSM96TUbQSf4X1W8Y6Bg
QWk+aFPOttJ3RlpQL7p1qavL7tuqfkqJJQXxTXUu/vRqQs9YYeJebKluWSOd06+R
9/t4C28QpHyrqVFfcyb9f2MqUVfFFqVITaK8CENJdka7b/Wwbe6Y8JDw7X4cFSyA
3dhaTiB7UMwVE61s0d1BJzmqR6LNjo5AtGEqyWceJqE0gOZGGr06aGvCseAxcgjp
Yv/fC3RDHixfPZV68xzoVh56LyLkH89rl7Fa/LG+u/qA1iTK0DyqWm1HJntGsMyc
pgyb1cDn5ouiYiZlmGJgi+lbLUYT1OmSPx7W/wfCmKvHmXAsF+zzS26VH/UYdHlX
tZpDBiYTJIbwhrf04bebPK/1UyGM4Lqk3WpoGmdfeAupfDnVCzQe7+vGSd7TCfWY
9CWp1pnbNldFngxynqqax+KvGQaMNjWpKkzsKPvlGO06dlD4n5FJ/IpG9qzdw3rC
gZDcSs0JcKCs5TSZUQf1uKZLmPrjc8AQWAdPOAA16u70r8030mApBMM8AY41IpcH
P6rkv+/upbZ7hC59iARsM4/2YNpqR7a3JljIaawyOtgu7/H6apPI82XJSugY22vd
7TkCaeCw8k/smZu+SgPN6LSErCPhidY39JEJ0ViDu4dPykJ8llsH1+ufefg8BG82
0Ml4wxxaCS3uGYL1pIIiqMHQo9QBXfRWR8MzKrRC8hREwojKBAJdzyU1vIOKvT4T
QOcKpKzY+5tNgCA+49ERRyl3TNriRxWSWIWXAx+FQYf7UCiXKLsumYnw/jhFJFjz
t/PEzaHvQLacyxgV29k5SaUyIsI7JUP57aulUx5c8X5MKnVkIAj7iz0dkFS5OQTK
JO3hdHWK/XSc/6EzeNV/AC0grDotIPkpXHPJn94+TZeGFGxPh0dKRr+m9zHE0rWK
yHhmUB52HOXgOOfGveQc30Y+IYBJBCjmz8sxacErqNXQiO2tJGcjsz4Jq20mXcqs
rj9Ii8/jB9IqtWcyhiVEhi4CMtR4hGyFyUGExQeUY/2ujUIC901xfxgi3vFrv9fu
31YjXnnc3mMexzoFonpA0sWXMyQ5B4mnWGm6YHkTi+VnCOZ4MOR7IkiDVgD5Idhb
uAkpZv5YajHM3uNcQEnEm1ljqgR4kZSXEHAVgVlY8ELfdak3PG1QEGGgkiFKn3xG
5Ekb6PfoTlB8evI6B7Y3wKGQ/VuN9cCa/zNSSuyotveYetqM7nRTs7rLy59nrd4X
Ak+MrPMa0gEBBkniF28NQ3QHm2+odwpbl6AAKvyZxJqiQf49XHBtR2CXc3F3SaOt
W8badi9Z2+EGMDRJKxRAZP/BQs86dCihHOTPC3Z/yxlnrN6l39jIuxT0LNflygX/
8PEfW5kStTnbgezwBSusAaQ+11eI++UmdAlCR8j/Cp6lKEs3xbzUiLzl6sTig299
fUK6czN7QcUaIQET0lNxf7AhfmsvsS3qBpfMienI0SYllfdkbTBT3wiQVuqOMzo5
eD14eH7K4VcTYNfqoLiY3YZsMPw6BP9a9muX7lQ6/jKLEJoRchC5esaLEHj4oPOs
QtxdrBreA3490Lid9a8QCVykmsCCIDrjaYkGKydq5OmFI1VrtfI23l5uL7yKVxZl
drktvkqRIH5WNQ94OiiUVLRY1QcqaKr1sK8/UM2Ci+bobazmusBEdbpiG77oqskx
OxargXe0zztGbhN9MniGmdthsfbGXKQ5sybHdHDLqpauTn7oTIOtz+CJ61raRWP7
Z0BeRz6pmkmL7cIMSKbj8DTBc/vZ5S8OkqQGdC2W0uqoNgwwDG19dMAp+wqExQff
Vy5Fz/++fnZsBrs78cZTeyJiaCSROxyEHhvoERKtAsWjPupFhPS3T9PSYZuDLQW6
7xoLQrtGAhj85CmatM+BMF/DEYsYdUz1HThAiiv6hicEKB2BFYHYLHe9MYzG667U
pZugA0x5v7bvgoDnJUpcixVoT7ZlAisl/Wi58F1CBtNSDQ94IR2id+nyAze59tDt
Qs2iDi7pE9h3A7zxcW1RWCpjWJkKKbE96Sm8Bb+hhjZnJ0pPEa98EQy1L+XzdsmJ
Gl0v/p+ZOibsz7di11/Y1pA/jDUY2Z7D0bH16JMeboOQVrfcy7MKQpvEWenlInPp
PVITU/3jGLftpwNR3+NDnWm1b463rqxGc9EWHKS6cnrJuAplYYICgBwGzMOnMUro
SluuCaFX280zPVcNDAsh2c8+Sy8DDrOruoD6l9EcEMkAHg8+/OdN3ipQ8QhKt6vn
VRw+mrXOAYcCLh1bxxnoGgdyeTtzvE08/DNiiK/DT5kur3KhrDdYpiuhwX/0UGMl
bbjL/M1NZ/UyzgFBhX932aFVQGwMmi9z7XucKQiP75WztYPkkTd6LhWZ5eSvo6Nt
wMX0Bm63q16rrh9XSrEGDNOJUxldI1C1FTZ9dF6OFYv/OCOREA54xSIgBX5S9OEM
dgPKv7aUIHAkH09Rmk+feDlEslqDn/faKgvB0y8nn0H45/WPXQ9VMzsCG70jpD8r
NtXr8R/2MN+ZBWuhQfz9yWraloo1FPejKzbFG54NpmYsABNGomw61/vlhXFdaDQV
hNADk9IFfina7CpTW6OZeXZ+3aGAwWTV6/ZI9d7aWOsl4JyMPp18T3GktXfvNXwP
kJFFPjSAGPIRYG59t2akVf5Joz+cqhwlgmRpYsyf87YjTLzyjcIUDquOGQuTIIbA
kcz7VN7glBcBoZO3nVsFfsxEgHMcKimDBucCodHJv3BWITbeN2iPlui637gOa0SS
DlpVaCaSzLcLVFm6zFS8bm1jYzCUzgcjNnung+8Kv+3i/IpN8lsHt1xc6ZLrSnq4
J1RJkQvQsnOSJP99h6/J9pZ+JN12eY6op0DVQ2iBUO7cOyWMeVVwqpUrDZyIX8cf
jdLwOWpagjdf/rlAaH8VTA1LZDHx7iDeR7K6rtlnAHaEZIP5p0nC4kbOgpHopsNn
xoSULk+qmLQBf5bNxdtMC7daiuRqi83979nQwD2Rf1OPhtZeFaUDa48ep5/HN6/h
gtuYo5JirOlPgX0WMORVDpAF7D2DUPq4GhqZQt59H2cYI8cEb+8OieEOL3U5rEpB
yOTCGNpcM89aNJS8J965+rJXUFOzMCeryOXV3Z+juPU6vPhFPYCXVJD9q67ACMdW
34/kFvJ3A2I4G4y/PF9v9fK3yMrBMBsZvDfvinGQ28zUL4SWyJLhaAIG/VprB5JL
DebVkE8TlHLPA1bMXWAWWp+FI7EfX6v3nZJhBZgjY5o0uDfXExvYUX8HtmhR0QJe
0ero/cPEfkwigcH6hYlos4VZgmqpaNJ5IRG+6f3rUQPbHSeBC0BhnB9wRAGZUn1v
pNIEgG2PUAKgtqQ55+IA887FoT2sTlKzf8kIp53J9Rx7aZXQaD/UzpIhSa2Mp/ZJ
b5f/Y9VjbAVyRIOTonzQy6pkSftVrRd73qqcuRHKddyzgiKN6uoA+Sx/+Qctq4C1
QWBDcpKdRvZzLZ186QAGM1aThHsB7IFHa0C2CRBalsq9tOLM8YZvuWlKbjws6X+j
k0lHCf4NpdPaSUCoKJOCaF2ybN4DmlryJdZRZcPPA/leE5AHuWK/hrDLTXTMPjey
PMweERHtmS/k4V75GZAPxuDWi7KyCLe3i+hoiyvL7mI5OdGgqJAM2JYMhSd77obR
nf7FC9B5owO8bvKUL8vqo5ejFtkGPab4XHRfVDURMKn5s60E9F32iZLYxJPgK892
l9HPvOE26+pff0xuseS8FPEHRMP2m1njhTsXcMIhD2CsZ9eoigCdIKSvI3jqKtQ1
3dJ31FEhopTPMA58ZMWGecHS2vkiIWEeUiTMPZ8plY+V948GTQXH4BoshoAOGWM9
APt3T3DX1vKAIPklp6xRk+dq5KsBKGaJ91EBhcAa5/akrTtEu3bckaN8FKOe8uqP
7VVQ/KwuoxAnEIp8BIOf5zYtspYrwovoh1lLTYUcbyxe9aZqA26vFsi5MUajc47/
FoanniC0pLOk7iDVE3fmzB6e9Ydq8FAgGvPplKyrz4zlV5vhuj0UhvuW2KftOeNd
PwN+YPu+/6LJu/Ros15cs63HTmg6lxycEowZXuHClLNp0MFXn9OqwufKN2+oiubt
i4PWociFUT2SEpjm4YoxO1S6XdzxkxHOK+povviouON7+kNzXRRNjMZJ9sEQahav
837qud6jr5x3PukogOTlVui4O4jqfhnnTn6cZ61c6tdlWhoy3+3Sp2i+wqH+pwtl
CzOQ9St9tZlKuEIvpbrOgzA+mgI10gvxpykfEcDi0SIS2Rcp3xgKqJM2X805etqA
KFvqCrXKdXcgXARF9kklPj63wmnseYd2M1+0aPe+QQeWUJK6Doa1FHNHTxlKbIrh
DRwjW20IQl7Sdt515guRJIw3sRkNY7qych22t8/6wSbr1UM273GUL6Q/TFa9MmCS
nan/NFVfbAzi9zzIM6N+uKPezrpEy42gkMy5C72gAO1PxMEeQQ9ViNoMpVyCKmzx
+PH8htwtxGPS+XVac2D54aTQAU/Y8SIFjeRvFyw1spOx3segoD5rf/m4a1tuc81s
7TYvKCzx7gJzBZ4dyFbXGHjhdCSsbHYBJSbRHg7s0xTVc0x/myPWgE6Bt6iPeOCn
9rEXA59iLAsn7gVdaKSKy6LWLhp+C0j4vmputUdA7Z4JTw6rS3pEQEXN0DSNRQNg
ni1bVSoTOPfT0rSfDhpgbs9rSDOaeBeoaqvoS23vOD5hRAoHpACMQeolpwEszS8D
5mqYjV0AwDYKY6yGdhIoAer/0N11YJE+aC50DFA2VLYPDZbF3xRYYNKsAIQoyQQx
Zzxfh4MgeJt0aB9WLP9IE68Dr8qmg5JiB9imxUHt6BakZGZMVE45fgDCSE7ZDent
UM1caGW48Cl0T0UzG9FJLX1/2bWkwdoRD5ZIXp+DMzU+w+x+a/lkz3alyV5EHrTo
68FqCogWIlGwSt6ZkK27sQSwBMWZHzBOuS3U7TIhwRk0mdBZ/OYtGcCnCpgWwCR7
9fk8r9mV+OkK0BU6cd/8uxcTc3zsA6hRjk9GDpaP26+5xrzoNM1TOEE5qi47xUl3
zkKA3M/k6OpEVG/0to42HLvhQvXYuH2Oy7S/+GM12WCxT7SLpTPf1bt5csfAN1cb
8BJK+/SKyqiT99CvN00/WUKFVGgdFy1ttMC/qL2e7f8Ib6F+vZk7EA4aRj+r+ZHX
f10x88RxGjZLXgVE3sVj3E20o8vLfl2zuP2bFBfWxSihhnLCnGJvHKQjrtsDxBv/
MI81CHW2abwx4OLiML87GuO/nqjFdre3T9d5JnvpenFIhqgPmffzOENx3GFxEXAk
sNLP5xX/OxulBtfzkNvDaSeNiRskiGUJ1aC+K7J6QrBaVIkVU/jh2CVHZj4HfRxD
NFhxa6zTwae0qI1YOcyAJRdoOQIOy70jfxEnEtgRIMMPgIOgWAoetN2eFTudkOJs
jWXUUIJMm4VuLYrLBZx7UzoUTgf/g0w/HzM2hWKIx3iz+FMV3uvBuxDTCsQLXPR6
Ge87Wj8Oq83R3IPpfuGZ/jvrNj95/vntlj6/xxSJpzsjOhVXQmt9ho3vD3KbZjYM
I2lH0vTO+xUZCz3Ucpcht2p6dt/Z6b2CVY4z5rWYUxYUayXNVTpt3WWoDrhYOZcA
Xxbu7x51PmfumL31cqJAIvNX+fDB1FefC+zzenzktngwkxzymkCdRGJTRnPO2xVG
HcIkbJgimGFQe5vDbI5KzACUrSkiyvwpFlEiqtZUF2JifOadBx8zVhgA37gUq2Tt
7GUn0gu6YQssD/ua/7iu6DeIgKQnBjgm/05bUtJtg8EMyNE5s8jQoQpva0BWrNlH
BbY1PR58naIe0O+PmDC8a9HeSZ993hvcImwswF6B7bmtKkIBF7oSaADVzQ58G1Xw
X4MUlA3qAfK+htNJ9ZNglUc4740iTC1SENwFFfgXb1uHR4Dy1cW0dVOIPXDevZdj
zM80bqilIQZpPKAIELZ44dGdIS86q3WIRtrtjvMzatLMTC+Am3ARdOHamvqBRtJS
9OczseXSMj5fx1CCrXMyzhNa4j/8YAS0uFZ3Lp9XyzHCV2NQNDMeA1Kpqb8I/FiH
Rih+G3Y2kakBUmeV/x+UTCliI4cYvyMRGBNkxmKWK+lCtVYfuNjUBddZKvhbdUJh
WipdJlngzdrtD7OCTKuTonn6FlXgI+1QOMdFzyEiMY3zEzI7/CAl169b0feUDmOr
gZiMlWPSorJqwnf6bPxcqQ44Lf62bxdhM7SfN9sc88l4bglmLP2G87OZd9jEhO0J
mxtuPERz4qWdvzEG/eeJlHj8HnPb9i8uLr7wyBsmDVLIKal1Kih/77RT3xmo5ZjJ
dxUDdVyu/7P1tXCyN3FbYfOUzr2itufkv+jUEofirAcpN5esCiCkqLbOxxFD15r5
uuu969DOxrcnx+hNV9eqrb2Jx9XJJWgP55W5ExSmgJwSSckMZwQx4LbPu4iyngGq
50JrdrfzLFrfnnNNQOTb7ylyBQDlap9wME1LndjyA3/3oLLO2bPSzWD+M1ckgVEj
bL8xaICnETc6qqRkgfRZMVLDs+xbj6yIGKHp6tRTB/e3dDfucIfxee/3F0SBi8VX
vc29yc1drzv3wG86SlQNEDfAUlWnl/apX9Bt2WBQX32/6lHoMb17/aDx+tq7erIf
y3quwAQKMXK2tQxWHSTpO53bQs5CkacB/1BKzVbYKM0iXbgmW3Qzeb0i7gfPR/NQ
EwbNhFlOdOYZvFqu5X8k80cKuXpGDDdTocRnycp/LvYBfu6ulExsTusFuWvn04PF
3Z/Lj5QU/I7zE63LM0oREfh7MDYMeGLQ1hA0H96Z1apALoc0hxnh27JKnT2hJgBe
a7GV3eo58aqi1oBIrLOWjcdU33QOFDbnG79dLOelj3PPpOTOKp/gGQF9Y/s7iEop
B19nmM0p9LUbF4AZkYKYGCoEGfwS+LObeYB1HRoYQpzztx8JwnAw8J4FqvEaOH8A
kt+runT9h06YgmAEPc+4/ozb/lV23vS4GOoJCAP7xzOwSJHqDfXG+YrxTXzNprzh
G9gzlAjHbMuuA7ucZAKPGUU43tGCScfkrNzeOl2lEYuqHdIbkJRuqfzVt7DVBfH4
lheMfGnCorJkRcDJyCiWS0gkmpY9iDl0SH4QZz30ZTWhUwOWUwsgK5VKowG372aU
PwuNTVjmdrXbCzJBLLc3n2P+bu1qEnUKRTfyBtzYWiLBz0tCHPyd/LuYv2c/YfI2
EkFVMa+hh0JRD0TJ/TDRe6YhHhagfsKL5FoEGqDcjZ9qijz9a4PFcNQ8VnToptur
z9FQDGlIgwERucWRJax/M2IoQi0DdDCX25D12Jx9xCfiSHUjSaPs4TOTmBY+1U7y
CcgkIeywJReWIgxpxMKF+zd9+iRMT4qR68cXPPtwg63BqSl9SyDyzLftPwcCmGp0
wAqe6vh2llksaKboMNi1OfGeEI906HnapB1SWHz+IbdLH8d217WSX3Dhpf8hoK8l
KgXC48B/6VxcgoC8sDNFtSwwkdqcUU1xIm7KtxpSlb4ANfIZg5OiOCbY1ayJy1g3
seZprXXaEKG4kceGAOxfRf2DjrmjqY8upYcvdCL6Y58Tj6uAKIKzQfr+MeydPo6C
t7ibHnf68uFc9hoNYIQtHnk6OTWlk+9qvgl7m/EGBnrP8OO3OF6gVMjYUMFXaPtp
8ghS7wj7A+IAolKoq421j0GLTL9mj5iXBBWvcynoGT5xVULP2X2SYHrr38zaPsg7
/9mpYyzLOVLNBQtjJE2ao7egouRYZuV07U4AhQ1cEunhjQ/OqBvn81i1gkx16/Eo
F2xxHIGM9NfWaCQL6+fmsN/qZv/rSSwJtsIAffKp6QqjnhSUVELX/YsSJIfaHQL8
viOU07bqgZVACVoE0jR8ODpkZ/whWTEEx2C62zPHYL5QXrCSF+mihooY3ec3nzfS
BY5jP9LCx4vktAhHujTHy4wXxmZS3+xudmUWKmYjjAP0mj0NyIsq1BbY/gIHQviP
S/huKd0ZbLQ3pMkZdvod5b3LAXZ753UX8VET3kkFYCvDSqx6ofikZ09kDwY/qi2n
NTREGy5lwbm3Rff89Jf2B08r22gYT5sG0U6ErAqpBjvwicLc36IWHFCG8ATSfoXa
FRBifg0tCDnDiXu28u8h/CYA1/m4yHYt1jOlx5m1mWOoUHK4gUj+6kS3D/28LSI9
D/ZutZzlluKO8QLr4lTVgF6dM3IS/OwNBdPUpFzbatBxTEIsda88MQyNQIN20VFG
7yhQ/fc/NGnMQm8kgKWYQg00S8F9MwGTYDkUk6GhpGo7DxbcajyVCGCz7V4a7vuE
gHOsThPr5HnAiTgRveri6p2a2UY12WFxMp1dKpJserHjDGFJ8KKNp0MXMCPjVms7
TzlcUgXy9YziiP31TfMCXK3UCqwb9Co7HLB5PWUCm0+A7BLXvJX3qw5d+0ZvNtZG
BkmxwZ1Gh9QqAgVWNj6pSkvD6AZW/XqDty6kT7Av0B4NBUUyGkwh5o/VgOZgZJXk
ogDAbNpRlK1Aaq5m7n7enjhGIsbiI2AG72lAlMytR2HHsssDyzofAjxY1W68H3Jp
nxfxpqz87ivXoVho9sNVjQHxLvDm33A4RKp15pUhsOHqcmHm/T2H7UYHqxji1dR0
efr8Maj5XrayZXHcVY8Y/Fhn8Zb3XkWQNFK7bKTBcXkgCqnzM01oGHPbg3W0+NCG
2Ha9aYHPFLmAHqBOApVr+HOrjx/dfgpUKE13ICokT1WOpaPQH2IevUoYJhH7ZNIU
ZDHj+RfKHUi5BFANSOGGy6swFYGv8N7YE98/QHbk5MN0+JI5rXV4Cqdu9Su7IhjL
ks1T2VzYuga06ehAixBInJxapJ4raOQiS2Evl/Qoet8elo9PoINwZB7j2P46FRDs
iA0LuuVC7XzGkGVKhJ9qCWZ7VcnB3/x76RB3I1Hr09eHhwnDyKunSkcjfXW5vGn/
dzht5wwDa0+cfVksgMWxRO/vYa8w1eC9gWXVysdQuFaKK2hj1CVlVyprXupBmPc1
+Bs63/vWHI6kzmV17AfZNvUZZC27zUR8ypGPdE6VPtnlvE+7KhG6gBGulMx6WW3E
mHW4cYtNx+wwyd8nsUGh+jJgH4ngbeSI1n8F/Xr2lef6zlrZFW6npYSojD1HCVDK
6E3k8ywzUyR4nIbBLdb7JfIWe3FJMH0YNlhUbN6MmAhoDYsVwopGV5Jevc4QAPaZ
mGvb6WtQkDzhnIvoazcSMlH3tUkRytS8bHVAkKxKuCejdPXpHLlqqkyTrK1BdaJ7
mv5ApUG0/pvyTBiX6FkSlAmrvLLWBfp/Hglp1lOzJDgoRmUiHGh84/Z8qMBSBXpf
xFFDwQNOufW/o95WLuqbUchxKiKZlZ4wiWPcUrmNudHvd7eiBTiG+mOtCJhd60OE
m6ORGlq1wH4T3OlcICiJc8D9BYdWfHnvEkl6kL3PkgIqSyYbRBx/Z6tQraAi/2Q0
rJWIiSYyvNdlz/lv832b63C1soRpwGmeDkaRpcG5MyR8GewBe/nZJ+iY3dEip81v
OCEOeusO5UM9httJZ9CsOll+jQ7kXh56U4jhf5chr63gwibP76zTBMMsRQtQYoY9
0E8LJZ9eaN943OleIPs4U99l9ZTxSagFGXWJYABnYEwxXDAmfnnCFMz5fgUm2ann
HuitxTTV7oAgtZxlqO3HULaalT/w6+TCEa5KXRlkQxT2WVry7LuJdMyt9rpZKqwq
yGjTL95Ab5jD7VS4WGNQY7XM8Q3qgY62uAsOAcckpWwIEHiIIS67vKKDJdUdz84Q
bGHhsyXgy9fnUqrpYxON6xhv6cRqh1wHyTGiyFxDZhxBmKsFmFJEntSzI83e3fCT
oZIxhQwUi8EB/muljLTq8uSbXtiNIV8e22RY7FJnI75J6Ik67swbb5/ViPCYJtEs
W0cPX9LSm+7XbklHaXw2x8cP22rT5zgeQRKHzyx4Iu1yCFJEnT/0yqlfn5Xp452O
mbZhLbmjyAD4yUEXGf13wOs0tJvmJX+8AFgvYDFQdXBGGc4HUZ1Ne7s7Z+3sgb3d
D2+a+8gVMGMbgamrRpXu1FkBLKQi9Nf9lsPpqXQRnbdKD3VMaQwlgxRbYU6fG054
eH25ispRo7k+Uv+JDtR1zfwHNJDrx69QW96zYB6EQ895fZDdh4fKlGnl/MGzGsfd
my1vT2mPRQ/2k4fjGXuJwvn14fiREl7e4wOh2eAy0B/+Ym5/kZhuF6p33T3bV4Xj
nYoC2puB6T1kZ357VGDNb+YTnlXKPQipGaWJd3FL3eGGrrxZ1MQRpH0rYysIDpOZ
OgdvOM6vK9MIRpuLM73FeVIFxCxltb3+2URhmhbzoB79mr3y6EUpEuSR1JdmX8DL
3V/YeQVfZhzKijO+tLixwfrT3VLBQt9lEZdv1Iuc2u8AHlsuk27TW2EUnnrqIRNE
AS7lkqT7ff8TMT73LcFAQAn1B9ESgueRgkvdWtomYbEHd/X0ROrGdVntSZtZn1rs
A5/XiEkug9s6dGq5glzJAsyF4RD3fdJ2srY6YflvhEuJ3z4zU2e8gYGJgp3pQtcD
hJPvMtkdgI0EJafU5t3zhUZm1boGTAtir2J2+f2K72cYOTeb4Yt4zRBoK13//jBf
noX0/xAzkGSCpLxP54ebooOIGQqFAmbb4RUr7aHtqgy8QWuUQbywpZfV1HqYIUfA
wyIWgS7bR80/yMLFNzWmtj5/4HC/jK0Qe1VHdvb2nTyET5OEAMsu8on0ImFmF83D
8edkqnTWtg0me5ECcVbhYa8W1Iw1Au04Vup/IcgUawqKjWEFd6u3NQ10RnKepxwL
0cmDLlmuoAtB7Pbspb/LVgUq97LNBbpoSSqbCF5i7VjLjmPVFSAjkrfxAnixf82t
vXpBlhyycnYL64V0XfHKmSz6IamKNF+FNl/d57MSSrll+FndVgT1eRxywxTZbobz
cIAX7TPVSTzYV65Xia1K3702IxX9gmHd8/kSqfYEUb0rnht7C02wAnE/BYLEOCPY
Ugj2gsU6CphKy26EwivHm4mmu3KVrxtJvB0TOct+pRGDMICAzV27DUL9q9cbfKRh
6XOXSnS81JVn0DjYIZsHd+BVPKhgLlJJrYDK0+z6BnTNebcMz7PB0EabDyzCRqz5
JJ833rqfXjiBUYwedf/X7uGK8ooXHKxXSBkBW2sWgDIL13dsVKGCjQfxoJKM08g4
zOuNDUeeQ913WKiE2AQZej8VloBrQXqTUwEejcnS7iKhr2w2+6FGLs6GVyVsQfmF
8/r4khyJVuRqJrVrj9GFI0jMLsmC8OMhZvqG0meSmZvwbYdSNTnMdIq2+Jy5x4Vu
bP/gxboGCD04PxkRZOdAHaykPuuR9m7godpkx4qUoB/jlMUFrld4f5INkjgY7JJj
Z2hCetTsaZmpJh+G0mYXuj9c/ynpdfCVSKbdGBOHJeiV5Q6aNQFXZ6Fc9gewC5lc
8sG310JaHeF8ksuJaYjFQuz2sbyQlsTE9EDUHUC820yDdu/WzyPvCC9o1hMAi71g
57VegSeeMEi+L4IFT3hoMDXSJUnYl3Z4u384j9YlUeza+fkYRPV03MD/6hDwts/B
PKmSvs9nB+NUh6gMfvP8c7Gz3Rk9G3A7m4JW+d5M/Ir3SezDYuKkxeWGqOO0pQrT
Ok9UUs90yfJGhZcYM5TRvkjNXLyfZDFCi05oMU3tloi0Jx+/mJFqh12l7SY3jTKl
Q0jrNOMhpLmEljmqHFTImph4q4xVTVApM4SDH98Q361SlGz1IUmuipycw2uhU4b6
Ch1YQKWWx5QgAWmVij6sgulmqeQKrVDZbqB3LER/vix9sjEudOdjfc6wpyBR3sDj
UsS1u2UpAEucY1lQa6gGzKxiPM7tOHsXAChOYl+8HyZrH5kKnjT5FCVlwYTU6Zz4
LaNwsVzq1zs7tHd/ejIyX98sEZhSStzG/b+B9HH8lGmDrTaw8q++ZNX9+vT6+0WV
WlVCBEBuRgHczTv3UgiAG9p9DOnk0oV7skhqKK8ktTBkESJAWyoxAXjpyrPQ0UiR
KTq7NvAvnqKWg+yj9ES/m/KZHcrUnXByywh+53Im362fNM3qHAvfflXTMo0SGYcw
vFJ2RRaxIrrR7JexAorMSYfZKdqLL6ev9B5M2xTl8XjFhddE1YBuXEKExJiO/OU3
cmGSQwm8dQ6qc76HUGm8oAxkl6ZYtVz/KEr30fkt+E3oIL8dKoTNZMq8Gi9GBA7U
nxqvsHXo4y1e1FIHcQfNvQtHrXsI5pnW24rreCQ2gPgKqY5AOWZl6pYAyirA0ku0
u9iI/swNKtD6zwpACgrdmVq9RqkgR0T7aIgAmocWhPWggNC7/ZywoKDrUfnf1937
SbB3ievh9yych1xvwKgej2RyxAEaHpwgv+m+olXlmYkR8RBNkYyBurY3voA2CMY4
C8V9odoCr4Lycz0j1eyFyNpV8Zcx9CAHBkFD43Eyze99UesdTADYqtUGDn3fb11f
isXuc0HMptJcE9cgKM2xcJJynwDYGUzREQJJVZH1KBT27yqQn9JG3wyjVQ842AWu
QkMgtIWsxamSfqfTfl6tkTAGT1P/fGYdB0D2BhGt92babzvYrKw7UPIgknyEqK33
EhPpKurVOUFqmYQHzIbL48Rzws2qyfBLgWvHCkURxCu0PJpxQFmSZNs9D9wUXFu3
qCJSORmYKr1QRgD90H7CACbFX7XiTuC7CsISBTYkUq4+OrjqwhYAcqUmxCYWVa+m
a907Gi9mgYMhwk2kmgMjodoRIB7+/U89uPcqFEqllV3MHfkpPldnteRXiI0nxzbd
MCTsBc8UKpVjru7rFmgHRMEpRkqqRc9mkNp61+OK1SMWuq9DrCXwm50U8LKXfiNe
fj592LfNlp/nsowcCPzkRZkvGSQEVoP7hlps1qkKu7yF/qao1CD62Zm1Q00VTfVn
+XncuGgTKnbDCR37DjN0WAZtddDmuTAf5Bbo0QSg7sIB9/bR3l7iYfHbUpC3/iaU
eFprvMg6W3cJpuIGTlTuqd0Nw6U6cDcRwBoMl5da1MRtvhAS9Ha93sEndsFN7P7u
eFgZEU9zijndGFoXPV1/k8rrz3dpMeZMrXPqTdHZuclrb1bDthOH24oti+NfJllC
bcOpKGIcwjwmDoQPiPbfzecDZpPWoiVDGiHrDfYmEYnPWpEuYP0oT3HRcfe0gGfh
YY0R75ysK7d9XjkTBjUrq5VCjW5MIzswLPOTLVj6WshFm0Rbj90wQ+dc+k0qRxtC
bmv53SqNkssCIiWu+AW6s6Oqry+90GDcWGgOV4Vk/62SU6v1GgufqJoSZ+ksCXj6
RYHyM5SCo1QIoL5bSR7draD391qNqdrVRb+wpkIhXUdfevaqehpjj4eGsBGH0LBg
2B49WJ3bFjrZg1oUaQpekVrTXVFvW7ty449uU72o7ahXJtDWzgFggZVTQGJVj+uC
Aq/NKx5XRuZhPKFKnByWwd+UzvV72vY7b8L0nZBOE0S2MwVC72/tP5jiVoIZgd37
IP3ECkC655241+Gtxs9s6BW3vIH417ko53PKHxJ1ArH5kNDLKFQbtv+laXvTygVw
hWs8s6fIM6ERTH6TVnolLjjgZC5U5xdPvMW3b7OVig34dB+B7eKl85/iS0FV3Ewu
uiKUDV0Wwn1lIgIkksZW4xKn7S+bdaLNj5XjKEMbq6HDnZ42Kon0DI8yiJNKgZgp
k6xfBhL4W9RC4jPSbLcUUuO/hADoPoMqAwmiEGZq+SLU4WZ7I1/cZado34b+W+Uo
ER4IAkaIkqVcAjORoTWILUU7sXI47kblrjgrfhcgoaMTtYWO8pSjEYvDil2VodOw
72hkvetnpWWg5YHPf2SnIeSchlWBn7XPOX2xfvMrWri/JbsAi78F+1Gl2vIdFEGk
xP61LWv11T20aituCqqd4o7/gTq17W+rapQYBpFrumcKh/SIuUSdRTUl/S1Zl1PT
KN7M72rz8U0woUBWphY8cTsi7ROYExdjgBKqKt6+P9LP+JL0JHkYohoRmz28liQs
F9tnKF8ZguGxxESdqnlwom3UHGgtin3jL+h4es84/nRGspkTNsIYY5Z04kCe+Q03
VjQQw4VH4iqsIAUjH3O9zRvs5jSQvVTZl0WaVhnqA/RWRh7wZHVIVZ0WwlV/csNz
Pz/L0bcIVPMmJUumPR8P1Ch2TfSpuC3uNTdqaV/MO99KcnGlTcHlkiiJkTXMLOk8
CPqxfjFTxNk3TbcVSASNg5NBxk8mRJFqKHC0Zy9Hbbnosm5a5ASNHj2xdG7+Pc7y
pfv6+hjo8n2VvLzOrS6bVnI8H6fwlEXmQVNArJQbu+Aalbq59i7fJ43iD7Jl92+u
I8EoqS6mlMuRpC7DDfITqeuqK0SCXGLkPIduBpOdK2rS/IYePC/HkDiWmbmsE/1C
8QdrQw7PKrwD1Dy25RzsipjQhlt+h1x4J14wxat348v9mY56Q5AwaNrHwHb8l2/k
rPXT11gxkXXABdJLMv/lD886m9u/7bT+FMUAe+fUWMYztCi2fIO1iK+B9Dl4dIbr
8Y0ewwHkNXXc84uwQftrwjsqJo1GnEZlUQp/9qJkVwIJRbKqeUsglPzrpw0uvhSw
1CSOcNtBDU/oWBGEuuAVn8yuLFwLahPyJ1SC25HcwV+Bw5xpNTtm+8xNOXwA0HU+
OvgCvoZbNmKlxP7biXCUKHfHEH1sZ0IxxHSuooz7UvcID8v2LkYK8tvpsccIP8Vr
FIf+NlQC0zP/nOdBR5Hi/SpUTqCR6DS0GgI8K+fJx0YMkE0th/vm+9MeLOEMfNaI
Sl8ZlcmfK0gq9HUDDnn5U5EKzZnypdpGGrG006i9RP4iQjWvs3NnhjRORty8OwN0
OrxVJjFJD0862S7XtUOr/VGdmtMvEbLLvVwUaVgmz2pnUxOQgPqdENGaRx4C8FCm
tSaD6nrIWZz8Hf9vlLe594yWEcw4IAwi8S9QTcmmYWs/0HclgpzdMpkjZK3a11Js
osryMQJY7Y8nkaHrbw5VDGVZ1npw6UzqrHTaKwwra+C4cR09RsFO+3hUVOUE1GJ3
mrwW8JlzL+AmRvjtoeoOsQF2zQQHV2V5ODYX/oRxv9Gw+B9Wn5rgWyG91X1gWg0W
LyGauMnSU5uw1TPeFpBdpaHyWxQfJd0tOI2TYnE5knMdLjSEUJoK75MBAu/2YsV+
PT7FfEhpUqSaUCeLgIFZBTRpQa9p0tNQJYKoWlsYBYPXAoB8fDR2Wkr4whGFjOCC
36zV+nnHb2//RAHoXN/s0miKngun5D/h49RXqj6Gth/qLOtCLUjlNHwMtX7OwLnX
yvgCQdvDWos3xPFc7E4FKOLIWMgTzpYBbX1ezEbp/UjAQfODt3DKCC1c+Yx/G6cS
epT1R6BKdPHFrIaKXqhCVH+0pO9rl4UBp0ObXuA1CjRdb3RbRCfXQ0L4WyQVHgAt
xtQP0mTlRq51guLQ/q2FEEGoPZjFfoNvFDxCmkLO0uh+RxbsaXEw5il3z8Sf04YJ
wgokSgjIPgTEn4QgYvwTLzpXMFBVaqci8g6vyBqaf7x3AKx5Q7o3RVQI9/jxXcdh
nuZ9kunL4j4hoqbYP3G3jSYKDBOwCjq2nvRjNDV63n0/qhvZRgy1t2e2xvsuFQKe
VhvFJ63oMy1/b6Mbtb9Tm+WAPZ5/bmgfrgPAwGA9dTk=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFqXGaONc8AXxJUtXjgX2SgmVwW21BrrR1JXix714zqJSkfJRnwvOjjpGlCFphwm
g/LNt6Z4YZ3/WERaCFaQLlosLQFI0uLoZDdXPAwCYG/E7LuNyMRc6H8Wu0/iLqrh
dbQIamu6q300ikOqpjrknIa7J2wbxmj+m9AjkqTHQK+1bt8lH07pzIHcAl2l2DMd
fFrgEQnYCKfET0+bPvb92tkxgtEp0IvlcsMrm0qc3lnEWl4NHZGckOliLQNNpm1e
3vFmnlDNjS7o5cgH389h0s2ZDhvm5oVJxZk+nYcevqvoZeI9mIFXZu7+Ekc9CqqB
fZ6ZLYrjNnF0eFzvJzczyHhUFvza89SDHMFgwD0dAL2Eg5FLuwOnXd2JMhGJN3gh
DXSpU44/hgqORu8vvkPDAcV6DHMgEZKYWOLjjqyc50PijQzrShOctcQSiQ7x6h9G
6G0KF8W/CtVMN8Yhgz+ffeO/7UJ8wG4YMVztlUFh1MHkXJ1Hpmjrczd5EN0+sA08
GlsAUpdkSjz1tJnA5mUWBBK+FLMENvivZO8ziYpAhz6eDuRolfWm1Z6EmLRBnaeO
AV+/l6aF1Dl9fuzNNosflG1jqiCokxY3dCWIwZtcAnnj+Y6aD2XCqT1HuYHG6f6C
5gOnrxZgm1THjq6htZLe0E3u7bmXVy2VKCMgtN5786CiFOUlc5dtofKqLEwvlw8j
PyRKOhIpjgt1OZNDgXxof7jFDN1E5OnBZv/1q96k2HQyOqZK/UNkPVTqTl31bhsh
xkhzqQ2eH7R/r8EeQ9xOWu/zfAo0gTZpYv2q45VHqobpPXJn1F5oKSZ75lpVbG9Q
T18Lh2KyW73YmbO+Sh9JdKv/5az77p8iUV3lCqzquUYgQHI4wjENPs27Vt31r1T9
OKt5+fwPZ3/ySp9cNmlo5CnTxDOO6s3thwdMisdpQjQ1vmCVJESMU9ZDqsUz0Iu2
Pikp3VDJAOrHnPaKEJtbrIkc9bnDn0V0zxK4A3g9+CxHGqhPqANqm0Vtv/dyifZY
BVC/V+pETG9uSUiy1i8XAKzW2XQ5n4e6iec9JIUIWXVFyRam4TuuAWtLzLKThrS2
eTcN07llkeEkNsKNfL3sQkMct5+Bn+q+lXacOyZL6974RPbI88VZxS2fifaMIRzK
0LtAXpArk2LUMFaWWDli8dgKuHL/Nc8kNnXRcha4DnA9FDAxFdygWuNY/JGtCf3Q
1anH/xY+LmM0BIaLPn5Rn9qUEYNnyUa1v5usPYiHe6X9Q7PMghPvK7hVqeRhKdnE
9/UWtFP5F7RPM8zOB6HnoTqp/gC8hPy7W296uJBBXUn5NsUfW24TLG9shPfxWXBe
ChgUy5CKhku85FlNVzCpE02//RVrhRWSVPi/uXhBSnc0y6IJADbzyPdUKQcwQAnt
/DwVN5B1aB3oNEcVzAHPHuQorZtjp7UEjZV1BgvO7ZGmp4cPgvjy+9WJEH6ZeuBy
JSEqc+1tkv82vk2OE7jIOgqnw7PSucPqY3vsFf2Z6qe2t6MoiyGKDZTK8dCKbBAF
n37aRmWojNujTgIDr7fDbDwMO6Lx6q5IU6MJ6AJgNxzXcEpr6PJFHkTjfYU86oN2
MtkLMMJzhTWIUrHOv++MC3hV0cdMZtv1oB8XISudZOqO6ZIeIQI8NuJXw9NkT2c2
hp2TwmhBOJRp2uHiDRG0i5Ij7U2mTZFRHroyVINZ5dMQ51n9lt9rzbZ7CkDxlsrO
3Cnhc/t1PFMrH1i9UT8x6Y+4LcrfIVEqbCjZrWKMwXsyfnR14PAnmNBg2dcLPb+6
rn4waYT0Te5Qv62u3iiwBC1xToz0Co2C+Rh0uSe9sPDyuqNbL7AQvv2jrsz6kq0U
lM0Ihl4Dx0jZPvpuIDaOS/+mGVca+e0/ygyHtdmUWce4dlqvfwOBqZGZWULz/BtN
wDUHNkLZirxxYKFJdiKc/pXShRWylSpFSxCyP/nZCjufiEXHAdQ4/UN/hhuqXON4
4rTIS+ITdO9c3iOVnBuYL5/mQ3Vu2JSzbIAZPoFwtDyYFkrx7MLPQXzlFnVCL46V
b0iWgtH7ZOWlknngGoRd+VvMeoLIrA4ZQUSck2erZiO+3UzZpeBUzpbY9yp7Vcg7
tGeonXIAE4L+C6qN60PK2w13lNn6iXRwZDiimbpZNWABkcE5VDsTXYCXTBX+KwC8
eYlL2b0rDWAGscQOJ7YxMdhj4NhFjPCsyLCpg1KY++xPTOIdi1sj183V8BfXnpk2
zZrmX68rl7s9HAun6MiaHl7MStDsWfsflIS627NlFlcRnWiBWShg3+/ddcY+DMoW
R0qKTgBjTjfUbp2z0i3Z6RxEpKmTQL2iqVd2ugAAEUIsJo8bNmuFO6TX2ZU05CsZ
tVOH2ify8LaOOPe1ezbyFz+tHu0eMszVOJISGwDntZgjZvBqpTFO7oI6DcB9sjzn
s8wr+3DJE0h+/l3pgOFH2Viw1+kvU7KQTkJtdjkmuWOs/qgCivDusKguT2/ZTzjf
q9uU2dNLx4zXlrkQF9atiVxilRIi/HAsevNK4bb05CRzTJdi4LiEQFKLcFLtUNIp
6ptO736/10Jo8sAc1LQQxEngBqJ1QYBi4v2ogKi5NmDpj5u8fGR2ktd6PdbCYspI
KFuRw1VtMnyqhf2tgMbUXH/eKbvdd+j5TbRLzaLJXr0ggvcuoQ/IeGGnMfgnv3Pg
jeGfRoroG33Qub2Bcq5K2cbbIHTdi+ViJsmTey7joTbT6fKj0i0kMPFgrsII9l0c
H3TU/WpMAhpIS4gpQ2tTC05NYAa9aV3L9loi+tikJ+V58h72KW8jt6Qnto90p1py
/yIegGgA1Jw7Ldtpz5yaIbTF4y/UxWoxiDiQ+mK5k521Tf7kjlb1Z7oddAfuLAf9
ZECymDvCqEYCHV0cr0htgdnjnBLsTYt9QkpPBfGge/vPQs5977JDCdusSjEEBAI7
7A4ApsY++6X0SssQtvmRwY91mcf50xThC9o8ZpboHUJOGvygdCGvMtVzD8s0d4F6
Eb9usac2ZVhnQOxtaBwok7gkzPkqyU3SFUdWrNZRJoi3bXW2xZxi0K/95ivVA+si
bbVIOkCuwXEsO35lFPv0EYDD7MPmVnh0vFfkMj/FsJpbhE/Exb25+DTnyXYRu7j2
1MIghUyXzqPKoOWdARs1HNu60B19ffe5avco8L8LbeocpsYCrFyTV3G+guOfizDj
qgdSD9KOfaz3A2K2j2Olsq76Is4euoPss0jSxMqgSlPW4gNbYjUhVpRwHXMedrj3
5o+Vj7Kws5j3ums22T6skt+jtlzwb3AjQftQ5XG33uTnM7Q4vek9BpiN63mXoXzi
fdNoZbs3W3+FHwlgLvqMjZnA1AP1algnneD0ZPxXt7ONHki+4ciZetbwqS7MT6Kd
pTU5rhm3z/fVXRZ/1HtjyhO7m3r+/6+JuJWTHlyWFN7/zMW5TunbwXpvr1yfW/yO
j2fBmQIEqOHX4rawGaQjfHpw1oimBJQO5MiigztvlaOHrt7swhe6DxDAt245GZI4
9mfLtgbI0mlrCmBzAzAMoeIUDTcdJaaN3XAUCjdw+9H7VydyiavXP4HR7bEA4dsT
PXW6eT2tjm/aHSDRDeJV1raFnRHmgnKHIDqG/3vRFXziArK5eh7wL+i/5J0yDX1E
eV6MiGpNyfPtKs1tFY9ru67hoMdzRUfAzuOpk8acXDkPHawoyNK+iValw2K4x9Y3
+ICyc31QoFt+Z7GgdSDCSo9kkAO0vGv0Nb+L1ccu9BjRDEmXP5j+W0gRpeVS2Kyl
fLL45lzFDxDeM6J0gz6gmCak59qswxLhHIZ6cZDuA9L0OxeJd16U9W7D5WemwzK7
iKSgm5aps3NeiIFDxFCYIWSCPQk36ncsahx/QNMwLIuvEvyiGaLNNU6MTsbThvM2
Gfup4PyBgadYHnYnImLrQ+Y6wLNQUSvx87k81ywxlNCD66HYrR/JoZkOj/S6WgMR
1MUsn64H0hPh5F9JsXQIipCWk4kTwprkCO7CJtXfAhQ9nDtDy56j/bLqsTwcvhv2
4m1OUxNH0faNnwG08mftsJpRwydOSQfBXMSaDdkJYH3M2qJ23M7hJjeozZXvl3kK
ZULoJDqoThAmWjirpdhpsJB5qIYmg7ZnaQfcrqzgG6H1PU5g6tG84rHd645PFfga
StipCjJuohpnXXx8vBc22MTL52xx9Df7jewGZbNIFBOe2x6y7HFlSU8E1PifguPp
phR7K+6Bd9Zwm38sjYsWlz7dwBkcR3GpOlq0MVpZCrlEabVNOAu4w6qwkMJ7wTxJ
pNQ6DhthBNL2x2/NVTQIkLZl1nd6zhr9D4veyiGy1ntLpbCzB5/Yxw5I7xjaRrIO
gTrKTZgP2h0JrPwgoC01ds51U+J3OSvJpAs4H31ak1ZMvhlTm6ppzBc0Z4gAJDLh
DE1wyJr3lPAZQlMTPKF1xQ88p2M/tzl38XzBj20+J6rb7vY+j4IXGYQwbR/2KIdt
+0SCyictH2fjhsn1e/UWB+ShnNzttcQ1VXDv7CjDA5yy2DcxyxrnoQqhicsZk0mU
kR60whS3NPkzGFrefkFtXC1IQjD7eUa7HT7FZMwa6RTcJkxYSRX4CM/q2BTjj2pi
Cf87QFNZC4I4aW3u3Zyl+jK2widIVrcLasJKgNKytxVOTlTA115nF1vQVQUl0Ce7
KrqTwD5H41HN/SabbzJvKL0+CM1IG2SNM6yXwoBmK5cMu1U4ORF2kKhbxTfO16+I
jrO6zOdbkjGUomMTMqO7zTEZp8bVUgtwGOvV/MQR+VhoLiTEexVmqTw96uD9oUZQ
2vdw51v1yrt4WI9yclpseqIyxBsVMw9y23z56g1xN6gNWLxAtUPrfUGHH68baWPw
Lsrmsk1hn6R4NAkpghkihXMlzYgLtNxPG1lSfUknoliMoAviLdDD7cqOrMzsIob9
OIAvcOZDa/RApqTMUs0Ub9Og/LE3+5aTBhz5c7kiff9Ye1aXowgD+YPcqH2SkrFv
Ss6GumR1FFArhOj8qTBHd8g+PI0L0spmVZIZI14i3SzkgIQOx3A88J5KorXnKB3C
8REsw0mcPFbzEvdPyfK1eCVkSNFwMB+BFHQ6VaeOWqYFBO5c6CcYJZ8/GGItCbH7
N/kldlWFkJcW8AtTzjuzlCCvZBvakrOSMay2IKX3fNyfqyiH09MKw13nMqKy2YZ/
0lywQ60pprBl3HRKbRnDgKVYm3a8sQDw+pSjeTHfHMzM51u6uGWhMDNKqkvw5sxm
WtgHGr3eOo0KtstkUf9rDFnJUvcizmmaj+HkOjil1m9Dvn4JewncEWxUH20IiDu1
Z1zrXPsAwQD74MsscGgliVyIQjWt4NOdCDIg6Lb2UhdjnK5c9JUlaooEc72/Dboh
7g9CgcUsnjAxunvlIpHbthjyNGvt6NOJ3dWsP5eTN6ybxYlcYIat+3zNaKLftl+5
KyNpXgmFK7vxEZzP4zXTk9EFWjPB1+q8SMTmQBv1UP/g18oDdtOKmKEkLLKbtO9q
911s5g2baxPbZFZSpp9YXerO9QSqxtIqzyRdPV/oTO0x5tLeGPHTzlsBpCGoROll
gKYx1Yh/w0Rjysk6uSc9Kx1CD8gwviRlK4Olq4FwDa8FPG1qmOMqgC+P9bMIudaf
JygNjPwqCtlAKbK7V5noCCbmXqkzs9MevbtltWyO9VAXQdESCejRXI09QMZ6vS1+
lQ0fd03YO3aMuAmyCz4kLxIdImO8f77Fo9uI5FRgOG5EyBn/RkIBWk/DC+kCHY9I
5bome6lCWtt2IHvMnuLUzJlhmq2z8oXdPFBJm94VNw1CIOE7P2hfHjIQj4bCS3op
+a2q3YyC0SwOUfGrBxYgyMsczGM/HDqPceOXHQOlOUPR3Kk4cGyM2PxuGiTGJef8
Y1skbQMgnfIT++GM3tQflMldLcLl33EWGuI0MYtHDgtlujDseKlF1NDDzGvWxul+
FCaCSTvpqHcdyeS/MBBl2mVb0T7ns+uH8NMNzeZ62vFEC4jnwunPb7wKgS4LGq48
SzNy9L4qUJiGNEylyWAneVoIymASbyVP3tjgMWHEt2jYyrnL4+cWAkjth284GSRJ
JFoS/A8Me89H8MObuiPhVxGR//AV75QCMn38/zv/kVBZVc54whx3V+CstIn3phGz
AHBrtzooce869vi8vi6nkeanywcgaRCuVUdEmJ7fgPmUNME6ZruXNW9YGywIjh+F
reu6NEMP0tpIqZg0uMcLdpDVbj0ZK5nIrfYBtSdcZM2g5YB/Znm6YsQTLs2qlNdA
74adlF55aUGBm2Hp9QTIb7qDYAdOGeiuTe2ER0Oloe/Kvc7WzfIANq61RGs9uBOM
vSBR7wXB9JfI8UwHaFk5KGtKYmCXUtMmtvoeNgeM2+J9UPc6UFRU1anIMAXg1Bib
QF46MqzTEVYrX/D0xCTtBpPv0SjYWkhIRToue7nV0I+3Z3LpVTkLd3sbw96ug23q
liFEAiGHAAi7M47Qy2cp4UU26qOMaoyYLgzUdyJUP4q9PgQpIu9ONRY4kDFffH6c
vq3U+i3Q2M9BOJaCIcgqvDsTlRgnaTcmKUbA2AqwGCsklDR7QRHwCXVqs/+UoEvT
WZoN0UZa64PHp9N99viYzjywWQBCXg1grgDVyXo4ZyFqYpoxY0WVp2Pl3lfLv2pS
eGCmMSbqGJ8sTG+fQo+P1wyDpaMJJOHIWtSGHvS2H3bR4ryYkB6ib32EkMKvOCEh
/S5gUJat2mn6nN3PsP7NCHtlm2XF6hNcv8eTq8V3auQX1qHaRcJF2fK2GlIp4yki
glt+aOA2FBvzSZKF6APryiPiaK4RNi2Dchf0UA0GY29UpfiYslqTuNeOBSiogUq5
VM6TgFypPjFeC55g/FDa1soFOZxH3aC01e1JzeqvoZRLWnFv+j1mqi0jJD93/GCT
pZXsfw8P6jimlpyIzbC/Kf1v6t66u5jsWBO4zzIzAbi6h7lJwqimn5Iqeq70RUI5
D7tWvSxOdF/9kuLkyKxiqtDacO7QeNELfPLNN5vabRWSWrNjlI4E/D1QFbgXG0Go
D7A870vrLCQhwI3G3DIyLCVsGBc2EgdlcC9Rit0iPwq4HQwQlEpIf0rYuqn9o2AG
CzZbXPw0/jPHaekO/4+ge+wahxLr9NWDFjDWcKIsCXsfIfhB9nKv1IZ5oxO0FH7P
uL6TDe6QIwQQ97pBJVllp0olrO6+RJfxBuwcFLxFOTtyeLy+b/L5UkMH1iCLGTe+
jiNaJl1ANsxcPWatOI8x5SsJsKkj5sgjkqG/OnRGFM4f+/yuJn7I6BVLQBC98ihX
HwEcVH8pNeHTFZkERgWh/AsuE7+P3DtqZFocDyirrl0FCfvwdIY0myqxdDA/gbxA
DBhSM9UZrrs6I8X0Q6P/0zEu8skRuLICtTSbODJcJLsRbsFCRE0KsfqBE45Byz2B
ACi2ktBKZonJs7+y0SfqoXSThMTVqR+EmsQjRJi+3o5hX8rERqvItISqDqwrVYnB
DGctlG2ZajzIvnHvtwueE2Gm6vCH8BwGVabMGxg3CRemuEkfpjg0tbHwjJAXLdGF
1iAlioTmlNENzl9aGUt8RQxjI5Ljp1R66DEK2IfTjZFHKC6peXWxekXViEdvX9Gg
Q46zmAODHXc3dhXB10FPIt0z8qqRTeooB9feSZnYYImXAj308R+mvZNmGOvyu16l
3pnwS5PERTRffeifY+ObeqNyF716/gbpHJuq17Zjdd5ozN67sl4pUCklJT7PpQcg
OaivH9cD+SW3KUl48NJf8Bxan6BdJBP9JaRZbQoYCFjJtpxuEpa/X84eiFKEUu1o
+7BWx8x+yKI5Zo36sjesU3Bi0HF75le9j5TTI4938Wxg0keUsySwEp0PHR24Puq7
SoNb6z3tmsMQxcsNZrt9HfQWatRHsy+aPlgrXdzwfptyO4kha6x9BJfb2lyL68Hv
3Y84CgZvkk7jH+UFLz1ceSEBO9ubOlt0oUsZTwk2EXlgMcBV9Ex92iSqHN69ecOA
1aD0OYkKeUMtp+Vvnt4L/lxj3MXUkUVU5qrDkK6h+OXKkFjo/thVGJvxDoUKs/2h
S1OKjX4eFr1zCpji0YbqwF4mm5YrW79Lf3J2KloKDSZ0MXYrd1VY9FM5iUOxErY+
amXNlwngeb7VS7jpeJGPBGolifsEpM1dE/qytL74hEFDx7/S/wxp6JM1L9cw1WB9
nYtp+PO/5EYn4O849AVTJ6U9j76xpAAgW4xLpCK1xdTCt7DS2gpvQA1VsnW/DgKU
zOBcKFzr/v3swhtfqum04OwWWMfKvz4MNcOwPqYO+BVYwvdTeiz08mwzK1BOaZwS
bAo/ESx8zpCghdcuq0Uvnm6warZWqxbzxj+RL8PokMJX2WnXcbzvBfcRUICTqlAA
ewhLDMlgAMxjUUP/GYF2W5asROc9hAYCAnm84Wt+a37nsMcAG7DENF8FFjnmtX96
OHkbiQ1007lh4zWXj2v3szadxCAi+XXbMCrewXg+7iqRqhJ4v8sZ4JJl6oDTrtgo
ynQCPH2rjGlMrnEO20mc3TfhkhatwQL59V3thOmd1cH2mzlFp8N3mxpXOP8/P1FO
N2jZFUGKwt/0thz0iJ63U4p0PTn2MwH6w7PgABU7q8wPyx31TKqDq/WAduBiyXuq
BcsrLswquqYKMj3NjiuY9SR0N+syPthaOKjwX/9ELTh51zaOLaOwhpln+KTtkPFk
QYrka1JFuia4BV2mZeY0n0+bvR/pI5jvaLQzBby8kLffQI4dfR4WilaEpAd+xKw9
1TK4RmK1YQHfJmuOmXq48vVMgBaEoBrGFedRu6VMUVK7kSr1QcuzyO/f1bC213XX
xWLJsgD+caOqObZZZi71OEtQWobiW30GQJwRi0GzQ/GCTX/21yiNOPnjv5mjcpd9
kcRqEZtPX97bPi0owuv6slGg63spAswLdQ38NlqP+E+X27paH+g6aFna2rENX5bS
uhYROJu/RqaX6PSeGm4eK5x0y35eEN64B2cVzcsXrXMC1qFG6UzSC72pttDWj9yC
C/HW/LCIJm/trDpoF9OgBGVOpFhjsFhCX9yM4atjkYO0YzhGC6l3VAAg80H9cUcN
Y+h6H5KHbqL2Z9TSqeHhplTT8l1aeWvAgVOnWp7i0MtJo3kft6/EpWJBv+/CaIXr
eK9qXTSlvm/v9jiQ2DO0ziSDRQC9KzOUuwfwvhbTUqR6K4HdM5tAyJm+jC3Q2kzY
yj9V+hAsAqdVOYLhGmsnnOMCpiEDCIjzcB45/QrS71nTKkua22eutz7Xkd9xYGWj
w/6T42352dSmL6NvcSh2NCkW6/5j3y43ILTWijYJ1E0KPxKM4YPS7/lBIi6U6Lqc
LKpnR7x28t1MBzszetMSjtdZjMFUvRfq/vyhghDqEGxXqfyimDJ2rIxm/q9aB5bR
ZbHjHlZW5H33f2kYv7f21GBAbm7vWBg260hpyj2/nX0HG9zbA1ommo4DPt5XFsGn
Xgh5+1bIYRs8KE16jfq+hQLWYLHus2yBlv4zKtHUinrtirofzd+fZRZan5HNutaV
CvUzz0l18s6tSswRN0Dzea/SAFBDmeSaCMheJJLluNMmLyFdOHlUfw+KKInRtkvn
FdoYaS43lw7+vvM40ozib9pjvLB2ZAED/9gN4coPxtsPGzAJJrx8vUtycW6F/+O8
u0d140bCL+bV1h+Ku54oDfPgYuE9wYT6/f6X+5tU6MNW9WRZlHt5qeps0ohytnay
Cdg+oIV5SWPZuFhQnssPyo2Jaa2kl3GPj63KZyFtxcwFGcQGcx35nOjPfaY3gcnd
GD66uHv5gS877LzpDlXdSW/+2DK0Tj/r4rNHHgPZpcD+IeSQNcIMOd+lRDI/jQLP
q5wLOk57no4dZG5KID2YZy0F9zZ9AfMZG79w7x7Yvt0eclwsj6KVp7gbjo74PqKk
1Lg66nuqVpCZk9hXA98JmKMSphlkS9QHP14YclG7wZAt1ZA3JkY3pcNnojsPV1Bl
BO6Hq6Xag3kIYc5Ww2SXHiS4RziqCwUi+oLQvv9QnK66QPc62a1TMViLa5zdc0Wx
w+RCWd+uCCSJH/oYKtlLDfUB4YfzqlFl43Hzu+S6gDj/y4pVAc6oBjayS+ZCrTgB
uWLOozkPPPsvp7GtViG5YQyLl3K6hFQgWC3oT3lPTQ5KU5z3G116X1TQVc2TDjHU
ncXH1QM1I8WpL6lx9sdbwALpeP1fKJBi0PlY2IeulrX+vZd3uLfiqlPcO01NOwsX
kFP5/hByNfBnVre7QY3drv/+Pm5ijz3sGh6diKed7wLETBdTTS2xhKHKTv3LnT7X
wZ+o3ItKq0/j2hCnx29D1IWrCj8tOg4k1HrTouJVn8+AjHydvBIUjDUrrkO9ycdZ
I6MN55Pu/0XWiXgTdywwvwEvi1gZQmcJb2PWnZQdmEXWDCNVDnae652CpVXtaw9S
V5uvhXo45FmYDFz6/cw00dSn6iPMIolc+MkgTEkBbLaImEVHFyyP9B5kENzIAA6d
GNBDWT5S41WLfDT61Czz0XHDKtetSg6/ijum3u/pI0vwsTrdq4cXc+I+YlriVvw1
1qYQsEqCWithYr3B7qjcwPPNnitcNmJ8yvN/jqH4wHMyFKtCFIHpiwSFlkEVYkNn
vuOTyulcGcJtiINA24TnnkfOZlQfH9IbLDtR/eHh85PNN1bt8C3T7jNIIvXuAWfo
1ym5SdEWYO+nYJlRQZcvkvZjiK+AxOvOV6eplNTyRM9HXUzDNbRMFD97OSpc0Tk6
wVcfV0ZYMquf9oVzZj9YHsTMsgIDGwmgBaqlcmDaS6yZ7/jnxj7seQ5rPP/bwqZp
nbvEUUVkS/ECrdJSaIHCenLPyF+aAV9DAeVxDCl0j5uRKz6xBXqhTR0xvmvhLFKM
Uq7tcaai4NCTVO3GMcOr4FRREJkyI4/yM2wrgvEvqJ9TQq31M5UZXBfRJd/M7CXa
7/iJJIJky7s8uZzkaA6d2gkljNZxbtyoGnCCW/2dDmdKEvTokd2ueWyefyBR0gHI
Lkv7/Agm40156ZyjWzsShsWu/KH9FaDRWFyCSOmvf8Z/EJCPNvsn0+F0dH/58Ws+
kejGrHriEcB0+Z7lc29pmUpXT24Bwkg9PGpl+K5f+WjMPosanqWl8SPZgiI7UIEY
sVGN+rtH/bKhpJxUIup7JQlGAx0oMFvl1aV8neZVWXsQ3C0qhQhh1aMS84QmJYo9
HhIlBUWRWesE4vghB32uLT+Ti6Q8JGqt+U80IP5kJi53DAqFe9dJmn+deLTkcUWj
smaTU0C2iG8mqsrkHXfPxHxYEiyZgY33lmC1QSRt5dwslk8Sd5L7bCLMhGFdHbuc
GvsvJPWWpAaUnGY7gZd284GZd54iRkeO1ZYQp1QTRW/cyBg4h3HSx4O9zKk4Avq8
HA3Ynr2/0jBFzsUu2z2g1KHrbOWpAod3kSZTpenl7GsSlbnlCPqCG/0vTgSjq899
XxmmUuuHf4T8KwwFDaZ7Fd7gUiZblLYv5tuu9Zh9+M8k1eGBEULPHqXH/hHF2RW7
4fsLpiT8QG2urMxz1Oo9I7Q/412p0iW+BceYGf/k7DKG9gf1f02y/I3QtxjvpkBS
J9uqQzxUwsGfvbtxnc3v4j6Stx28i1+m4tnzm2SXnqWRTrehAQ7tmgVvJrITCpUk
htCpG+vhroYNJwDjqBlFG71k0EZJL7Ys3Uq3H0k4UjXntrGzvcOV75nuPsh766/e
AWWSPm5SnQ+xVpaSJvx2kOwqRNyPn7JrAARweBERYk+tla518/Ao96oRShBr29St
z6tcJl0WXylBJuRzooSxdNTWFYERSqqHkJJJgswClX6PMmqQi0BNxnvH9s8koFYs
QhEb0FZInZQrXwmxYELBfKZYTWyf0L5IoGJ9F5yC1sxX+y2/dyl1zCBdELM6hNBn
DyRTPWEnP91ETLTLnG6pEL0RqivAO57foAvN99Tjmh4rSz1NJjP5ipHeMnI2fg1Y
SRr19uE/plPOCS2pD03Ikh2es3YlUzHoYh9NO9KERItJofiKGXKyKpt9sV6UWKQf
pEhKyGMCYPM2g7kP3KK74wr3TtDSjZBaMp9HGCg0rsuhJRKWyDygpRSvluIGCD8S
SlqmIdz6jt3i3w9zqNgkbV1MQWGhIEG10iW5sA0vIaIWDnYW5UNtxaOOlPXR9AJ2
Sb+TZpkTj0V58vhYf8oV5YcggJuSFIRvdQMxKgcyFGNkJNdSYnVdjJOjzUwfym3o
plmntPwwLYr6PzoZN5JXIPPjeK/RIrJHt8ws4H7x2gzYDw6Ddyyrxnu2wDUFHWRQ
rNOrJdlVDiry8hylKNS4cYmN/4cpPZZv4Ew5Rca550ltpWTeXtoIKL3S18803KLv
dOCEYms2EacE1m75+BitkapkCRATTqnrMTBH1wLglObXURJzWVE55A5Fs1KcWsWx
ZFPwqD2+62KatAmXU0BWyHzpLU2UXRfxWa2yYQmAA3VrsJYnAtbJKOB315bqAMyb
KRaTdw6xVENLnlBNwJLiMHP2HOAVhab3ZUV5Zw++dML9NCp7zlNFJiEbgDHKebip
zlJAnYSwSGEKPQTjxckes5kAX4tsF1ZKM8Ndb/FiV5tHb4Ksm6YoyZuy8rSwYdmd
49nHE1WaC5HnPMQSn1X9q+Gw0Q4Ze7snydY5QUhaLcKIYYAYk/YyyGZSeu+ll403
JAVvsh1xUvwsIQTqz7u0yBN6ZPbp/TZOqx2RBUaV02HvpBf++o7yqwgI9yEEy/vd
0n/sNfgfwxW+SzkE9OVrWD9B0uNzBhXogkYNtIb9m1nbI+1WZBSFWmc3UaceRjtE
V9f2A++UhpFy8wGRcOi/XGFNDKWRBqPqXmAD8ei1CRh7mordZvzBSR10IYIRHa1S
VUetvDdLreaYczEnLd4iR9XnhV/cCiZhADUx/aUCbB/IfCq0/PvR46/SrkPDxXHZ
i6qk1lIyWIbE+ifYby272vE6MFSBFluoq0tX1yX88zI0t6A0Mym0fXQItCV6WtfE
kiKyLmfopNFljwLIwtFLKYvVqxzczhAqVWHV4hNk2rswGiEjN7yLsMb9/Kihsj2T
rJF75DtDNAsIOo5dSgee3KGJkhX+tMx0vyZ1W5Pyy49PtLI6ALKUWF93byUvuqdz
Ueg5VkkgInWwohHfut4JEWMeMvrXOtMMAgUWqmwu4Nf0ENttc3B8gN83KQyd8Iq/
0JfpQHMNihjxvzHizM/95Cjx9a65N0iUdOLa8NtLPYGBIRJSvsi6/iT66lrUl/Na
w99DRIQuJnajAZzQTQs+EGsi93+Y0hg3bkxY4X/rm+HU4snwiTUTm6I5SqdX4vR4
A0mmy6BtNhXiKZZY++mGTarOU8RSiFW7JcibnrGzmjmQluxcRYLfjriFOt5qaiYz
+AfuFF3JhYj+MizlSOVIiLPt8ULr8LrO3RlrBDCBml4yTOoX1kqbdt7xNRFbQpDN
U5aX4BH7WUCg+ilBS4U7GDmIHgZRrYgYFhklAsH20KgZ+3nxi+snUz92czGugWAP
zpynr1hySVUFLs8pEOsuOMRpy5njgi3/kgUeqEAB0H71dCYAyKUskzNd8poGiB9i
MIMip9ASlJbFkQMMCCEuNByURN2soQkjHHdIl0nCku/FFXYNPMIfkeY1Uo2Yfwv8
wrF66tHZassjPHmBRBoeJsMrDvCFWqmUZm3yhav/OvcE3j5b3IzDrkTF1M3SEw0C
H50L4j0Jpo7YcSQMlkwE6sSETogkR0tO82NNLv7dXA3WFIBYSP68utVycZudjKMm
FSJGC6W68G+vYmeFfk9U0HHLml1kWSkj+YPkT3IrXmKx9dQj5p2QoY8aJgMNEzI3
6p0kZt7waKNjY+4j6PBnAbc7U49/Nb5gaCxrP/6eepuzMKG4bAMjMMy4uG7Dm6sW
xQAAfA4oc3qyRyRzL8Wz0nZTJqgrM77iV2J95LZ28VuTnioo15qAlVRKnzXzIOqj
KAHWHyXvS4iBLWfG0Mjg69vdE0k+SivAgbS79fUywiyQUpm97TCSRbVVE+O6oe/r
jEkdcridZSGeKZkqdbqGd30QQ+iF/akX27T9S+pHL6+5O3g4zkDsoYU4mJTWGltO
VPyFiLAbQYHnYHTWZPztwMSfa6mnoTaFRs1yYrdy/iumEgOhpN7pobfC72gBvPiX
srH8HAED7J/5wtTQNi1xDNyUyhAUUZ70eYuvKy8QKDCfWT/qKTy4dnCodHGdqY5c
+QU24GL0bmktB88hiKxYcxoIhqHW90EgdXapRorvBYk8EIMJUAS8t/TgJjl53wNO
44cndkfoGclSJl8Ff0uAPObvUavxgOlhgQkvcWmFFgcvx/Nfm8o0/h2qvk0wJ0lX
29kZmt2RJ7t94QwI/LDKDgSF1MIUt/xt1kn6duSOwbzJr5otICEeABEZi0LO8Q1G
9QkRmTSWXK8TSRlyDN/PENbPMuIosaUJhA9HmHHX5WUQicZYHQzeuTBtWxalZcU8
2St81ff2keBVlZKXkdvk/yszVSSu94qH+DE0heBpy3fFstwT55zzU6lrqGwtaiwo
R3ftBbewM9dC37JWeF3xNHZNbqlXZxy8Gn5zK+LuRcVPiic/nLhYQZp7kzNaLnt/
n5dQIMmzdXUVlGx5yRlP3gJw8RYJVlebHhKWDKvPyTuxpDjgSnwM8+zYn+oDwzze
RjDxLkPO2oRGRdoBd2ubaKr71bnCd3IdcJ6Wn1SD0wMhOtL/i2NwlzhWocbXIVa0
jGHNzon6+/pzB0LDIDkWLM1QNBqkDEmGqAt2Vkwz0UIh8VZ3q7F+GtrTKT1rfKXP
JgwHJsP9tMmjT5yiZ30v0f65XtLMHcwxug0la228IESHLt1lTpPEnCwb7dyG3HOj
4Jv3OUPETWPK9QCQD9G3bZsIguLPqdB7j8cdxri68FlH2oz+f9hRUmm90liN6nOw
B8oXY48mXGuUEsZHaBH08TrGJ5LFp1C0jzsOLVeXrgd568MyS9aLTWK6r2r90iIe
ugpYOXbT1BkwtP8Jj/3GG1aJUF8uA2BxCqbQ2V/eeT3a5sm5DJAI3D1rXnqf2M5Y
YrU/6fSn6f8aLpry8KgL9Pe77T4gPAhmxSliCYzPeSqrPEos+sYOkiObNMy0hY5G
c8WU606SNsllSqH2R++GOgvfHw/GZIoku/oIOXEExeFvJlgGPD02bJqS+J8Ad2OS
6ZQEZwg3wK23yUfmR7cIaOGewCZUrIwpauJt9avRwb+/eqmdMDqGBVeq4trPrsaT
PxMpnxs48TRlUp7pR74GTxyMGmiF89g5Q+VJEmU8I41GNSCM3GcjWRvKn6UikhvS
+oXOvWBNnbgTOsSm/gzlaT8NCa5iwOg8DUoJP78uDZm4lPgWL9cx8QsPcmq9JCxW
BI07+9ZgvI4shuEqEwObidVpEt8ZFFSXtqq0mNH9fksdIokcCYgKYy3pf7VOugWf
mHCZ8Cng+0Fsqxqh2Q1hgvh4pBpM4bnW20s7z3+6EIyS9rqJgPaCWa59/W1HMKq7
kLkLtUPpO8b/25TPwnzIwU/x2XsgQmM337TVeV0qLHiBeOu8CFWav9/5L61vPrXK
XZnH+BZBDlSoEAiQgmBiioXF0CVeRXL1iQO5FeTLgcKLUudFRs34Wfvc+IUSjmZa
iQI5Nc/nGJw3trXFlxPJ5tYBggAO15OYj4i+6VFmI62iZs1lzcHJjbg56UScarv9
7OgZQhR0u9LSMahWx0u/Krq0bM3gx8Msl0MDt8dtM8QHf2p+n1AGqV7ONTMar3qK
ekNwlBktvpdbwDMsZMJG2o3Syh/6r/6lO+Ykq7mSrYRKjB70x6UrkiTAxXVBP4v/
hD3xj0eetX6NNMFtCBgEq9svxBhfX/aEQthS/XGs1Q9mAanE2AfSJHjqwLcK3pnc
ojT53KbL74VYve5cZNRdlrXS7aCS64QRncxqHHmVhV+QlkGPT+5Ab2JfhmHXHLeC
6EpYZrEDyzK25ks2HsyQMwwQug5y0qRMpjUmGrRv2mCx2B1YyQEC6lyLa1ida9H4
mIpx+WKjyg9d9TlnH+H9EkY+kC39V8ADyzM03LgCnLjwDPmLDGINcqXbsMPu2G2x
JaEkIXwW1PUghwkQ113WNV/iUXYxsz8sgCdyj5AZdqb3OCH4actN3GMpWbxiaont
Jb1wMXrpq7/F1Ov3I/OXFuBFHab83HZjvjSbtY+TOTCZaWQ56qK0EAbgu8aDEEFY
fgyyKbC/+5APMYhSCXJn3KhtpL9CUAcwAPNqholoihmuLjBpl5QKfMg26/7Gdsoj
088GtijpwZqT+m/b3VAUwtRMZ9kZSVM3IAijLklRb7kCl/Gggv24Z4SRdJycR2A9
EvZs0uvUHqAYE6TWebPVgA/vvEXprz+WqVGK/yWA7gk4j73zSxA6sJ7LzUtargrW
ItU8w5AdBy6Zh5KcGiC8Lhqsu3kY8pJ7fYvKdM/UyZxiWOWYJrhL2okU5HWxplqz
XZcukK5/wSn32TUI952iOElKLd7761DrlBDPmun5gr276CwczWLFCCn95S06yKm6
+ZbF32E/9OCi0Q82IzA+v1qeiC/ZCgMev3TIfaaXUjS41zJqSgUKLAWVNdksWjyT
EfCeo345oX75gh88yl0SCdp4/YHEYJlcsFat2XD8igK3RYhWUa6eCD1+bUb6SKII
DeRISd4hGlmQHmWVm0rFoPeLvSGOpcIKWt5u7iUuSC2wFLIMvWlXqffKTvxvx+cd
NgSa1n6kNFmYWOKLlmo1DZa9UWcrLsnkOthRCX9R7b56k8Q5/VZpbE1LxOCMkyAM
GJT4ErNi+9OOXqXFJ2pn57BSlke4DCK/V7c179wArMYrMvx4VUg330wmRgAoyY2N
PSWx4MQOtZVNpMwn57iD4twj6P5YSDuKXYdbaEHiN+mm/vMU4/cel0XT9uPpcCMI
nu5fy8Mtr8vkdGaxYFhFFBWKFukI6f3FlOXgxLXn/T/wsGE9SLdwx6Sw+zmifNEA
tW2Zws35hQqbJcC12MJ81U+foQPB+SXIoXyYLw7nketwsoo/BgW/Lsbfw2bmzxIJ
8GPkdOuYWl8wU9LgY9LaP4YLLG8SgPxrFFKHg3v8OL979a5+AnqSjhPmILVLmxXq
5HnG+L/B2jKqtmt1J1ZJgcXXm8QBOfNv0a+bXD11jdcLq0wevVsBYo61HAXQPBwi
WQPHhx4uMT90m6SJWymaj5Eoino6FYsYXYkqEA4ePX9PH/z9cfxGJl1DCpIhHRSN
nLi9IBO21oPR2iiIKenHFYCj4r3gSvUaaiLxElbrRi1iRgvQY9g+7ka5aSoR1tHf
YNgtG00KZS1xhl2ucmdRNbrcBSP0vxrmU+3FoO3TSFovIDYMrEFSKzUVs8EisVKd
pEWqyTgBpV4RqjAGWeYseFTW5nZ9XBukT2JlzW8XqM1Pa0gUI+WB9UCew2pojlR1
s5UPJ/pmLtJBJK/HLXO7+WuzlMlEdUu5JJ8X/+ybyR51qC2NFgjtLtqGTBfC9lKI
ooOqSkINJt5FJwfUiKRShdD7B69IMR9UTcM9LktSlko9fwdNR7yUey8DoJ3qNlDq
tPykRG+u15tzvvRTqcFs5mnY4k6ekio6MDtIAMKPwkp2pL4g13K4qIRv+4YfvKlW
a0Tbwa4z7YvO/+i+kKw7A86pjSXrA8OMfcEM3ujkJElBq5K8CqrXq8fXVAW/+A0C
ZAMh3taH1jI8NqkzmRKM/kPDnaD1/umNwCQZCjQhbOpoPGssh75UEY7itpZGO/6J
tPfqEDmC8SXSDB8iU/vthUAQSpN5vwpnkNijYMvUN6+8jEptAq+7gck4GcwbajFk
jTarsBa41eW2yo0gxuDt61uBnxfa7+qJdRbQtSV//APmWOKkFYiyl1yK/WVUITnJ
/Ihw0ztpz0L4bUfF4CEvE8B6TSK96KCIPEjnNV70nNuTp7y90iyyrwyqGx1VNpmI
hdMHmrLJs82RdTEE1x9a5ZQbr2QOrskgyPN5GV4iLHBL6JgC/0TbbUDnKiz7R+jR
Mkvx/NYpIUNGU9EAmpXu6/JQTtH6SVzo2pG6Cg4cmEVeOvschuwOcxJZE5JfcQ+y
Abvrczp4oGAy28T3lcwtq2wIJOlfAtey6rJI0CNWHXy+Jmnszpm3VeVkscUMwqAY
Hnl5qPgD9lR7RTQo2yJSlGyLCu2slUwLzVZRB/88yUZKrAK8AE3Axuid/5prC/DM
Ihbo2mtD7aNRm6Hy40zKTYdmdV4u7MFT4l2t44amISVk+OA0RyQCss3RSwFn4Ygo
waOlkaDHoZjalYECwlLVPir6AodYgambcW0Y5Lcls3BDJHGw5OMdBFbJOXW8VIBA
6hWVc9f4+pALsX5OReAPXTRRvZ5SGIpmXmveL/1cg1uM75kbAMx0lYjHZiDbz60s
0BMmWSrKIw+18oXVZvGrkvLPSaYk1yOhA4nsBLhDOPiqbmK84wqrYi7xZTWpAuEC
tO909sK229LP71O0BxIAJx7BUbd/njnryoDy/OPtCr2Dximvg0Dicvv8M7QCHzrF
L2EyBKjZmmZrAEoX9PFHVyc4iPtSu09+IZ5wpaZn6XPZ28nLftuYSNASWyBVwS2Q
bVdBUU2KrHfm+fZ/E7p/DNxZQP1wKUXwS2IzmdAyXG2TCtOSjJsSKk/wYwXtB8KJ
L7UrVcmOp1HCfwq3bbJeQ9UfW5FDan0hE3pbQPQRyjqPbdsLn/VId52uxPupRTzp
8PLuS9492GVjBWffzIRVpdIC0opcqCIf9BKAxc3ZJrElApRsPlXacSnykTHBqc7g
NOMYeYeOmgN0zOy7cbJVtpB95uPtovYSZcWIIrG5pUU/ifh1+BZKFrsmN7bftquY
nJ3ZnoBqZPgqSD6DeJKab8zZoGEMkuW4GG4VUkCZ8+to4gYOBlHgsATTnDygHKOd
tceukfvsadkFjOvi6UETjigLqeFTOhVf7ZJv1fxYsOeXe/ihu5wWMQvLXqjJ7O70
jXe/0fwFLqw6Uhp9/DgGiQRzUte5yh3n5VD9NrbjUIpqZ1ytGttxHXXP/Q8SATx/
g4xrD8L0c4cXtcuNYGWHwgSPK4hWh1mHRE3v0dz79z8+rertvDXQgGEUOVgO5YLG
9cVwJ7WEjp8I8cVeMpDchSNXRqnudFSWuYODxUnsCYeghdfCo3ZTvr6YfwBHHYzX
wNxu3SrDN0nLpXoN0hmG3GGy4sAUxqhfk3MGQKdrOtUHKnB5KQjbvlNrGOu2TB6R
0UF132BV5zcqDotKjY3dw4MTFMkInHWFORQ8njDvtIsbAVlj8C3EQOGVkiu0d0rN
+12aXjWSbtGgIGwZHu1nWq40IyeF0aNyr8cN+gyZa8qdk5CXzwn8vcltHNkoe11d
ZTWbwfd4spo807btfS2CLrllgO142ItbPc80EciugP6a/TT8QQdFMF8OQ76g+cAb
nh02H9pf02X1OXdKdhbV/mtzXprq2SMzChbLhThj/hSWUjGfftVhNTdPBXqqMQ3K
hMfdMRaZkztLxNnv/LGM17QipAi2PVaLyzUxZg1nDSQgIH0kna/ODRV6v94STIhJ
Cq2p1H9ymrkiK+Cc3z1zBPtFUx+iGkAwTJbseanYqGUCASicdgRzS4Zr2HHyVDpt
PpXVYSDXXgtm0cdaYqCWoMvzrOe01SYPcv19KRH2gycQbGxR3OMHCU3Zvg6Th+dU
hzrbrjS6wPflYgXrr4LtbgVdBfUfNqwQhCy3MtkHxsuTjwKLn0LB9bX5uQOJPh28
1Xu8B/rcKM+PonPth0e9I7DP/Nq+iUh6ukqDl08SlorQpLmC21Z/xyjQiz7lpeLI
8HnjAx2AGEs+DtWwbcJgLQfjXh+E9WctoynXQSFu44franloNKF4fg9+m4kK9JgG
+yjS8wn3i49lfiJosqznNuPIkxd29iYhl96vFHadStvoFL9MMUKSNJBo6vEVkHPJ
ZM1YZdJCKirD7MxYZHqQIlCjqOKgwHr8OPM3hxZZAKi+e46oM3g7OpI7JnqbbVXv
9WwBL+r76nnSWV38mYH4UBlVSNfhbU556GkFzLz+68CtD/J9Lv/lt8zbi9UtstYB
8M7ABfMnB2rzbFCvhlFILiVM1PYFteX2ELRQ5+9MoKNkqJSeqCMwxg3CBYQdxijP
oNVT4ifwwviDGU2hwzmjboSgZ4RMw809dbEAV40AzssG+MQjjaN4FAruKd31n+A2
P95ZmqCSTq+di1Nsn2d7e6KsNBNywYcZ2GW7qBAOeTTTcCwdTSIvnTG14Y0yot71
pj1T3kmI8UYpaDK5N5DFUs/uhgJr84UI9kM9AJKR3bYqkLPFqLgtWGuX5L/FmJ42
Z0tzVyfebk++SbdInX6Cbh8M4F5iefumXeGWQXDtPt8Sqrlh86JrXFMd2qLDQAMT
AZ53cCc/Uzw4VUo06j/FVz4krBM/AaNkJVrb7OLrZjmGAXjK0hpDS0T6y6DLyS/E
urKxnIv+tjx7ZqoBik+/uwZrhDuK77Hg/SVdsS9ISH67GVeWC1OK75LielyKM3AY
IwXaEIAikGnW0sq6Kl6/IGmTZF1qi9hPUeYlf4OgYXm5NdmrQfU/NzDgH6hyqOB1
b519/QCV6/w9yADQwqaM4crld017ci4MT9gzK1VhYAZlNIBVdSwDs16hoJUbk+0Y
s8/wE6dvy3jkdIvvvQk1S2l1Xa6LsrLfm45zD/VUL2GnLYrY8zIQQJEdlvPo6oV1
Wci2oYc8+3UxkLSPmX2fkTl+gs0wMWeUPBp7sWkWgU5pV8k3n6OP0mzjgE1d7kJ9
MLe81A9WmBQIHqM8pq53Oi4vo6Mq8L51RM9LsfF9Bq8RFnVzA6Mz+zwNipQnN32d
BPiNVto+TGew+78QlD0IOV+PJ6E8H5cf2z4xR3pU4GDVfcAaBJVRp0jEhwzLr1+C
jvRRX7djL2POHTT2rkCN51T7/KaBSdh6c9AJQvL4jywmyf4IhEy2ymWcnApgOFnp
0Cbw2AU5VS0WEAtu/j2S6rn4HCG8wY3j2RtrUG2nG1PsrY+C3IrWcPHLSd3oIQgL
X+DWBmUxYao4RhlMCUCJKER8lOUXcoeNXXQVpj5739n9oP3oc/pUzbo+87dmRB8x
DB7jiRuwQ7x7Xu7TNqKT5f0fNemkqAt9aIXi9Vc3fnyJiRb5is0LXc6Q1Rcwmgya
h42fhCzOURaAzB/2CJ32GjBzegX9CF5w1i4DE1Wy1p6l+yohSZIZwLJ6fFWSUzgK
V1N3l+hQnUzJsPXzpWiSsFIHm+LioRHarTTNkr9mMTRRycDA7152zPK71ze/C9yD
WKoy34BA6TilCfqVREh0xskSSxtcScj7a+nE8yrPw52FHmBa4obZs9x7ZvN2aIhg
U1eij1wmozfc+iBqNMD5ssdBAq6w1CuH09gNQiHqZWyAEopoQGyAKe2+DKZ0XojG
revXKd6xyFCda0TDLlHIBMopDvqKCHWqzzr67kgE6CQ7XTGLgWTo83KaofvZWhua
BTN/FxdgnQzSBefLqzYYap92dA9st4ukkc/wtheO2KnQcCuRRvhI/gHIEmJr6Xgb
/FsoE2oiub+5euZvxyYNPTML8XTXXvBjr80JuOxGETXMfY65rjzZQwIfx0a2JFUM
UpXUR8QTIaKu6F2FtjTk+2MvGKnNylMlPAw3tPIwNQXeg3bTn8oN8flUIhy3SnSi
64EiTQomx6aiUViP9fvfz9Z5WGdKzDSvwFcCZ0k7cNqmWOQTb2W0j8/szQHuyhUS
K1bd9vwlColpVrn77MZYO+ATzzbznpoKGb4DwG0Jl3r5migS4nJ6BPbyBq8Z6oil
p+TtbI3yFMYmanHKevzQen27JWI9P8ZvV0EowW74dRwb9gJbGSYK9xe/aaxxH8xl
IRSHbAqNQeWtECG3Wf8cxJU3yK1NmnAVztzwvB8xY6gEawol9nfHvRQDuDvJFdrJ
MGNHygueaJCnXO9F5NA4V/CwS968uzejVql0ne33WAqIPShEiGWvys8yL7ntl1UI
kGqXuir8GYZiybhRk5K8Wqlt3P9+9e1Si5Tn94RR3+oedJAJzz8BipuRnHVhKgM8
08CTng87H+kKoJ51l+Oslc3T5/yfyREn1bv64scvVNdBev3uhOcr0kC06d5KO1t4
3P+12Ud7xdYfG7gKvUIfURR482gTKROlusAN8vN7Jdzt7sLYxv3ot6yanVTN1yoo
jFJrMeh4+3Z63GjeX1yMdgZ6hiH209IT8cTpdRO+FMhKz9SxXwBo29xpn4xWuOYP
DfdeBr1D7oJWdUt/N8LF9iJBX/6Me7Z/E+MpnFSp4woIcgHgaAOY1ntGhCmWmwZJ
D2zrR1gIGHpSE6yyn1tKXRAGuP49xhHTdG9HqM44oCMXXTnHOYB3XZIMfBzvH4/I
OyTq8c095sOhxlPHHssS5/KvFP9EyCi6X9d9BC5raP3yswb4Em4iq4n0xh4isHNi
1A4Ka4ZyiIqFAA2i4TXz7a9+spH7ArtICaqE3ZcCvitNIzwyaXgVC8fWcA4CN/7M
hLtRQD4yaZW6saYyXuYTouNrT4TG+/oQGWzknAh2hrCRCyS28f2wl18piW+HJOmD
9INRn5AyNF05tpO5Ty4CxRu1/pXmCq+M+BH0eBi3Ei2D9mUTOtWruRPJSANh3gZV
AWQnc3X6rZQec+Y7Ew9XxJEMSVPBmEFxO6OOAr/k6+qGZvf5U9hAO9owFSrGN0CY
y3rbop0Uf7kUqhhqYcJ60SDKjzuwtjCSYD8SXkMa0uGHRdNio+X+jca5jo5DzXW5
Tfhbmw9aGlF1GBPsRh1tNW2yBsEnw7Mon1E1L5GCC7ozSxrN8AOEradYNVQlJRg1
T31X1Sc82nQ+64N4wYs6nKyWLdn1j5mNMzhX/q0SrmdFiYciOIBZSEC1jQukuuWX
oXF/CNjfZT/56/NH60dnl/EHbAKTwxeNfsxqwzss4hHVDwQSu5ghMWnryYacB1tC
gQwNt6C5PeKGxG6JERQ32fCLQcV7f7pinzGMsR5Ng+/JdEP/vnL0bpA13lSu4ag6
Kfw1uIQWLs3RaVy9Kwz63sGqteebo2n6ZILeFGTG0zhLmQwIM6Ni0RGMl46+vVGq
vtTtLjJKASCPkd8tG/4CHEUdUc11osvy+l/yC6Qog75JPS6yrt2V9Q7t9oYmNCwD
yEGDKK14YNemrI6bnafqp2kOJvCBl9DYrGOmT0BcaL4wnmuFJpxd6Pzod4N0RJVJ
6ZgAEObe2ROJBqjh0f27n47evpcd+2QeFxPKo97XCLcG53pxepEWmsXg3wuWgtp1
7TilMwL5JyRNwD+hvdc0NnVYZxpnM4zFLdlv33vZfi9ZGB7AjcfzUaRTEQPWIHmU
c9gT7QG4TVAQlzCs95HbYwdFqYO7GkLiuMctdB5z6vOvO4hN781fxl4Cnnv22yN1
uq2W0uE22L7pDrZk1yS3y2wu6Kn7mc9F3T2pnxYk2khheT8P8oJral6bLEnszDJT
krL5kznoqd/DuOkVvpxZ5OmLp7wkg6xmsOgt7d/YGhWBfNFEl96qq1Q8+Df+BrGU
p6lKlUYoEh583ssp/ZgLyjbac0VT8NzkGi9YTn37+irEbLEYyxF4wDQQrDK7u/mg
fU36AACq3RCiQoMQWceiVFcSntDcRV2LGd42HNdeQT6kL7vWeoCNfupICOJTweqA
7ePBVOdtV2lIpEsXemLD+vTulcyTwdipYxjhpHYJtboWXB5tBXPyG/349+TQU0eX
PBH5uaqVioNUQA6Jgbj2hsB360T7u4UaHKSGc2lxgTn6aTdngpy4sNnyPV2+9uYW
L+D1tCvPAkuAk6DaBD+1xK3dbJqJ2ZkXGHQjSMNTI4nUzeoKRoqr4G4MtHgpEC+I
xZtSOBTkE985Pfbg7d+njHBSRy8SGSQnvrxoNfpDHZuTWk5QWrMz0uuu4AjA8z4z
a0S/sBXve8tGaCTckyv80m744m8jgQUwZ/rImnO1l+6IWSPbo6xIvfkx7hxw+mhK
lmwSPFCeEUntSGwzSM+bTcywbaaz5fH8OOYrYUEbKWonxa31WQtaMZ1WqV84VUtp
LTPFXaRRK/6M/r+baalBkgrZLW9JoZzXGuZt9OQ7iiyzuy+1ycOlp4UXEVLKAdNd
CjKuKSGi0trmAh6hpY4QZy0yrqM05/QNPaJPH2kYnu67QruD5sKWbWzcXEIWd3TQ
rnP+eKemzqfnIzPd+bqF71BvFUNk7fXx+OsGO8PPM2qGJ8BKRvqVb8q04OQ4VW75
KP+0dnozZWaxkNjkZfHvG8ltSEbZxOlRf/JAX+QxUeUwPkJjpgK9PLbiskdx7w0U
O1lZL0GXpd+ZOt95sDfcNmi6O8Ocjen9NKPWQrddCy4HrWDupwtYfzyR3xsrjDfb
snsokmMXuCnSx1RjPDqz3KU2q5I112VNvgRn/L1KOSE05aYFYo5JSK26Nfm/wfPk
SkcALV7bE1zG68gnePB3Rwz2s1Zdy4QfdlYC2+UDMIEHvdYmRKOG3aEsCLeieuLV
RjiYVz9NOvotjUIbdYkoBzPyWKEYYn8IAhGVhD4LcGPDIfP74lteLMwWcULNxfra
wewX0ciy20lRDbBB+cV7Gmqd6MS9V7WR0VMsxL/0vQ4a96ie1WcP0TsVeOGZRVj/
NHQpLicGjxygVUrr9ln65JfyonKK9ylWVGOIAX9W/Svg1c2HH3hl0MaCQ3MvOUmc
Uhv5SmEHpBLfLGzNXXEeK8Uuv7D0SHwMnw5VK4ghDIJaKij6VQEQ3CVZcEzFo3bz
bHMq3bfhfFnBZ0OjgHoN/AtvZHEuEylGVmPGdgl2XxpyfXHMWjcuxRzToPLzSwV6
6DbNv8F4SePy1HDutXc5Y/RZtBgUVPkFm5k/onFN0oUGGZznqSwtRvFyogHvXu23
PlCDXJxLXQuHVUkISzqqshj/YGK3TEdS+H7pF9uqyF+KT5TgStMG56oKbKhxkZXI
H5bA4QBoten/VeeZX/tPfj644OS24fyyjktDKzGy4P9V1MkhoNz4dXilIALe7Ju1
0rNHLOZQLuRS0jk1dq+CxPXGVBUtY81zcbxLRKEGZsu2EUmLP6e01bFRQ1axBuIj
AnkA2N92PJoQnuYsKMG1MikG8qrWGJTBa8A+HiWuLEFJohH1BQxJaUV/NayitLG9
Uh99kVbSNrh2uSuxwn/GPf2bz9vs4E8VT0hMXCGhBPG33awPPu5U02OH3tKaSzPp
oA1GhFE7JrYJK5butxsj1iCyHufNeoQiqqTAnXK/VYtgkvSkg0mp/SiCJcYtlCTu
biS1GhsCgXzLlyz6PGn5GvYMSj9FmfJzAFDP1rvQ/9GGv+sLdCFzy026z3wwOdEs
DqSgLKVQ2vdaKZCdbJOYICCFsHsTiE8eGMnu7rqTEWjynsisEpwK4XsGihQNnR8g
knqRS8QWx7XjlIGSJnIWTUeoddMo1a6ab2xAPTm8LmD9OP7gTGqZLLHgdCDXhTIh
SQYEGLef4qe/sOuQ+FnD/BQ23vfIqJMq/KTq1E6c1DBZ6uyfxiQPc4tS6r+QGKWK
gSO29OmxTwl+JXvsw3Qa0wInMiBCUmotL6tKTrjfRCV9QO5Gy4Dc/Ppl4wnt84nL
Pa/FjYmqlAypPnS2kMvdTAOm640KzAf6T8Tpj7HdnYr9Tvn7D90QuB7aBzBhxMxs
Mv6ZVXsOO3uwZCshg1pgMlSaIwVYwpOUMPFMn5jLPxZmbub2H5ofNOl+REfXIl1C
QXwf6VjilxgrJTXIZptzoG36EwlwAaYO5TC2GlEKLYmX+/pZA1ZBPiQaHc9hy7gE
pj9wpYH2egkkoFRi2n6exzwpN1YtaKN27z5ei44k31XM3mDB8np36W3E4zv0RUyd
ravYqq3zVFJ7G/rA/e0//tsaRU5jKMdpVbOCLtJRvK0nScSzNPV29hoMxLdFHiaW
zTq1bOSeFyRJr3Qr4TGCAyVhUtrMO+cmKGUiuIRYhyHpbhdLo+NGzlfcEJm+74r/
BXXiWwLEJCHEUmmiUZ6viPAlyvQMgmMoHF2QGAVMVmxtiERIiM0Ald3TNQwmCKDs
Da6+CUPiSGpl8lhF5oyT/eMhrV+g/Gb29XXjzdHdw87NvtOR7ECQljJ5BbnX4cZz
qvPyIf0vljvpQjjq0idceVeVx9I87B9df4n0sY1+CsVttrobw3Enwx6tpCKvEVQZ
mNVcKKeqpuIEB5E/gJB4cZPmZxRbn7+yXpNcbUL43JNCuw8rQMNVo4vxxlTlTNbl
sdMZF45zvpjwDvubagFPfDoCgaHXY+so5wbrqgOXdlj6lz28riuDFMl5/73exFWE
q5qW7O94FVaH8Lq2NE2HbQ+S7eBoA17whzDRePRuAXlv72LCzpm9FoOaWqxuvx3c
t3qAIQTjJ2RmL9uqHku/azHi9p5EecVdG7O8aD8hAn8iSp5IJAdP+ftCFTUozGyH
EPE3/S9cJ+LZkfxnzcO059OP7oWEBZDipVWCImF2eLZXiArkEEwnjH092B/SuVT3
03lwjwWeNj0f/tKeqO9AdJENGdeYFCzR0dGha09rISXMpamwV+UZL6uVOkwbAGvR
q8CiEMaPUkIPC2H/m34FaafhHenViZ1Noi+Ap2UzxNsqpEyX0vXZkrRHhL1bI1wW
clgPLR8t/XCaSE6MJAUDM0xQAfwWSpyQtcON4h4viLmPg1Ff0596/3rSYyF4+Jpl
xIMRGk5WOvsTX/TCK8oFXMI8T+gThRdTAcovl21v6K1s/9bphC0/9XYM+vODu4xS
YLm/QrsRy+MYLwq2HbMv+P542F8Bt6RwJsSnpXS7H3RNmHxSY2Rm1+1PUm9E1VyU
4fdCQOakcnlpwfyKtr9Ksuw49sdDVj8tFS0bJutKr2e5kRq0LSwIW9vLrggVb+v6
JD859/y+dl8qe946bhz/TulJCWpeAcL+reLlM7mVyUEUJACmXVpvZRpi4ofDCSrk
hG2OIcjGAUPl9XpfTf6Ee5faQSLrvAQNPYvaYU2U5e1IiA6m1DlAK2OoND2yyJtt
6aRbrxFmyZN4R+mmX4EViPySOFrSgw7SP5rxisHOScFKUB4VEhje721YTu0aG2nf
HFbuuJUNX16MPdVnvBDg9bxgE9Y7wn9eH+Za5yd4gs7IHQUqFNwFZmP97APUMdAT
Hvd9VuQ/FEzgBcKV8PPb/0QgGGzPGoZcz504rRBtiVKEJObSjkU2CVa63UtliK2o
Gw0SqsC22R0mvOrfdP47/wn7pGUw/v8DhjNnJnhcmKefTLvtCJfWRvpVvZefjiUw
WSGY7+j86ORAQ1TVr546OMmaTlGh756rY6rcZsaxtQqtd0QE4vVxHWdcv7KcysnW
QZc0w8dDbcqNR11qmcpFLaWoq0MA2qGYPMJXAJdoQrWEnd4sh75OIVHRooHtZppk
2KnISB49X2Rr60VOWE9ggOcwKJXijdXZksR0eCEUyeQY1V0Jt4KO/MT/syeF+0Cg
WX/zMWQuv52dLdBuCneRxmmOO8VeEfGnXVEABZX6FNAXBgo/YltrJRJtQrBQ0rVC
EbhsMuOHtiS+7M1fbPyjZB0AqawARuRgVK1hoLCa2lCuu+lZ5j6YRkB3SwX14YT/
p7uVFQMxz1I7FVk9NRbJ+uJCvW59BPgKFltS0vaUbck/gvEg4+UfR17O6mMRX0MT
Khcoyv87mgRbLUpgYEfZ2U52KmmSQ6dRlohZBmZWZ0NEOJ5Bn4/P2Q3hmmclJecC
aMPl+FdkU5ex3S8WuGeeG7PuZKm5S9KBH1BKYf1eySx+Siea0nxgBuY0PkoyeHtV
nQD/o6PlAo4OAgvcJT8FRnBku08WpiuadXVFWGc2NATQzKdYYGx0XTQOutrH1N+I
F3c5wK+6+cXfXQAI1QQlbkL+Q8nJygVobR+3MtE+eoU6RlIsAgqTKGFj72uzZU/M
gr1o/o+YtgwkO61ICKNORIvV/5isXJd+Ezspe2HaIz/VvEv0krAcTHjVPBZ/v5IB
hltsf8A/eU/YOe3Y+zz1BM1xwT0xK+zI5sLb0oLinhF+Pz9dmpDnj2OIGW2FdHox
1thPAbTrfJQsy/+oyTRbC1xYdX6hajKk/y6PG8QtQ0NLBMc1F08AJnWTOQodGRSp
WvHGgSx6BH6axltIHzH4Hoc5g5EradTiNc9q9pTwEkjlnKcFdc9fJ3s1dMENXCwH
CKUioqUVRnFP6LJQidxEhN7hoRkT7yta36MArGD5Hkc5GnE9orE2TkT7YW8OO3jO
yia6aJVWOBHL1mRjEd3nd6pzM8RMnQ2y5QcdoLQSmEnRgcDG5fpDAn1X40urOSXP
82MxuWC5/gTKchf7MJw02VGxAwrqqRYBquzkE0jeWqAATzjZjN0m/2BELyEehFi9
UTns4+TjBSROOCQFrrGZQTG02GYIhpW/JX1PtuXLw1Kd7GdK2AeIa5WeqHArRHzf
et9YTPNNwKevQRcF964mFxJslRIr6vldYuoa3q9N+4w6b2dyJYhRDhkCM4SBmw1T
YbMkWDpTP5ValfYRWoZEd/bGN9b1sqMN8mbIvCR6Zi9BSKtPBtnyf7K4IORAkNe2
QqQuGFbuOBJSK+24lbRia0DUXY6f0n/SXtm/hXbLV5JYyzmazT+gxdhDkaDp3Z3l
j83wPblW2o4ksveuvTWsY46yADFPfezBzR1GjFPYGskBNtKt0qNNhljDlSNSIosa
bd3AEyMu2NxVfTwKTMtyQVnzeTjX7LWXQG7WncsfjpQ5IIK8qQRIJ50rExVvqWr6
6+s5f0Aswhl8DT/xhvaT9Dn51Cx750HAfGNQ3XSW5BJsJS/m3wbI2/xZpNOCoJxL
ZRxM44hokhvly79iKBgOkqijTqbuRUtX2fWGmzdj/fQZhCpeA8qiV77PnJJzXUM8
+4uO9TltEMqhJlj+7X3PYI2gcayPkRIB9tgkw7+fsZb129VLQdbGvmWipZg/n/zh
JIVxueiKpyXWl9DJkIn0DyTnd5Fuvh7Z2kw/0a9cegmNYg/ZP9zIyfCY3/WT6CLA
ExIZgG5GDdNZhqrLdCVd7aashS6yorl0gYvl8RgdqVeoED9Wz4yucaY7NTeFh60v
tP6vFWdBk9bVr1Ax3Z5daybgHo73t9aQZWW+cp6nyIKP7OUiKSbtWNGG4UCQBOJx
SzpPEHXrWAw7e6IEwW4ypXZFuykquBMsf9XtQTDJtjbf/nfuEHON8idLwTpxpzAV
A/kKa2zs76W+QBCZhNcCCGLtnrUty+8zgc/wr4pbj1bunC5qmA+DbbPEOY32MBtl
5lnobyDLm8BUpNQf6ViMui96TNgA1wwLKigfxHk3QtsaqSsp0dF8LE0wIg7oPpOi
PSpSjPt+/2xZbdJj6eR32iAfGqCj+ms5mncZII1salqNOyopTwC14nAmiC9SdONp
hkkOE9oRAMol70pnUCJZ55w2RzUyBb/WZVAS3lC+8sEXDLqWLjyJB0OtB63ZHr8s
fTo7lFbPxDx9wz1S/Zzxw8eLZHhrOPEbkVaflc1awblzpHDGZeTfDo754yQikACB
422hdVS3bZIRwcpTBI0skBaUF66smLpMGdCTz1N3nZbu2KrgnKbwyYlckcSzFYgn
VJAAPr2oMsgf+rsXW5q59Tit0jjLGBYIBMwaRER4e/eGJbWS4qJcwaR6xrq0o+oN
xRYM/WscXNt0Y1Ota/jTmyr24au5nMLpiIz5RP3MnvfPwC4kxyzg4zWEOc5I1Xjy
gK+aLAkFbHvxZqm/mwAAiyhHrtulwV3Fk9pkSxvEgA9pSpoE3ee4QAj/67G4mK26
ZqWji1lW75amFHTusNHr6w6Te9dyOkY2Izxp+K6rI1DxA+vwu1qDhXf09oP3T/OG
rlciDt5nrGKeJatRSKHkRkt10yRzi1lGEkwbRjhIGubGLZAbn8pbM4Kn2eGlghmx
OUuxsHyhLlPf9p25kj+uTz30xz9jFkgagluNmvEgIspVE0rsXCG0FleSJVm+axbo
scsya+6LS1eFXEyxP20lP41qjzOvYfcnyTY6y6Zuq8y8SI0Pp5PR/8NCd1mBojGZ
w6a+5bPafLF1qwWnX14NUUo1lwAYVtGlp/q4w41ayuHnWK9hEALgb2nkR8sLF2U2
pKE3NOVQ2vQyo/fMaBgZGbSdshMiHW5eDPzEo9HlyF05VT1tmRABgrZW+tp0GZNO
wYT6FW/XQShD/B+XN9N4SltrVVPQEIxgpD4zQxQpd6Squ0gxvFar5TqPJrH64Ge5
i5WLrABPX9gG3V5emLa+K8BYeKIB01dwAKAlcpXOifpUUZBLZqcFAOpdYJmLxK7+
o2ZO+5TsYVUKO+iNBNupvj1ai/tpEh5I92zIZ0nepoqoQoJA1103byeA/zm+Nh2K
9FHWRI0QemLFB8gUfVtxkRS+ZjGAFR5786OD8MeVvPquf/5xapJGjeSb9GLlYUKO
Ml5jA9R3iDMGectr8kQfFQTjNvB5Xtk8MgduwVcsHIgMCcNHMSArDn0hjJRc9SzQ
eJxPMHYVJ+0G74AJ6gsuokv4mwnftmOBDuMbV0ZEjxHBA73a537EfUVEFUdO/L9G
VAAmx3gy0AbXYVMPFWXFwNbyMSVKNsr6bztvUoHS003/PPddN0crMxTPu2W9c1v+
wsqXkyXbG7o+F+kRRz03lpgNX/ux70RAXU4qcspgkTXQCNgl1J+KZGv0u8zSzpfs
KnG9Ra9Vi359nRQOC4jpgOyXgPrIG5fc3ym9ik3p8HGwE2W04R8pA4BOVwyOvD1l
aUZwFNfHo3nCZaglt9ojsnhBfdd3muhVFZgxbkMsepTH8xAibS9w51UWYTdP2o3R
YWv/uRdABpFSt5jmi6tGsB29lhMW1DpnAwdanR5HHo+SwgRbbJxEwcODbJ9PKHAA
OX24XZpjuFqx5ABqFcvU2AmXkKGORD1ioXQynaZcMtHzdCDqn9NzGjqfGMHAY5mk
CfUe3rUu0pjX6bVq4imk2Aj5lWCnP7RJCz5Fs29QpoF2AQ/FtZFopyFpLPmKQFUo
WK421meeOdWWMkt/YvLyFdVqbWTEoVErcx/0H9c+b9EmmMX9wbyfzQWUO3RlQq0/
lq69mP0/1escQHkbcnt2xAsVpHONojLflFmm/8ylC7NuPiCQneXG0l6F2C2Slx3X
wsp/ZIdRYhgHcop3B3gX8Sf6NHlcnzIthOEHfm7PJRCDx1EY+ROylQsmkdOUz3iR
rUOySxnjd9TR/GeDrrkyUJqSL+FntmTQLVTj5ZzxEMIVafs8rKCcY7uEpRwIXAT7
K8tTfQfeoFcDPIP2QDHbb2HyLwD+sJK+OXPtC3ZdagBlXVprbKiNxP79jHlknKwT
LlwlVIGtaiVNm1FH+V5A90g/lKRkv0TBZPTN92NwUan1Ymz1pO/oqLNkXesLdA59
6k6RbnSqaSM4NFNhF1OdOv10uLsHwGm2/bJCUsT2nawOob/7piI+HxvRkq6n8Kcs
yDci9UUsvUe13O54onCdwmHznm2vL8qwltjgJf2fN0KamkwhHuacUiKKhIkoXCqK
u0qUIkYO+XCsuGm90oX9dUuyf7pJ5lxxbP+AXF/3ARfhkg2E0shMXOwQAfKbgYcq
xP9RTj4CpQOPLU4IzIUKk139mkTd73rtOwZvY/34IBPST/9ttZ7ZTD//nruy7REH
lEVT0tiZxgZ7BJMfOG3fe+dYq/0QfBMHw1Zc7qcBGgP2+eB3HQqlKMctexasgy4f
BhBM3aczC/rppMbg16LnNahfwMhNQXcZ91VDHDS3/7aw7sWE1ys8I6huf5DTppDL
oE9FQ/JjkcXCIdU3dEBIkwJM+thU1p7gXGRNI0sL+7/L9m6Wlk508Dx7G7BdqllG
8L2u9NeTfii57u6sX25+qh7W/KVvy8V9O9GCOdCVMitVXrACwTzYt0t9g5LrKuIr
afhmiA0CJKTBR5lfSouPEpq5B5BB31mISjuoXKtSnCBARzf2K2fvE4aoOMJE0Ckv
+p23UDci6C1kU3jWJ9dyAKnyVOqHeRVXW7ZZCPCQSALlWqERvcKOr02YahQs6Xg7
vg4+V/Q4FKoRVNJChbwMd/71klo6TTnWtL0t/EkSNEktWcj+iCeHjOLGmkEtl9OT
hiKLX1MdR09cfMENTP+Hwlj2RCLU+bEMoBF5gZCM1KkDrmF/Y3hYY+QmWy5ccroM
s+HQWdy2UCAXIxhRLPk0n9OzFUaQ0eh/ps7MjZUAo1n39FZZG02YOUf4C26tFTya
mzsHmF5E67z3IMEw5vhKS7Cyk+Ksepz9wEdzQkc5/x3sRm13BMM0kQ3MwFkyTCPb
GzT0n1J/NXDTozMMq9yWCgyyt0/sSd5kBKBaVt4MCM2ExSrj4sHn/bZTRWK/jUFl
BD/F11/BdORtdVG1+se1KBptY/3B8k6uWpZh69Nc5VJMAIe2ucjcRA70Hl6+l9Qi
EBL5HGk9GDtvugERyMdzlqQLrnLCfvNGCFUIBKaVQF6irLH57cUznwKNOQJ44aap
ayD2NxEV6ELpy0ImAEVnKICw1GOSsb7IpJDDoS5Yv+6mmMv4Mevb3qYGVkyOByNE
LDOubqFeucUwNVIsTNgNIAt4YgTbvu6btYDEAefhVsHrIVFisVpHucVcpb04rIVE
VabOYSFRUpW6TqDaK7OVjqMCDu84CGNWgRDNUxIh8Z5jcKJo/Kh2GjIe/aEBc87l
vp6FD7LIyWQXph94wnnoPwLb2F2Hll2nrn2odrrC9kDjpAUKm2lJRQ5RXFTFv3B8
jt1Nrf/FZBBxXD5lBkJxzoPaU4ZiheWVSL9cYWKOcdiuGvsTTfKItRGGdq1N/Io6
MPE9GS4He0QGznthfecLjOU+oP4bboE7J2hav3SxSdi2AOLZfuoyDPL0K3EM3tzJ
SjCkAgH19EagOhibPmQEIunNk51pyWkn9sbbBHQ4PVWTudqTrC0u3SKTgHXmXlbL
lTGxdgW+PPQyUHQ8UQ+p6WGoRYT4cLA8cokYvO6Lv2uTRVl7ieYgiK7mM/YKfzBZ
6A+cuOVgiNCaA7gOiOQaSXFJUuOe1uVHRQhy+AONP4zvTc6Mot/UOMzvK0m7hQwA
dbOP2lb/Gdmps5+84OgT9TNBQCn88WFGxHo0j+dEDlESaja9bp8rJ5hKKQgKU4vX
5QHnNjeVMfRz6IikdG0BE+ewuU/zfXUl3/HDw3vzZgfNWueDKibYdsEwB7XXJWyF
wRrCfe6bPFb+0P/D4jPB4QEwyfofPv3LiRWmOoDUzckBYoSBb9LZFZzQ+ZjanmjE
Z0oo300Q1c2dbW4x/oiv713+NJzZa0Xy+jjjnBl5AnghuPiOMI5+7B7yZPHz66lr
rvRhrgEHnhGql7KznR97/EMBIcDYeGo4FmdeXOtRLvdCwKrPfAF1e2Lu8pUc9DL6
qUxhJg67E/QGYnfmCc4m/KXhcuZ+4JVEJQ320zkOE5VmCiiuSy+7sJjmwsoFEQ4R
esDl2qDyR8UBFTcTrTtaCZ9ojiNhe/AUC3Wd+CsjRwOQQ6AHfKtXfoqayGY/6X9B
VHswQL/QbfEF2Tc+akxCPYJXyN9yyKLcBrMatYHJQ8ktqRj38mCmgz+qHkVTYO1y
tNMOtOD3FqjB9h86eFbf1gSWsuoS+OP64X3dC9aN19G/1tA2AxTKRKliahh3uExC
uOFAOWpqqA2c0lOzAhPmT7KwxBlxfmHtY3swizpGRO2LVfTf6c1w7mHWI+FFQelZ
mR5xwskJf2M0IWS07lRFrq1Zfcwhy9bUrN5S3QBDJA+oBDRpgtlASlHeY3ijsGZM
zZuicpwC34NG9wJ7PWK6tMUMELlZ+CJnRLQs6i042mgCt4RyRmq+7LtRCatfoxq2
6kIWC2aXHKQd0APq+wmqJr8iN0i4gSEQlAZa8BL4f5J6bzoU+tD7CRtfoCrVnelc
Wq0Wnh8hGiqzdO7a6ZtHcN8fwlq40iJuMxz+kBKe6ZYneAZjvIXB+nlKAuzvuuwV
igX3Wu+MlTqViVKG+Zra3HXg7kOPYRg08PVEPL+3P/jqi6qPPwdiDLXTL1MFEtwm
IvM1R+RJu+FtX2W72fLH4NYHS+B3FDZuEBxW6wPdjvB+1E3XYsAUvn4yLakUsy+6
onO79Jw8xTyn5LhDjylgP7RsrK5jvnSc/1WWC5eY+ARjju3c9SS5surywJl613N/
KmcxCJ/gxGRaDLJxq8MTqs6OUlWLhCUKniLJiE/LU+OqW2Ibi5oRaGHW0+GVWER1
r7grV4HLZZ/ZGJ0/5I4KuM2JK1rig8PJZRCEV2fO4bMUEpyStE4d4f31N+wJUgwf
ejI3le1XjiZwKlnHoOOpbLXA0RGde1mh+61IbIEv3EQtjXcez/9bbcok4nJMxJly
yxo24Ev3+jYVA2Fl6xdrv3rMHJqjrNIJt3mGpH9heoaGsfW+oshPO4UURF8L2f+8
3wVqh+paCmVJDisy3lV7KdilnW4rpaQL0vTQcxhqxTgKzbU+l9sldTlGEY3mJuek
qys7Kbe8VUEAv2THYH+i/22Wf1QVT/Tt/RGGtfjaIJKEMYDCtgfSURwfFC4yPAPY
3r1cBN8BfLCM+9GdsYh5LGd4YqvADvaHz1Vsll6cABT5XBmhuww8qZ3dOFtcDQ2z
YTTHz0uEvXV5003AG3CSRMrDpEm5SoCOfix23TxvpuInekAs6wzMklPOdQglVuQx
aIlbDGvSZ9zWB6IBHhEKqbQw4LTwehz4gZizGxH2Oc7SoP7oQ4bs8Yqd3OGR/SzW
qSqyKCN7DYxz8hS3bmUCdfk9QdQIX6An49GkWiEXnVYj2eGAkfdZabxS3u7OE6x8
ip46DTbdXGIrzpOJjbTHdu5jDI/KDojcYHOmbGt48h3jdHXCyd0UOkb1sTWCDP1H
xWacO0Vwo4V3+i/cCTPq7w14pEx9mNF+05ZS+UkDeiGj/0gD5xxsRDYYhIL6vg9j
b9so1T0aWkXYLmCZj59VAilTIJkVSF+7IQJsDCnXrIvByIIIY+xna+ouKoZosIXu
Ec+0wruhvTlZw7txh+EqW7L7k0GVfyylGnx+As/rajTjMF92Ermx8EZSnrpv7/p+
EbuL5yDSVUDx9ESPCtGoChdoYLe4bN1toij/VIpyfkgQnUNx3y0Z31GplR1PJDG8
l89KfQX7VWPERNLkgvfHIzS0pRLoukR4mTntZK/1ISpUErnwsH8eqks9NYj8gzFx
wCQMC3ZDNd+jdr1Bit56kDb5mD3xIAUV+FhN2kijv0eU18BoRk18QBLmEgaqklDN
+rdt/Cwsb1Vs1fIvAU+0iNQrUyEPfvFh4kfI08KSwFAI5T0Zs+NwJqp9CksLIVnR
cPBNmDW2LzLD9M2ZZlnFeOkEygfAG2cgNOfaIM8XnJ9gD/aJe4zNh8X5k552/i72
Dl7AjYAgu92AVpN9H3q6dNOQKFsnJ8zikcrz0wRLpg3P9//B8vTL5+nDZLcDfVmd
lkZnH3PP2zLECOoQW80Ll7DXbaiwnSH7xPsZiHRZvjq6CEZze21yLcMOXRV/XaTv
wA7feZnldhYzLYAvMSp+nzgEV3bjlZXpFmtXACTd3xOo1OaFr4KxRpVkrOXroOod
OyBiAewxvgAamCOBmMF942JsPJoVtTPx1upM15K9AiskOpDzv40ZGIli+EUsBV0U
P4qWnTAMcdEdg+pVzGiVVKz2/277Wzzg48+FCHV+J1bPhwhX7W1VE94Khu+GaV+b
st7kuZYVhzNkz/4B+3nOCtX+sQ42nSwa6pkzM9KSdJvIASgq1CfgLIfEG0QHbVJA
sEOqj/FNpcpdnYNQ9gdAmbrf5ZMB3kJ5W+W/BnCkbG/57o6vkPwDVmuvDDIz6FAF
dsihxGXm2eBGtOsQeLABPPeENEv56j4iX0Eeg2Fx5nMJOEtka6jr29BQwew3lFh7
16GR/HaHfin0oPd28EZmTMvyXSnvggisk1hJ8m9WS4s0lLbLGC6tVn/YIrowG9GX
j214Y7B31iaQd3MPIpTdvRhuF4xOTAKhMYGHfvXewFnRubMwBDNcQmsoFkifOGY0
sg64bxaSQd7c9wb4217BUvRdhG6LWCo+usEiIpwr4xHXS5QX6X2x90lpjhUWmMAi
gWJDk18tyHYq/1BfdKx+j1FPWrxWy3ivqp98jqpkDgpSTv5SHwm9pbIxuEH5Ocwq
rF8DRfbDCqDPvLPoy9CaE9AuStFcKbiC1Om85MboS9Z/YAOIRGj88MztSbdHun0E
8zjY62YDHAE14lSNN0H0EHuRKpcEvaD5rB/3JLd95y0+kizTBLqt11VSXLdsIAru
giROzNFrM6GfKtBcdM7PNBww6A6BrgQzGfS8q20ck0pzRcUmSTsXz8ji1Pah1Lca
KjLdBc6ItsUnjLxsrRybP4+MEMcHgbp9yxSQe31mka9p5tRvjZtvVYdJT1o+iyeP
NkTRR2D7hfEfNORm+USSBNF1SxPttZAHhHUyzkgUdyZMT+6dKVK36vGR+rBetUMh
1dTmmscgBEG5jGn2LSDD+iNFNH0/cGiRtxxvx3vkNLc79h95bPxpXqDJ/cl9MS/3
hbWIHDZ79BPOEHnKaataTh5cMyKD80ZKh/2RjrcVibW39xNtZqs42r/rBdSBTuaS
Q9ZAkO5hZIyVT9d/YWtZ5zjAw49M2AyFzHQ6dblhj15HmlY9xfvYrzbL+dQKKwbH
xUgUm2em7xl3ZaPBqiwckTgtbiPyG4N+di7wGZtRlxutjZ0AWd8Av4AWoFMZ47Cc
kSMzyLzVIfROmcygwhyFMQif8nPGeHQfJGd97Apwwun1gDKVlQhhJK8VssIrnNgw
Ol/cbN9zBxXp49aWXBM7M1SAQf4SnhaSXgh/VK/TNTrfnVkPyLQvrq0Yal/kDBU2
vUzArKBzwIBxRM5gbNgpjgZ729hI4cmrFWPhqXBC1rc2bN+/F/jLsjiTDWRlWgql
eETiGDg/Cay8Ygi2Mm3sNutcTSZRvMX/KeYvxaOMxboOWFmRk95ZZ+5ifk5WeLJ5
SkZLlzlf5xvqpK8fkWEN8dttzsxUNznYxOhW13ISy+IvWFe6WNOxVjV//HB0Q2tQ
ZCOOpkDLysauA+9xgCsQRHD0u6cbsTllM2MG9Vx+K9FZ/ZE9PclxLCID7fjW/oxe
jmm48Nf8T9bltLM35VeNio8z5OfwNQHzYrxMVfXcjA+KN4KJf7A2PADe8KstrUzp
ZdzAYpvfBsDQCuNr4dKrTx7gdum0QHCIevCPP+75o5UCvaVGv8C/BJkWoMBi1J1M
1ZNal3ZA7zdubqUNTdfaOuT75Hxk/+d42QduAdDILpNTEkOFLnfTtL6sP7H73dkS
qz/Uvn4IBBW79N2dERfl4BSgjECAWcUQ9gwMuoT/3RPHIP+3zPCdGS4O/4VYUHdD
PHkYVmq0qx3xrU5Qjl5lUWBBcdcYKuMPEWjB0Eohuw+nsPteazqN8YhR+HPKBvJt
/57FUtusapFYZHVQcJsIJcwXWjc9LP4ytF5ZULru4cNsWM1Wo/QVsCey1GFE4jh/
xnSBkvQKe3j1zX2bXrmf1dmjgF8d2jmgOlq3t161VnecKoa/rMpplHRM2KhSHOMq
scP0YoJ71x0FSBHR0T9B0KTNT3WmZmq5G5lEjseCEHEP+n/TN9QGjVpn3miQ6Nvc
HcHY1aT26ucc1rUWTZndlj8/kVxKicEQBCjSINlrgF19ZtHHjOVowfv7XB9JTW4A
ExjvYD+mbKQ/Y/yQGPtOzEywqpmF0ZEphonKyUzKc7q/uOOpVhrNkaRtjShs/e3M
J1K9IW43/HDEQhbPcdK1J4ueumHpt1GM0NVhOfDBHyBP5+N0imD/z03+kZ0JCZN0
OigqC884l2nuiUWBDRYFEFKvq9QOjb4MNmz1e+AN8sGPOW+Hiv+NStdgPDHLX9fV
2jTa27MyXqFRYcj/RTRJsKlLwR2F9qmSiQhZfG6KTuGwVaDJzswN9KXW6mqaWNuR
aPFmh8mbqJ/dj5GrvAHbr69Bag7+VpSCEZsPOSiECpvk9n+6deqopKmIDpuOFR+v
aIlhYzURObfSi2ACJ1qRdKFo8cKhlGyC3yrn4K2H0oVpOIsXVa3C4r0yExUOVlTk
jtUWylzhQxtuhC7PcLf6iJ4J0b+EASjNHWcqaZxrmMLE8ajx8eoKtqIHub8oPuPw
C2bKTiPBuaa2XD9kxGkN1ByBN3Zk9UtzcSrRR/yresjeBv4k8Eel17Oj42pEuU53
5JWF/nKFq2QTZnef/vImRacI60tgN0HNUguN3+GktCgDXCSmtg1pYYPF1mgsbvbN
Stg3Y7nlaXBhI6jBGl22RVE+s55lcPOBlcPPDAdQ6KsVytXCYqb25XJXNraIzPx8
Jc6DmbxbUkRD9qagWZh5hOHd+DgNEO45c5ngg6NjDF1oTDcUPjKhmOWFyHI+kDWt
QVpk1LbA7ugwhvjVfrCHNKutfSpFuQGE71PiicmZoIXd18GN1b6mMA1dvzAJVxGg
BonNSRSR6DWOSBYKR7Izy9R2mEV33Wnnx4aK3dMLUKJYlx3Ab+SVxxjcSq00oNGS
FYfjc+kBqDMnUiOto/ai6i96tRFkHOUNd+uGD8G0pJ4o8RQ2HhR+rLTuJ0Gr07dx
gAMcNgxtpvoq3OCvpXgdZZzRB39euWPW46M432wHWWuCmRIKfegx//NoVISKTHCG
MW6A9iIuWHASnjLz4yV0BG7GkZwen9OgZOXS2HM1p84vJJU7p/9irB7VnJpP01qH
UrekUQqGk+0Mr0dBxwsmWiWXL+Zz9cGD5sP68LxwzMcmJm5uGmyHgx+67OcqHcvT
WdbCwu9xCJnEUryDJgyMxfYQbG2KI0HFZ590TU/ynWZLOH40fGevdIpha0nasgW/
7l5OR0re81zi3YBm11iy/E51l5h6lwltxuHU4azAyMpqQG2DqbbJ5xiaC/OVEYMP
s9rV8fObPXgszdMudWfzexVNx1qa4HRoa4feRSrYRLdWh2yV6j2GAWl4RCKDPNeI
P7bY0mcO7VgL5XcrNgQIv0+eMNTqda+w0PFUJVROYJ3AL1fLr6VohPqO1gs/pccw
x35z2510RG69Rpr96dMeQeEArgi1v7sQrCf2bWACQpoKWDSH4IoTu/lU42hHiKCc
9+9EwQiANaykBNAJP/ha4s6HTlvfQE4ji/79qDAC84yGx5CxviyMzCi7oMQYkP3s
/uoOuzrdhSEi7qbpNM1GkXRM8pQziSQbvAHeLx6oH3Q97DAY2MRVuYqA1LPaNx3s
cdHOtsiVFgEgmXzCK9xVI+9M6srb3G2c04/XizDRhjRh/e8PhRyA5pbzB8f4t1o2
43TvlY1haF8NX4AUfK1ACZ5Q/QRJpRMXE69Y1S2sFxShacSy0Cv+7nSrU0Aqa1+u
b72IYEZxlPxtxeOAGFxUxVK1IstQlYF3Sb5i7lXQWqfgCJ6uCrHKl9vEswqvKi5F
uMhSUF/dyVWJLRrooV1yc/k61NCam2Fl+cnNha2ZD9TIY4fyQKDVOr2lShwcZzcN
1C933SWPuYpTOZom7Z3RU5M5zb27O8C+j8RkkltyeYUAb1ijadlXP+bUANynPBrz
RKky1NAxED8lG5xDmtEImeC1XfinG+Nt1kRQX9xoOb662ByfzyrA0TtLbt2EH6nZ
NBEG7c3ErPlkjdmAn/ea+9U1DQdSkeEXh4jfbXsJH+mllv7uspj1tcW7u9su5emp
1+swspfuTROM6mhH56KkinRzlyqN6umJDcMiKm4yAZ3CGTaO1yHu7sg9yZR+CHX+
XWgpQF0xg7q6IwMLWL3nCt6iInAOLeHNwxzfJl8Hc+T1R4YmmfyxkHdOL6UgGR0t
xM9fC8UKV1/Ppk4MShRs4qRK/lUSqvLCRzfj+ewkCUKJtZaoKvn8VB6cP2NGmp/+
h8IBnN2Pvgubm7IcluzAhdXoFlek7z/TFIimu/Yd7HY3xnTJahG/8JYTZDonREuF
pnA+vX67Ptvt7ai22x8s2ToTlb2SimVmbXybIqe01mJuduZZOy3nIcK2qeC0R8Lh
3MJBivw+X41PXBNfqkhTjHw3+UaQiks4bXG1ZeJNzMN961brAhywbTjP4Oi5iaKR
/gr3Hg/AWiI9VnOBAjo7ZuIkrb7DosGLDO9WlM8PjBf/RBW8D/ZC8IYVr2xgKb+0
NtX2qm67u6/fe/S2pXT2ZwRVLAWu8/7o74fWpizslSJehvVFe5fX6BgUgsFf4Av3
CfMJeyveGXw3/pSzaqn1jPZ6E2FStWoNwI1I6ABvFju+Gwzez+5anjgNLWKGvatn
oQGG5Hm0i7RiAvxrPYmyH6veHa/8yGKX79rHiDmslCfnJXeNY7BSrMFHXw6qGLPC
q4OY/uIIOPz6TKacTGB5C6Xcc39FVGWtzTLuPA6g5tfKFdocBiJfK+TUNHnL09K1
VWDI7LHHgg/LUSLP6Wkig3PB1Yqx/763dBIuJg3jWa0ds0c44qkg3C0yhz8TTZLI
kwlDYk9lBOnwwgy7LlVz52vpZOEiVo5+fhUyc8lqde26iAQWNPsomJ0cW5vEp8zp
n6bgATKhEgjjEaVwQiafF+6LPat58+txmxfL3JhHedy1tLao/2TmSvoJlf4LoZgY
wdocgqN7OK+sdBM7wggjTrRFdxJ2zC5N4gZHk7DDzrFZt5zV4oZtzVZWX1EMbhO0
Ffzm5M7Vm7T5E6Iqxk7j1wAXB+r4I67CBzAXDf+1V7eUA14WaIZuHRMTAcj9A0LG
WDL7mJ25ddbKmWxvxgU7vPd70BA6kGLMp5qd/a2vPnHhuTDWK+9LYN2lcok5Uzgi
IraRhcX2N+eR8nh08S5NbInbYBHYe6VMJT6fBqT8+lZhm04IdD/CFZNriqXmGZPd
hKioyhYnnZkpOoXzPTipJs9RESFNLkuqTIKKWyjsJ3QYJts2HVirXAnMgrFwS0FF
jv1H4oSK1j7LZCe38xJFGqP9ZIYUmyTcAxbVRM0nznv5ur7ObBrrkIr6Qh7UiBZ3
O3s9rrKEn3WLBviJu/wI7nfJ3pBgcqrXMBZaQyr8+KpN3RqMsiIwKua22PD08Uq7
MxCZW5tPwp8lSinBOM8YJh+yXn1MRU1aXyvQ754/zQKK354/udOvB56vDryKWoZR
t8OuFUZyJhiEcOBqaNiFY61uaER75rCjVDIejBkBEbnp09EuIYrv9hKc57KvchLk
hgwL7+ObVwKZxqTDzJXv3RglpmbyEzKATJyLzMK+sGAF02t1mDdEFh9HXXTd1zRe
V4OFTvYVfTELiiR64Z3iAf6+E/Gcfm6apxwLUN7LCPKVAjkp41mOlFvhWg9hrxnY
2Q1AhwAkhiqE3wVcKLphZ4MUoFd2YW/1NHINp3mZGX8+89z5maZf3umpTKn2/vj3
AtJlzY2zJMOOi4WDKVmT8CXJEkSo5F8SUQ61pR5ycmuG7y9HLOOwyn5KdYAX6foK
7SPenqKcqEHITy0+CtdX/nG5Jv7Lji8IarEvMevK8XtojeLxFH67UoiYEw8KtO/b
O1vCc4/dboBIMRkID128nHMlf9c1tHqaul/PgdXI1AY/xPKidiRi74VPC8P1wcd9
ZSii4DnuRcaISrBEWIj4FUnGzm9HT2/tkAAOTWCcLunvMb8gWZv8xaKCW4G+NbiV
XKrzkB8qz6CDS//uFTTw79jxjn/992fWjCH3KS2q43Wtum1ij1EF11zY9+j1BADz
HjbDg+tiz0nhnYg6N41qjN5KL+618ovIP2/a9H+r47k6/uYHe8zESJPv8t1N6ies
6MqM/mBJBIkqkuqEBqhAY2DUdy2seb5BT0mixDa0k/zjSZuggeRMd1pQwbBFMwgB
mmQuXWBZGFsO5Ly40OQ1zqt4C/ifojWz7AkXuCBeSCE4dfw12dux+85YPcJZuIJS
dGVYPBWLBujYOSvDySVDG5ydjqODAgZ2PnLo/IK6nO3aU01jdXQ86V5DYJNbdpFg
d2DEQCw6E8AMrcAa/gS++uXD2xSU4xFABv8Zmfva6VMv8xwCC2/c+r3NDFuTsaU+
Nnrz8fIMaiqre8zdELTVBBqccAC75/+qI02yOsWZWH2JX40TLLzo+Jv+AX6OCf6V
PdUFt+rh0DkITXbp4SgbRcge89uRqrB+DKOnAVdc2iUB4vhS11wvZhXeoGjnla7R
iYx6dgrs8YQlxnznh7+IlNJi1Q3O5up/Cjy0CPzgv/QTPJzpnfsAwUqhOEtOKNCM
aCG4ZjEY9PNxJoaMXkq52vavK96oUZn+cJ3PdMkFrqyl8y3vhHKBlerPSEGAXs+/
8VV0deh5rrD1sVHEkXBfKOkbJYWNy8Uz9Gza2au4Hj3fG4nTtk46KkHLDD6wCt+Y
T847wKCScTtpCjKh4vYAZ3CSF/NH1lF6kWU70BPzL79QsEXJXi5iFfZO7OIqFuGp
ST/1p7k7khf5yl9ljVETW/wV1idFUFO5Hvupk7+u0g9cblHlqTRAu1WYZsqiB67i
IxMqjnu+j/QCvWV11iIb3sreR551EAJv3DuOv48cnA3iqTvxS1+2FhcXFYCe5x20
VOqIzqie39bAtUwvQnTWCp5+5VbWpwZHfH9td+k9PEGPGAveL1hRdCS+Nf3Hbiin
kbMMK+wt4Tu+bG1Evh8fLL/zbjsQgJF/cZC7od7FhpvNGOXennjfXYgXP0Q8+euD
g3jiMQ8arty4YUSkbHeI1ThqyuYqF81Rd1ccozqSUIH0w6agY9J0tlW3tBMsYtf9
WyFxHGj5p1qaFTCi7fwagtmMuZtgrB4J7z5Zupa2+GeARabTNbFxs82aoaCv8FKL
YwGZfIHZWrIjEU/C4wUKhrescSs/ZzEGKLu0YU1Cai2q6Eiiy+t6jNolSHUn1oE1
wbCPqor9jjBUv1IMmmHzVK3HMMvdHkhyk0TShfAFA8mcw5EVKuPHDo0SDNn43rUv
LjdANJy59a4q2z0KJ70AK4S743w92Wz1iIw75KJwXQs2GnS9fiZM8QE4R0WR3jPq
GVzPo7e/6F9Z1zKOm1z3pL1s1DOptFZbx9CqGLBRD2jTt/cf74pRRi8WqPdVwtxg
Wcac++rJqpea4z1DUgW1gQwPdWn5GBTdHyG4royOgsvNpnVQLlnTCaYdCZMQ3dMY
eR6FNrRO2GDVaxiA43qlud8R7MjFE/p5qm98lwvePsVeQVk+od0abpD5QgLj4Hbm
kDBpkCxx6AkzKR92rbEduP7xupMZwkkTdUHHZnBFsVysayQrNZmrJwnZO9GijDd0
oooKNF/aA4tuC4WNgFEjTIdNek0fQB0d0CC9QIHK+PKvPbd7Gyv3dIWRX+iJl/+Y
Z42oRdFExymYyZNnu4sdu6PEbef5yYRRvguhTMrc+cr/nlr13wlHSch6JIq8o7So
zFo4KcmvYIndyQ7uB0ls+94giqVEeKf28YFvaDlwTwvFMLVn/ep1qufFqICEB18D
lrHa0djFDvqJE/0fqMIo2UFyZeCO/blnCUqn6RsAgQn8oQIlmmaTvKwPe1iEIOWX
ciD/xbwmieM7oX0UcPwQ0ozzl0v2u1yr1iLjtTeQ5u17PUjhZQgKswjUOkGmlaFR
unXdQ3UUsAyX+IkDPXzcxyr7WqjoPfoX6tradSIZSCm1z4cuYuU28kal0JGSAbDs
CAzPj6iqt/9xsvMXr26I5TC1MvQfyas4z8gHCdtlItZ0V+rLt13Tx+MovcPge4Ki
jVsU1qphYWeOK+sKAHpHRqhyMaRmN4v2oBJwsJzuHqvOWAbc5J7uoFre5MzD7FEO
fBZ3BZrIVLiJsVEjfbQv1zbdj7DtgXZwPmHyuY+4wTMV4NU4xmkAJaUAV5qd/TeE
04xuxJZL5v+vkxS1sGb7QGQCk6YDdLL5stZoUqm7VSMycY8VfxOGpS9yrdYHjSiG
/TTu92yLwJD3JFoYzfGpoGHTBhaasR5phWo+ZAOHF4ZtBQhokd0WQbDI5P98e/WA
4432D4DGHGmBCmUR/59xr/H5rzAnF3CYTyA1MWT1LXBcGFYy3yi2hRipRXKvtMfU
WnP1wazpDZMBN54bof0vw4Ol6kDZPFQ7nLJJkRR9ZqsJNOJBKdrwlpOf9QC4oMZw
3MKSKGZBLorxkGLLgQLX6MUv3iPbzw4HY4bAjg0O3AoPoAxscobRcwnsy50EWkJr
agp3kvdt1DHZym6fKnzI5dOk/4gqb/LRfe8yIK+aRWODI1powKxU60GJf+UxFw3t
hrWlvHtSq5vxoIeSEzndo4CUvEeofMw1t6ewd6huSMJsf4yGlfZLZTrahXvTt65W
ZGhmC0+QRy0R4fbW3w9JPT1NzOdxLDfj+aRnsAFkf9CC+ji8GV1SgYREYzeczEBy
DV6yA0Qos0+pMAIBVqEgL7JTUzAU3+8n0OXzCkfmgEB4rBeMgtHOCXKIDKlS7ZaW
ohU9C9BI6KOap+XhGZPOgT97/RxVtZT78TazgPSSZjkjnHXqVhAUryHLkos0B9zB
khtnos11hnovfS+yC6f+ItKxR33daZn4SHeLt0zZp3D0Qtswu5YxGrvJKhiIgdcG
n5z8s3DwiE3PDaMmW4jOfD/2gvobybKBeTxoCDubQdlxszKoi16z+s7ijtpAtM9O
6IFQ5d+TFYIfHbF31vKU9P4chw6FSC6XwxWVHAoEJGoMCSlbH3yhVKEJcSuqkGez
qrhrliXmWdrbzKKVALN8AMQKh3NxSHzuBlMHNXef9BI288O2YehMoSox1OH0xLGu
MwBKkuOYVQ42slpPi88ilOnBQfkULWoruMixvfVWLoIi+39k0eB0hwIh+wrSTcAj
YRVHAI+zBVcHY8URlfpLX5/JzdrnYNq1E7Yq6EMzn5fOBbmOftp7gNbA8vaBbl78
Tm2Evl6SIhmNkp5GH1zcFQA6UOtE1YEXwScTAni8nXPN1RUiVyAMeyypV6MkSdr7
FfiljTGgbvFtcn6FIFFD/aCjuXD9py8XEZdlAU7JkwvQt/5rlO17vj2vgNiqAS7d
hQAHSSjuMHL8rsVJprO8J53ARTQ1C543YwaKZRrqymOb9UEd38na3LwiMb6bEvKC
5QS1uDadJwfgruUKRjtHKRIC6v7Qq1toWKcgBmQrygYr/Mofl/xb0X3w6lNjU7fl
bT691zfpx2Sv3CfM7JeKERq3nHEcGtjoevCLoMSnD2PUnmZLyB1uthfjy0UnopzV
4FCd8wRFHFcF+dcqHQ0v1SevzIUM9vbccbH/1za7mA7J0P6I3pP5f9SMk4Duo3JN
TfNFH4WQBqUgZxSe9Kjm+WxqtEuOCXzKIs6iedSDHYlw23LrQQ62ZIIBKwP7Xx96
tCkfGYr7nfq3daJgem/fj/yGYCo2k+oGoD+7UEWkL2vGQQDkQzj4P/GrheUqyOEa
hTahxWXxzt4xYg1HIXFPCgItA/K7HWUc1n8/ei7Frb2hmIA145tCfccPg348j2oi
gdbeRogCniRq6s+uhgdd70lJWy/iNI1XcDzGrkaHlq27DcpKVOzXiPATRZ9eJM6z
Dw0UqHv1J5d3euRRlBJFIqI7ELUx74nBw8Lfca809NMXuI30EONPXnI5xY1A7Fzb
tuFKq/kLZwCSZNTKpAiFQAoBKTsheZ7+pmPJKZHnUkSuyiiTc8Nq+AfOxF+bUirW
lBzjfQ8EXBuwIvjIBwc8VAccRFmGhPpfYAegusr68ffVU2QbFAVzaTQziJkm3aYj
PO3Ymc0cjrqacvIXw8G/y3emIVQWV22Gh13iF0LFxUYFhWbW/9XzoeX6W9yr05ux
fB2rI+9wsuspMVTivpGE2DuJVbZ7Veab731ktizNa6AjeYD1NQDlAkEqCypkNlWS
6YMozaBLLrlQCBdG7PalCejuw7nXNJ7mSJqO2UFUeTuBok/H11Q6qT3AXzlSo9QB
4AxYzy1Hlda1bi6Ec6eO0XHk2fZoSV7cMRyrdSM74BdsXKDdWij1ikYZ8JtahRGp
hO0TH3I21pn6Nm6A05F7/CI+Za6S/GPkgSODEnetRBj29Qf2uLPGh2+aRKwfdjHw
LF7fs9569eBaGc/TB6Uj5DflpHOtwHsmeUP+0423z/0yJscBbglozm9UFB7qw8/w
9g/PDxqDpYBYPKTNkH+bg/M9hSTopVY+pFa6KAFKrPJxNa7mxqSfocUeqbAwhFQa
6TBOETArjwOEUYXVZ3FA6wJYr0rmz02HA0YTG9wXO5lXhz5z8QZ3CJItWX/br44B
3puCIjT3vePKPog8t5gnuI2YSJorW1pIYA5m0FhPR4Rm9m+if82bOsGHSs4sXEwK
H4lgpkyXmoF2+DO3RXTEkY1r2ppJeJp9Ru7BXwJRfwPGoImYgPW5mXEe8ASSZhTm
UqIKgBgfdOliu+a9lsRQCDQDC5oNpF6UffxI8KCPgtskudOl2g/rcIVWyL6UWE+l
KACYLhHNxk+lgEgDUip6eQbTddKO20XeYmH4poCYkwGSiwW1ieALKSwE23A7wTTv
qObdtJs0ldcbakbSZM9gnLH7vnwOOSLtU9y6sUYbTuYln1iMXVWGlxKswvEfNeay
YIpP3Onpa+N83X2v3evoyM3He29v/1vwTnxTB7AbauY=
`protect END_PROTECTED

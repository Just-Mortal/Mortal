`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2Nv52ZOqH4UeKKaQR9x61WSnBZZeqJIc39c0pwepUYman6PExBwNHyViyAPgRl/
+byXmLDdMlfueXqp7BqFxZB/oOptBYKZiLSuqJpnhdS/V3JM2W3XdgvWW8awxZwn
zY2F9FQeJqTZ2WvBapLf7kMIpWQJoYr4WV0a0UZ0jNg1QRibU+qG63rVXsLChSLJ
RE6pLftgU+LhX2lX6Zq+dr/uM3DyP4FY/LxsjlNv2tT9Ck8ci1MILawtZWg7az8h
81QnLt6iA+oXZUV0u+ptc4awuON5jhdT/esOVWQfYPvrO+vN8r+JpEZXoJZ/ZFMI
3ObmmJ6izsQ+VElFliXqw1795A9kFe+MI7O2hHJFjkUEm2QZ48PgRgFOHRhjPsvw
a/gIlxStZ/hvmWOmyJn6HFjKJJkbi5YWD+3iyxkunjEGrwjQAKCkgCm/ufDKzMyh
HccgrC6xOrFwS6QiIo6bm4J+Matk+tfSeN+EVxnE91x4ITL2Yj2BC2CmDoT/JQzM
IVyMGHUgXNGUAYRFahoLHA89WGCg09uJw++VgDBaWW20CUoLDxYIiVsE4nWYQoys
F9fYaXGa6z46vvNTLfar+PgGmBdgOzMpF8CecaZU38X/2kysAcWPHvMHPL2jyow2
sbEKD/Zl/DsWTW/ge46OXMwZ/p71fFHQxFtF5HD16U68UMD2D4NZIangqBzVaz3s
73OP7NlPVJBnp101bBOzzoOWX3M4AtNvMk17DXxfuSY5DfcaMWrTJV6l3c1tNG3O
0UBvaoRFZx3Stc/zaeCmZaN50MT6SOK37LXp9isoXouoeaSvZKIX9uG2zGoIRtHk
76gsWYh9Ims3F5S+Yj8kwOivIqw0ZmznwMEErmmU8KyUVjTGWSwBCA3eFUjNfqI+
bfVMQP54Dj4wDqKwL4qjeR3IqxBoAFf436UKkTCEWAnwd9rYHMwndXwa1eQ9mpsl
NugnbpFEwSp4DvY82sgCI+zudt8XGqjIM+lWzqXtE0gcHUcXzzTZBgDolcDVodG1
AlHmyffJwvl/e7yR+hqYSPBlnOo4fIp/B0DcLKBBQgzO2eNiyAqlB23ePxDFmEgD
qlGI/lIkASlCHADhsZVcNUEs4Jc854Iu+T2NI5pmjv9+CTmA3siIvPGEUHQwm8+u
97hn201mYSatE/gy/jS8ayfUvdvtcS0AIoKYLZhoOQpS1O4lqhKWLx0GgUe5JMcU
4tA6YRkeduOxnzI2+AagW95vKndiyG36UJ61ZMByoGwQqt5LQ48uCi9TplKFWqW7
JE3zVSSlGqejWCPpC+bWdmktSv50GuvhJs13EdvD8BE=
`protect END_PROTECTED

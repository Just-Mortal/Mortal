`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EygHpGoAQ1lLYGHapgta9il0hgDY2ao7YzouUt8rWjbC4lHxeXCqeSq7Bd4FaQBn
l18Q1ngJbre57DX94/DdQcmPtEZYXqJNMfbQsQ2SAq4Wrko7xUd4UKV88bLRsAzU
rUS5CphSy5+19rMoavcqvmMiCuyCV6ALDCbX7k7YsXulKfniQfvXZTvqcjfl2zph
RB9trl4MdTMP81lDiZodGwP4wpWHn4/A9S1GoZC4nuZnY6bQ2PFr6C2T9U60gQ0g
/EkCk/j8OEkY51E6AjUHz+p3XajaBDaXFFree4djXdcfsa0DIbWpdw1YVG8d84ld
BG9g/4f8uqC71D8N+seCyV2s2H846CYNSrN8REZ+efgOGw/xo2yEHDNBbgVHItUx
mjWh7xMOh8fXx84MIm8o1Z9Lqk4suHl6vr5A7yv1NrDXtlv12jGesuwM5f7h7uHN
hKgfSX6/aWWDIQ/LAwKyqjrWxBLTC5+lHkZJfjT0kgRcQ5SKiawM9kDBUBucELNF
WejwcyWF5HWRQdVo2pglymqCl4nDLAT4zvacbKO+zqVa0mOTApIrpvrfZ3eaZ2G2
dSOj0TzF70CsVCXuPekD+o9nkEuTSFPcNvirIIyk18Obf49k/wYLtjwIszQRqo0+
1EjYdmwJf4B/kRjSmA1NSl3TYnV6qoBKvFj8v6bdAgNNgM0GhlE+XUJ8ITh7qupd
o3ng09ACfrqrY3pbfQ52IOdf7FxTXFkaOEZ+i7KGRM7Yc+l4kffDHqHHuaESTWwV
MFqefNCnr672l0hMHyhlJv0DkLHOVnCaMHY2Uu3JfwM1Cez8Vb4KaCqRphxWSfaE
uyjjLHT/+2r7VNGb9aNeF+EpLEn6QTkCBt1mOR3cmAdCADzl0/MyJ+IUwnmomnzu
uTSiR225RbeZT2oVzEezRu+89bTuNRIuWtCQScxPfa53Kmgju0mxsQGXx3+U4QTv
bKlwi9yM2uE4uwFIjHTV7t9UDlIEjNg2spMjDNxb6i5hAwmnZDbbMP+4hnMIQwXM
WZZYCeuqKV852uEEXcAE6MGDhyEjxYxkZHWbH6LcPnQaYnbOoYsIJ31TkkSpke0W
kzXJZSFaP12WvtJQupLY3j8qQxLeeCl4OQ+w9fjgBDCELR6sz91cWf0u2xJ2HHOU
Vk2GY8ny6y5fW7a943TxZ5L5X9el139PdUMuXIE+eiqWmrAejYm1l56rBBMtv3Ui
2ddwvy/g0nSBN0b23E7g2EN1ljsvCzEdtpv7su85qwq/Q0UEkt7KG49zbuJH/SfU
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8+WGo2ha19DUDCEvcgGsWcLVj7cMSx8yyL2L6w88Ex3vQgc7Qc49UNea+fNggfg
y6j3zpr23MHUW6iJMpLua0H/qXzNA71xwm/8tVHaQL1I3XQXjdtKeNo/s/Uqi0Iw
ldfmv4rMqZBMwuOctNRwbpVvyYnb1MaPKfGkxi5cGSvn3Q9Wzsa3ft11/rpx6lUI
FwWJ0Ct736siPikOewCSNyPG+s2GfomAtqNueH1xQutxvyZ03fbFgjHPnkQxe3T/
N1qzfKosDsvexWeNmAQ7E0zYs4TVA3n6olds4gW9m7ChCSpJzuioNTG0sYzFvgkm
YcedNAHyt7Alc79VO4tWDE0O317Ba177JEbhLFvMdFFgVkwFjAzp1ylKTUA3Xaqo
fJHsTBiH4OALevJ+cx25lB5vja1RIzlCg4ExtnNN8zn+fvQuNBjyCXWrqn55Xrob
ZGcblLLnk4e9hTVtbJo99IJPi7MJBO8miE9NCuWrHJ4qVame3ey1zKPwUxhuxQMv
kitddxY6KQnxXI3LnyeR9cl4rBQ5wAbgYevWndiwyRUZGoAr7ZJPtcrHUOYaOPF4
3Hri22JsT7s1ZTmTEqLHHrKnxdY6Q9eOKmX0T2fxlkenedPCOI1hC9XD/idvDfpZ
CDT71GJI2+V6MNNLdDtgni7teKtABzmhNJxLHecyD4RgvzN2xM3QclOq0cuCtXCs
vn3kR5aHiyUf8140uINIYT/ApJMjWpJr9eB6DMcVK9UvQps8xv84J8xo0jg1RLtc
OOgdxK6zNKSqih9qI2tYSOhP6MXp4IdlugyAiJ6xrAQ+TIXV2YhuY3+zQUK7Qf5+
zZydqI/zZxZnKis8s+4DPzNjW/e9nbPF9yMi9MXA1t8gLeYqPDY76tY1vr7m3+/3
vAmbwMsbQKWrXzJrwHExFv6XRSkBI2g2PbyhX+GVz7dgE1xelUThrGp5QVRqdJtm
Bxuj9NQKRTP6XWpuZHhYj2fVs0Ux2mIxABlcACUmSI8Nt7nW01ZFZEszVanQZWrf
nyofy10OGZWWPRQfMB88Ixyj36uK06/3MxUUb35W8cwN0y3U+tMMpD2MAZd4NVsW
DMRyN37hcdLJ3vJ2nJJuVy0Ql/flYxG4IgRBEUr3oOoo4Jhdos1GZ2b9U3YDgB5F
aJ16EzOLNGSjXumNdpz79hZtxHpeyycO5qt8hpI+GgmlAIA7iavnNURoL2jE+6/H
tjB8vwZHSXbH9WAxLdrv9A==
`protect END_PROTECTED

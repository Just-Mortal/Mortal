`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXLnXl4GIRCTWNqL+thDcnwz4nmTw89wbyCaL0FHun2zHOnXSEbrGm55MpzowMiC
mq8v/2KzqUGLGq/kEhummhInnV15Sc4fbRphsYqIu7MVOdPZQ6r/0j4aWkSkZXfw
ypQ8y/B+g07xtpbTdnc1rzK6Ip+D6QTnuBKCcjPZbxEq53T4FwCcHIuVZZ2ZAYkQ
JDnGlBlVsp9cczhwi5liYZqHEeVCjiP71+hIcgKRKPzzIn3VJaFGUxseMBM4fjna
DrY3gYq7c1vqjuFWS+jEGnOfOjYm9Z0mx/cG6pGYf1WGbJ/5ioXhjOW+givwjUr1
ANcTof8mKpecHOG6250/P8PRD96bgmmuVAV877Fjfix8e3Gw1d4NWLhO6U5OoIw1
+M9IY+/mk4rm9UNCDJjSKzAzasrty/USO4S1UPM32mfJWJWmixeXMieoFHjhkvFN
vlzTq7JPULX/zYSSG3kPfcCCw7g3sFTqGUtdIJ8TyKg=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DSPR2tzNvlLmR8MoO4gYkCcCR+y9+hszHPREOLycBEn3/Byrf2F7nHgbo2z/8cWg
Lw3W2rz9cDQjnO2Snt2WhOKhq8y+0tysCDaVwzPnd3bYZlPwCHBGKFCK3n8Bchzi
B9FKCeM1C4ORyzVTSGSqKHTtSJoStiS73I+8/jUoPwM8Xc5452F6OihE6JPbYASu
pLoDILqt7sK6T5y/8r/IcNBdMTPWNfOQqr3e5NKFTZjD8lE0NshP3RaoFN6rqldj
rNXoT4vRWxQAV12mdv5NCcWUqyb/DM13WDTz9OiL3Ym6rSbdxldAW1Aqbixk8aqc
dOc+1kMh+Sg9UcHwwfeNw+WfyoXUo4ROq2e4ghme8Te/BUDWdSO902qGNGW1QXyG
jn8iQqA4AAL+wf1HBlC/CbMW8tuLPpWHSx6F7fJYkSumZ+8oGksymBlJr93YrPny
mfXp56mCSzGwEQFqWW1l430eJAXsLLGhwdkKuNWup3vejWHS+7hY6Z/UjYhYxywu
PNRoUAILa6J7TlR+iM3NnKPJoJBked0HOw0oeGW0oesIyk8VxfVvHceIhH0lhOvG
d418LMPHHBCXODYypRQ3fVqAcAn+KCftCt2Ob+sI1asbuAzYyRVvNqr0j+iF+X0C
5PPFxMhbRC6wac2cAScchtRTwjmZYXBb4N9nDF4Mfqlwt+ZG/Q7SsCm6py6yoBwn
D6+oUpHwvngSEX6ys/0kzfTplZ2iJBnxuBbwEHZUgZ1wEeKgu0B1IGPi7t7bFZJ+
ft4NbBIIhecfBtaEVRBl0o4eczCIfBe3bb7cuehw/O9xJpS2oCnaHCNHo6krUIdb
KvyCNcB5lcCtk5uYVFXNMWXboBIigLUxI27a2xlpBktE2IG8CEvt5hAl99is+XMq
SoyMG3RuDUsuG3feXmXWgjV+BG7TFLrILjoB0RGoSwa+D+qKZsP9lSLJa0um5uv4
Q6C5hKQkboGi6jMh5X7eXqkBWk49zbh/HJ8Bvrxa3Peyx6SmIzcJOlpaIUtPJt2f
6xhkHlFw6bz5xhCWbjgSc4/NJuoRRU6RCwa1PStNmhvBvhx6yhNMpzXR6S2lta9K
UbvjVcWPcKe5JbRwi/xPbjUa5hjPGLtjXCvft1OB3kdbePKF+0q4leILc8yQnprx
eWJZ+KrmZGVVBeIV5VJjKNQReSw9kLVlWdBPcPmCF+Xwug8mXYjf5Ab+JJFK2h12
iBw/KlZhK265KPiuriqbjrrQPyKXHMOj/PYOI4V+RmEFuyaaCPG601t9s4WKsCW2
1sPCLbj0XF0Bg8iNGAP4G9+azckeATdloNbDgekFiL7CsF5B/YAsA7pvtBpYriqF
h357VpxWlt64QmE6NrG5+Y0CQlybnXKQl07akIdattkzA+ymmconPnFF665WsevI
2Zjg51kOrwIp53rCeARorsTX19zZcMfeVkw+N537ksNvfDRKF8IIJjs4wZI0hCUy
U02EvkJLYbM1Zx1081qYSE+Dn3xY8YxCk9wM+plfiOVCFoGuOlwcx3pVnu3ORZMj
QpzPCOPhRGzQIATgWZ+BBG6Sr1iwgtgAdUdXbjPLM+s4V+8bcpOsUPPcC7fKTCQs
b/GhwLxySaIArwMVpgpTUyb03dArWOqO+TcPbA1J3XT66r8kX6sQd70T/T6e7Nyw
EQKpRda8MImrpHP1RnLp+Nk/N6vdzYCApqCwLLr6svIIicgzRvC/EXW8XJZ1yRul
0yqJdakK+HyO60YyWmAIZpGpyUSHj079nJB2rRyd0wxrru7C258Nq4rsev4HLN8J
k81K9jQJ35SJF/k7YuR9azwIbqKND6VoM3iEHQkNOCDKy5lS0tXbZj4ou5v/Epde
M0vrIsqLSm7kDZQcLg4N326+rr4e9eGf7FvrjYNMnzcmMR8iLTN1362l0HxxM6DP
je9R8War1oXNJtlkkbRCciN+YOU8eohQNZvFO+zRmBQ3XvnW6scykAf+iU6oiwzm
hYzegw7GVrTAH4HNsVzZMmVnNDaBD2ErwTCRtUy9t0Q33BSXI330w6vpyMu5nGwl
dfZ4AM2A9bVs4CITBnhFMTw1i2fCCFK2mQWmQqxQqusfhJwdoS5rPoDRt5rxG1FK
TYSzI8Enj2agxFooNSb6wzACcwuaapQv/M904sO+g5K5j1wPLAPqt7fYF8yBSovE
12dJjmLC1/U1R2feJo4xPGq5I+qz8EP/shzWEqrUW2v7T0azcG/ai84FeAg+bNXV
OCfRcti57dbNYEeZCLHTdVEMVQ7Uiz4PIXGIuOYI1bqmEDXbhLjYfHdW7sN4fCOt
6tqt1lwn932mqIMsc6yhjzHxH6BzJjXjAeLF+bei3PSRLIL6SA7MbxJx9xIFsOmQ
IqHmSW0yn0ZR7HImhhsoainzP44J/n9JtTrT1KI/mkWj7hkeU76m4Y/Xi42fieCP
mGsVv1ESQjZCvWcJ+5YqhiOTvRh9n/BKbo/G0T7VcnT4RTqiWjNEOaOLz2ZHZ9EU
T0Yz+4Q7A72gpQU//nPq9P45L4NTN+xmHpIoEYcLd8iT4bMAA9BibwFO/XYoMWul
T5Anb9D+d0FjAj2ImSfVCC6ugmfigzxSk//vc4pwlD7ZxkMRe7CB6p1oETzsiABb
/IhpVU0vIouuZ75qlPuiaWPQlEJOsoYGVjKDY1F3OUmbSh1qibekEGzpZ9zFZcQU
kNoKNEy9E8UMJlN+FHmkA/P+UpncBP2Kvc2XHmNm+naJQThjfaW7fJ8V2svKpKjv
ns94oWGRBvt7aon6TUaU56Byi9RDuDjLSfhlJ9lE9nQS2X4/9aEEqL5ml5caQLzW
muJ766ntO3XK6picmmn6PEblKxUnJriBYcSuutUM+MeQyH16K+1trDmkg5GxubZ5
2QSIPXJX1Jrbdh3gK3KVofnHPaGZFXILQGO2Sb126N7zBkrdjY6A4618bl6FK1aA
pARIf2nhQQz6SnmGhg9f9rWTrlxtpb44N/7MfgVy3DiAycoGjCbiwqpYmAH9826A
MYz4qEcDe2cDM3u8CYS/HmJiusvv7jbF88/W1pFDcsrxeLV1iToiyUkZh3HXaVe3
kR9BP+toJ4KaExe7jEBrRw8vyeRH30oytL9R7ROfgibJxpGgvV1y/EyhTRl4jbat
lDxUHRx8huJXOcD1tfAEAFT0yAwaawvqRtZSLIVaF49Z7SIvIuOSELSV3EOH5eKH
0xRVPUw0EYmQhNS9c+gWr/JZKe62qXkfQwz8kFno8X7vmI9dI1Bs8c2lerbAbq9H
u/qhnDpqbLlbTSxjNZennTPLLbcppWLaGbkQtDgFvHiOVfKc72qfAVgexcSvvBXR
1mpmeOEM+L0Wcex6a692IQILlsovQIm+sP6KIFJuUYA5BS4/YKJGElafTo0QolnY
i3aQVjSKhcuTguvT8ynXx3UtWbBEgb8TrEbaaXWEH8enkeTIsQ7D0+xeuVx/JaJt
rDmbJFYr5v6ctzRDhqKuyw8Jh9nY+M5WEMYq1yqmzlRBecQrtYSMXqGx/323mGlN
EtoGDsU30byOwRgcbMQQYho0hvHRGfajIyD9FAu39Xor0IwW4gwSfwlNLRLWc22j
naFwhROysiUojqDz1n0a2etnIeHfOSnKkEWuvmUqWVf0ASG2EaJ+yevYIDwIyAST
jfyVa4dkzmHvDcsLpS8ezP7pMrXhFtThDUPtxOFdmMiDnkHc3msqTZcAaPVE1Qlx
O5ybSHo+o8WHxYc4VVQLSgYSuuRjyhTlLoCwXi/y5P9LKDzjQ42AVWXHyjEQUZnL
mDYGx2FVVFwHErLbFdu9GO+gJyoCLce1Py6G7gENqDyR1Uclms1uaKleQPMOjAb8
FBSo9KSRpAQXw+m/zKvwm/ZaMU+6FVuwJUqdCE78EBDQGW+zWkw5uKuYlgevdiVg
w1a0xmHBTwlNHDB35W6QAfZmyZPhOQUNtMgQzMkCTUk8RACxSqTP34mWMtyclB+B
z2+0GZJsbGsOGPUKlirif7sJow8tX9wdu7dE+neUSKlA8XwTJo4mFQrxcfsOJ5R4
7XEAKOOfiUCW+q/IxmyyP4/fkFFWdZBSdfeicEJyAxHhqnMbTsd7G68JXtVgiQhE
+s3AgvbiLG199LyVYihTxemZrIi+Oq87ZzfygBP2TvKpA9NeLHjlSIy8qEBJnABw
FFU/Uf7zsm8BcEflsaILHSLAUcYaccWOkgHmvEX0o+r/u4Sx3Zf0HPmsnFt8WXXr
E1oCroCnkrUmyFjOp/gPDjfIIDkveIey+Lp04LhUCxGZOYSsrDh8nlXa0gpnbU9G
uV6lc3g2Y4C9XaU5//+3wMBMfhjGUiP9m7i1J6EYT6+VkkAhRjKI/nncveyAZUgA
Gs3q8qxvc6+3l/I5WJK9GLMk/cjFG2hWV5+ddkHNy8JDtbVr2hEnqg6rqWK1Yxng
x7p5qF2Vv5lHf7GarMo43Xno0rIIrC6i8khGF2ak7w4l0Q94FJTd5/Gzod69HH62
Jen4YeZdCFQCE8+pADpQLvGQ5Lq0er457P9NZeHqf0F7FOpe3eHyV+zIG18De1Ph
QTibhJBhE/LF+7IsnHYn2llMTHAOa4lFxgN/jY3HTp/ficgHvNCYEvTFSY3+cTSy
qGgxlyC27CvRXlQSRGtYEljCb7me9LOdSU+PHA+PzR1omnjI74e1ZoWWOp08cQVi
is1VPBx198btmvGqf63fQRcQdruw1BVj8GeSmcXCmJA25559uM9QqoRaz3tKEgUc
NxwhUyD2D6GhWiC59KcTDKcB9qlnZn2OFwVXAACj4NOX2je0a69w/g3KxOAnFjlx
yKYeUcWLZWvvr3Gx6yi1cuz2S5MYU7H7xIFQnWOX4T6si0ALxiL+WKw+RtQES7mT
+qQ5G9mwfjEMEYF89ElBcVDX6oxr2BXQ++u1a07OgYWAmmVobioMp0rGjMQon2TC
9jh//6qNDWJNcfApx5bCxcP7/j8Vch3XP4G69GlsZi/L+eSqTeiIlJbQvD5yRQAn
XL0pCANapOlBXlo8OlUnmJ1zjG4lcSzM2S2u8OLFcK1Uznq+1J/NmoJaFst5qaqZ
OfeEdF0LcLTqBSqBbvRgZ+CveYeOEIk2GvUOYoh03JRkYmKW8CmYPpz6UwjlQ4O1
bGDa0LpEvc11JGTMJ7cXQQpClbMLE+gkvfwzJk6bfW7XyqzgN4bUjIe4UtRRu8qb
zFi/fh74qQpHFqs57MC0ygMZqTKTp2iGQDVvp9FBZUQA1ZcMdt92jNEIYxPkCDLq
D0pOYfbn0i4cNyv/n9Bn+TRC24M3S65wQj9dG2rSOvyr12myJYbRiHNUTAGuhxRK
dH3hfhl74qYdPU14C0dhZRZq8y8z/dxdYL1Igsx5EtzDdI9SaTbf0HZL5YVFS1e8
zXLvBIMoaETv4etfr5dfMygwiX+HKEKNSHZxb7Iwfi23jTgttxhuoE0CJJZeHrr1
ynv1m2MkPcLTy1FtxiYbDA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rWVsVkQJem+qIxn0uk7jDi8VV1dSyqFD5PLbiQ6Rd8WTI3Gvu29X13RkVA7wT68r
08GmVHNMdt1Y4SRJb59OVsxBIXf2/czczMvHdUJbeDy0Y7ACpjeQk2U2Lp0X+atn
TnK/C9PPwyvRWkCVEjjTnN5ta1QDUY5XhXMJM1tQ1wSqmGFamAjT8MAgX1BfAsSw
B3+8cZYl9Z8ecqPSgTl41IIvOfrSIqtoOfeujfAdQQeWadZ2j9w7tLJbwi8O/XHB
iB43EdkH+UFJ2Li14EhBlWBZABN1Q+79gNNEmuKjNbR6wnZG3Yk1pQyi/g8c7Q7A
z3ezS4u7Pi8aR18iOn/1hmyXTInObjRTt82TgNxZ2Gfd8j+xT04J6+mKnMFMm1+K
jo/h5lzZkY1dvdAt6I6kr/jb3YGp8DZ52Rlk7c95+mERaZVVvv5UuaoB6RQIv1ES
bg1PAVL3ORJ3EjYVQpMdhB8SyFnzb2AyRbvEMeqF8ADPttQAmj6DlU89586IgB3/
Ft7G5fqFcXdQgAvpRP5sQCf+QtfcwORYC8Qg7M244FRsL21R7RTtl8EBhUqy9X6Z
QMDnVWUDqlTsHwQhXs6zYfQwXx1moI0mMqARjosTjg2CkEtdFaXY50gJxFdK53aE
H3aZtY19sawunst41a1K7g==
`protect END_PROTECTED

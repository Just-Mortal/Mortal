`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cSd8Vk0TA+sAOO/v7wsUEDVkuVQmFUJl8JTPTE8herxPkwixryQAVSH7GlO5xLzM
Z9XzBEjDN8+J61BqGw67yPw8FQh0agQhI0ISp3ziShhbbd0w8N7LcT+Vq03JXwOp
qu9CtVsmmJYbVa0vonEGKz47lLyN9NOFEuIoE3b6aul3OiOPcENdl5H1/Xwh3Cba
FdNeJEg/oWt8g+4eK8V3wvk3XjAnJ5kwRwrZl1/EYLi6VprQ+WF+rL0UVmOXaCPQ
khQJxeFXJPrNvXNmdFKD7NLhH9RqbuU6CxGvkUwmvrYqSKvCaLYpHPjiSyDz3bG4
k0ogvgHVjwo9NjLKRjVrY795lHxMYd8vrM9Gx6QYQLd5xiGXnz20qKm1tMm8XVOR
wr6LM0TY2Sywanvf7qlqKHfGrxwlLOZHPwUj4PfY+jCzMg8fV7zVF8x++EUPgTtO
OK3WDnGTt0j/Ax4GAAvmOvl0HPAeyr5VupYsoKefpZEHO6W3cHoqC45EKkEpYd+N
OySNBKesQ1fMRZVmoz9lOXbQb4xX5jRnsPE64evHYj0NlTH488YRnvDwpy2Tfbl4
x7eAAquUXSmlYl3G0QzmJFC+TiVtG9dyH8YWPbDNxIOiSbTmrs2p+oAA52W0Sabn
36yomQrRowLcZzJe75feOjazhaVxQ6gXdRyEx6haD6Ew4vpUrmDegv50hT5KSPuy
av4YP6evHWQy8QovXiMjd2x8/NA2gAE6z7suJUS34UswDA8DJDQTOqPMzr/vHCuf
vz9woCO5i9TqUnPc5auFHp65jDi9oNxpiLfDQkNFSLo=
`protect END_PROTECTED

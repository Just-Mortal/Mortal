`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FJ/x3zT4kC/cEGChNE4c96gZ53hoGFiyDJyoaCYoROgTUBq1ZRPVQRW5VL9WF1XQ
86mxKJl0EGbTU1+UPD+luRHcwjYhdDhrkRWJCUZQ3YxCQ+0oZyQltTbxCKtOJs/6
MxlrDHRBinSroTQDG0BJRDbiwtp5Cq1G4Yswxr246KV3LhfY3yHR7CVSO3gdJGJw
3FT8/ACGi2cS+3vdubBhTqxPGADdH3m/uLAvSqLYTy/Fb0vEc+EE9tpG88JquHzN
5BW7qt+epJ9lTtK+4A96VEe1wxIV43Hakl0IaFUNpkGC1kMh1AVgDpBLyknmR/z+
lcfnHcSecMDAeWW+opyoYU/NUjJsEA4G/xLLlVGLxnbJanD5QdT0H9ps59IOZsN6
jDWDg1uzW4KAx1HV+jpNtxLIDWmxYS+5YpgSOeQYRHFsGc0Wf1S5LfpE8AEDjCv0
tBaKSSRtiZAcWGyjaqKf81cJGouvPi34II4UEGC/+0UnaywtWhRDYjb0JE9oDJ6H
HlZjyFyq97emzpUR7pHRlB2ENZs5+9l6uCA01rktzGT+g9NodnpICxyMslk9fKPR
Ng8zgpGkJXQQNzuPa8jT3xI1yl5ngF5wzPGr5Psn1qLroC0BUeHRZ0rouxKdxOLE
w4aqYTGH8YooeaVGZ6KIORlcPVBPCvAqTBrFUQPv+ZyqfsftEPWl4t2DP92NjrTN
+HKBI9Poz6KGEUGabX1hz2O3atqp+JdaNYEyRgDA4VMw/MlIRXwsYTqcfepmegD3
79jTX1wUG4mNgVJ01C5yLO4jLfREBc5943bBRmcpc9w9zO1NczvgP+1N5Y2kh7Ag
XEth3SAk8kMOVEdAG3TtXul0mL9MDLRTZZUauAeTgwCNohp48Rax1MGeRO7mAwoI
HyJPHQXGM1Bcn7DND1jTQpEHgV0rP13YEuC9+mD7M9f75UHA0DiOqpSEXRIxHQB4
wYnm8IiSDrVA3Z2y3iJwCeStHur7rCp7dRl+D2klZYfNXo96HQHkoO57TV1Q1ALP
wJMeWWtq/DCHpLtLR1/rXNna20WpJlk4zdP75Jpmwtm79MScAhW9hupTUaDxy1xd
r8BY/ClaZkN8qaumO5vv9dKK/1//G7WbTkwbE1Ae5ShH1EoODiXOJpJg3e90s+3z
ZAIn7/ublI4uhTONoO8r9RkEGusDl2G0x+nUMxWxD7HZkPNURWoxt18HJRjcATnM
t4kP0Lz9m+6kF0J36TpjXRYsz5+EVmDwRHgg6+vGJJ17Fu2UxpUAjBcZuA2IpWvL
wRNHH8WMXP6yUSPojAJ6TZZPsCantZOPMO+N6OJNSypN2XHeSlCRZi9LmaTG77LK
AAvP7pxaKSig9AhvVGnREte4y81NKbmWXtVAa9HxZJ0T6xVW6mTPmlcbcYRbMGus
FPrzgEQKdIrYpwqxY5K95HXe95C13nxUGopTwBL4F73/B47f+p7TrDpOuw7bFUyD
h29QCViwiKyCBLJLWU900+sQPlNnxctTRwen/1juSyUwrpq1/INpAHbQpas/B5gG
mRZ6W7KrpIj5FojNrFGf6jQjOVzLEtKK2K1Rk21qv5JKG/2lkw+65ykcbus/3sTR
osjj4VRz9D2X8XkDV4GmSU0qC87OmiVpwQ7L1vy5xv7PGueWPzefqubpOPHBhpZ8
anUBTUnndOUwuQ0ZRR8QdkL/SXcWsuRtj7vh+ROIHONrSW0DBvbo4NZGN0eaHTeB
rzyrd5m3ZA5B3Cc4O1hFdOWVt5ehzhutJNo37eYuSUFjtm5O+G5SGk/bI3b1jii2
rmQeixaplRK1tUnCuoVpwJbRlBNGTwYIQhcMgJ+WojfPNx+kwSjiOvqJD6ng1Pxl
AHCBaEK3KoZe9set/T158yYN7yHNKrNYshs/Uyz30GNSPsu5DtwGha6pzhQBBOQP
HpU7mNwbeHNXrD/UnZNWMDRjmOOg36n0DbGfPIzNPX/jIo8jt+nQUFK1qvo5i6pW
rLVYrpf3PfXqsxISbUd+U5IoW8P5svpM30iEieM7AraEqZZv0dBKDwb984HdIq/e
eJMtoe8VQ3AsGLZCDZHqfwH4L1LY6FXO3JxYLrYd3FyN6LsrysmiyIpcx9nxbYvj
UPti7DbVmL4xQBb243Irh+ZGn7qM1K/A/Dw24CM1xY9Srg2bzT7LlCClRdn7M0un
Ovc2cjydFReWhxGzQfOCP9TQR84DNldFPBlAiGXC/5j2l5n99UH4oc3rluMU1kz8
25YZSJ39n96sUrKLKwuPHctrCfVrREzGHsrbs2jxwJ+E/7P9YRHziWRYeafM0uTg
Z1lYOwROPtVP0cu1tJPtGLvjgEmmBtJubL1EC+EGi21jgwEIskJOYnNuvrGdK6aS
93HU4+2p6N7tazqNM7Sm85pJeEZW0WeZ7MQkOh+vsdlKbpXodnI4uQLXWMbtL0nO
apJh2td79BVe4s2zjkZJgzPZZ4WkwMVg1vHzpTxcApGxDGU2oCnclSzB9K0gmrUF
JNziE7Va8J0NEAlBGZx8sSS3IM1tOog6OJhOJ6GurDXcnLmOGwzsJscTvPuHM6T7
sCq+VLF7UQr2Tu+aXgTYr82AHRuQUhTXfZUwjaEa06RgVgHtxb+VmAjDgNaRu8gY
GJxmEemLWEn2sW3qeofJMeG8OkPjLgj2epZv7KjkbBY3Ida2A2343KdQ3rLAEt39
4StnUNdIN6ud6uN4rjanobMbaYERpSBQAdZmU1i+JnbBeBOlvwH6Ti9G33DtFYpB
58qOCatbiAeMiWN9VgtEZAD2ifop+w7+lwFSac6VuOf+ZtpgqeNq+bfRcW1krAxf
vzpXOLNqa4264ovB22BMFGgoq6VHnZqONzf7ckH2N9IssJGAhrVxZ5Ku+IHOZzP3
bqhTw0nHhw/29ghZwxkeK2CiwxGZ95kBj0uxCV/Pc73NMVmr4BW/saIcX962o1Kd
22pGkCT+KJbk/ShRBezC6+qJIg+iIi4S0o/ghwbKGFxFVZvuaOExpaZAVi/4RTUN
4JjoWW6GS0oTOyl6NbFRD6vSrgo111+cTN9+pYk39i7aLkr+Wln+15hE3GYmNYoo
QflZRvo5VTQJYXJunEqm4HKlXi8TIe4dwHxMAN7/ioguuwhJe35u7oIuFPO4C4EG
J94/mu7nz272ckgdOmVaoWsaVShRvSudpte19kok8otrAg50m79a1uM8OMjnhs+0
FVN2Q3gPuIxQjjXoR0MLXw94tOPpo5xk8oxtjqnPQVemasSjUa/LfrL+QWxVpMlJ
qpf/eKj8amYw0iv3GCcNFA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VGta7Nb+onGLV8f79sdaUmtZm3INm6rzV43uMGipTG98RrJ4MtYJM6Plrmol4Lry
KZfz8lzwLTvyisBJcO0nxX/XnwJh8UIDzQbs+bGUOmwIon5mJ4ZvhUbgI64cCgnW
gbdxgOswwt7FEoxoY8VbxvcP/rCMDObsDVeLHq0h45lSYQYOxLK4UKEnk1j0+yRk
atIxImngi9RlcpSDAtAWFFn/+76MzOSrJiTE/7ZHMeboTKmPzETjrAe3VcTa+LVL
M+gNcn5bfnrxoYdqhAFDE16CpsRbOj45kMK4E3MgVtZlBA1w0hPHypMehY0PAvbe
RNrCydhSlfg2jDukcr7C0SLnqkUG0zRbIMLg5Y0y9VR4P9EL+yg1khFN9am+kGr1
tQHB3POjqj62ZzSccHFavAhDpHS9EMdF5e+0bCgub8yoOq1SwFLRpn6kZDU8kLbn
ANrgmdQj4msZC+JeWv0VEpKaabkTtk+CBUZJbJxE9Ydjp5M7TLB62HpVtE2bQvT0
KL4+3Yl1LZhnTKms/oTVtKb7YNodMR74COE1WRTZVP+Wy3Sm9ohyCVXDPVGkwHHW
7xyZ/fx0sYbwNDY4nR15RjtqHVFP6sSr8Ac8iWXJ2PK3at4esHVfkEpiyvQiCgVm
ai/M2dzDFcRGaP7AJ5FYQ5wuXyJJP/YWGyaWBn8BQN2ZncU35vEXVK2RRrjfCfTY
HqfO4woAT28u4NwZsRHmG0D75uvqx/SjKdjnpsGnAXznCjPVtnwq/Tmk7CCmJH8C
fNlxLvsD2dcPFAixn6w35nBAkfAfu84pcDUezdj5vVPDuFBObxFEHu5MMh+hFsId
rzBVNd+uieEqC6ap/QohgaOncw4K3ZYvyMoDcOPXMYDhOjY8GTG3HvwYW6hzzkwN
owC+EcbSuAfFMMeqnbCJQ9V5El3vOBwk0fjQt3BZuIItjfpIGAGmaPWGCBHairQb
ywISeKM8NXJLVwyUYuzWd7QV9qZWAdX6cNeOpKZZlFEGO3xSNWyrS3+M125kEVwa
8XCTejZXr+53ylrVxuMyBUItRn5VuRq36rMaErUwoFIla64ZjxX5OaFcNh/l5FGf
djuiEs1a4ZOJHw7tIHKBvGouXgRpUcRn86gIWcudxxp/XTv57+bvinU4XA4iTGZ4
n9aouBi1vmkzH0bvc/rn1hA49ijOuh/gCpqFrW1fxR671qgtzDBnoYWtFAQQvkue
2ZK5ihjdnldboQCKhr6RrmDdNb3A2ZqIjePoVITS6/ZnetNMS0J2z8bjm4h1YwF6
GbduiJ2U+pAmxhVkya+tnQfIkjOkP+FZnO8Mdm/G34U+rop4GIdCYAYQhQszJDLS
4Y8JoM6u0AUsRoIPSb0lROCSl+/UCyoV3N+bwDnGsYRof3xL8huyw/MbEheM3JPZ
DI2/iLZ0YlDVkoVKZ0S2cwcLhBdj5UQAmqAWxZYHFvZMf8gL+ctoI1b6P5mt2iq0
Rrd/5/fQdja/xIa2YKh3dDAPtInQVDDq0gAcqh1ypgZj1bMPWABoFlUO2gVr/jN+
YyIGhmEI4zWshUPE5Mwy7Vc8Xu//Y4/qOOsbnIfVnOsLO+3A1E9HrlaDQeh4Uyfk
hwdohXfj4/nTBWempTmtjn41/xp1urUjcUzKsf7KLTuJiWjmT7QNYNciZGNiVvOZ
SwDtGwdFfaQ+BmRuU39fhyHZDs+7Nhhvnfvz+iyq2uSviwiVs4W+QsM2dCerTY7z
mY1u/BpGrhljm71KXstXSRWDfPnGAC46xSY6JZIXZv/CafSQpm9jccL187a8hgRi
7Xf2j8w52M91dGvOEwHg7tmjTBxrB40h12d8GT0qbXqywFshxwlZVV6IsLKWOzl1
t1xah3Ch6aJvKnB3jG1eNK3YiGKJVNIlINTrkfbUEvXfwNCotf10ARcE7uw+QzuZ
vgLV8hjUwy+qvqsrWzdw5J73TMH7HMqrjKtNuSLrWcnjJ7eoUtnamrMZtEikBKP2
jChlIdlcSsIeJdgewKnVLKt0ItjaY1X8F2+SxmxyGod7ckHnpnkFaQVU9va9HxGk
KMq9HAJZ4a5pl4/fVdHiAngQnB6t93WWxZnao7Zev41Lk8ts8U7bMQLIlcCcCrBL
EOivGRTYvu/qq55YDWN/daEcEeGLFhCrMHninzyDcwBQOX/9vk4MFVMdsdWiL0js
TGi/E5RcOCmykJRWD6iGeSoeSHf3PB5OjhjXWvn00HbAvE9U/vHiITmgLtxiPewO
nH90CA2STYgDtnONeLRRahCWo03HyF0aQ3nLpmELJsxwJvEgRyPp9VnRfgqk56lW
ZNuPKsOcfnlVN3QfA8Zj+y08ZzG21dxyEvTHYyGn9YxR66eIpRPotwH8LvosYg+D
T2+eFPmdrzIy1l9xnDExdFEjcHB+/9DvWNYYeYv7Y0JT9Ncf07peLoZrgOg353vt
xSfIBckqZhXOCMc24bx6cIyODvWtzKrjt2+QCTZwvW5Fu+NG9Mw0FsSiD0syeK6b
QLT6U1hwDkp8UbSOYe8xrz1Ga7Sk8K/XWSuRfZAfsmK86V9tLRUYBREFFuoq36St
hvniJqRiNakYKv7PE/sm9uylPb2L6TtKMbitjl3aLbbQMliLhbplXV3Zg516f7Q1
a66R7ujCvAsQY5LCgDRiZcvCXPCMFZxQdooWepmISABuBhkpjpqUqDEdiJKBjqYJ
BA9P47bcwL/SipbDLlcfZVhFTGegaS4cqfTPqbGLt7VkX5lDfTCqnsxB4rW36XkJ
YXi2Vb27mtk3E6CVZUkdPyLy4DYesvuCLPV28Lt63q9MrERABN9rwcXxpMAdK/+V
iLYWUjlME2vTfe4GexUKHvixLYuuMz3SNRhbOH4j9Z2+RUHkQLU/uM+XucNTt6y4
rGp4mvZopauWuP0pxW9KBuQT8f4nb5h5oQ4mT+OXXqSu5xy78mWJOT20x6bfohys
z4ZmBxSPVUvJLJnt8H/Tw2CxGek6VUn2NuJsG8ldVlCu8BwB26VbYxO7X99DwDk+
Hw5kfxmk8mWUYrUwBEjThKQ+O/4PbJy/Fy8DOKCEXCIy6/0AmnrMugZlFep5rfLf
Au7bQQ1K61xGdgk/eRr8L59UxMW4doGstoaz+CDKkVECkYvcxjNRWL0ICD4cDhwA
8IiV80YOzQgg/QtVdGmYC2NgivKFahOoHmyLuJCcw8jMAtd7VbUh5hjHP69vYtga
h4JgmdV/n61s9KVXIAQ9NtG/0iClTyiSVux6LzJVczYC+egwakhwhDaEtrkf/CZQ
vnMic8G2htEA0Kd7SC7MIb+Z6zi9I//z/umIYOpSQWZD7GRJ17ZuCMdjDHAXNuO/
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4mNNEmc2XJZHjlf1J/wk2KasriC2fL/RgZP2eVHA88d0wEQ6gcaJMpDrgNbxL1V
4zfaEx3J0ltm5oBClAy6fcqTx09x6CemvFv/YnUixcM6uLhxzzrbduVln0oQDlMk
oKksnzbHNRVKRZPr6Hfl0eMqGb00gl6ZBfTSqXalCJ4QOwEfDCVmCu3a4laIXlFE
D/EzsRWh0Li7HY6yeIgMEzqn7PEQeYB2WXAAR1gGm05cFauNTjKnuPpfLJt8zLai
kE/LafuniUojpsuu3NGLIO4kRpHeIfTramwUnsAsAd6IUQtN0rK734UtDtn9F4T5
ajyRjlyy5TU4QyHteYkG1xIJeZdgkypVF8So5hDKBZprJYEY6MXTKjMqJ4CYo7w1
3DI/tlmuKFaGulDZSJbJ8xoexpXiUXVBEiANDL+O37Ykhwev4/N3la8GCHD30gnX
7gY5OkBXRJDOFWkc/5Zgaxwyc5JuZ7I9yd1OrYxGQch1ehEbi5pI+ysUV2L74Wbf
GxkrqYvMHZrJyBt1Zc/t0g52reXaRMuW/SdWiTN2giddPTq3xJ0bvRG2o82iMWwI
rHkHSF80lcyWYmx2eR6DuEjGx7UFH25u8o5bgAxkoWU6V7Yrmpg3j6O79y+kBSTo
bPr3dvKOMAtdvDXAxvUDl7cqTUIL5WphLAUv/M9q2ZPj2c5VTWWC4vElGygWG2+b
W2t8oh5i7ZB+zThFzMVrRfHyT0eywmgE/VX3AAIG4bgZDdZHf9Vx8OyKlWXGgfHb
dZx5LLv6iwWm/NwFnMGVxE28IJYmEk5kub/YEdeU+r9ZOBbo1l3kZhmUcWTJPv/f
FO1SGp2GRMfHynKfBt3KfjVNsQUvus5egKt4wQGN0AXmS+e1oBXmP4BJ9Mjo92Ce
CIDLQMV07UaAHwOheaZcD8sf1f41GveXDWAI1tylpZ//ydaD3Dogto+KE45l3JAo
s+afgwwrc2DPKJpv4Hzc2X7KVek+okBgMlB3+ND+01bNSkF6hAZ5mJ4PD2ILE1Qz
zUdJ774oyA7wOIvIV2MohbSkucxIJtgeCzLaNeE6UEdX2TVNNj1KEWjtYceH7MFz
csfez+2Ub9BSH0OQ6pb5SFunTHU9FCGc0t+3+16DQrGMKTIRdlkJwsh3Bb/1hLLZ
wdEeVQ+akmtbxunyIzHa/i7h8ymB5SScwdgM+jvit4koYo+Z87AJl9wVbNTyY+sr
v/+lF7TD7ceTKUHvwiAfBf+cXBo6E3pWLCiBiCdTEBfgwC+j6zxFvJ1WDb9XiDUT
l6M9ZqZTev988TCmwxDMucE3GCw9ak1mlFzvGOGHlFgAGpaK84RM1/JarwlZKqBK
Bzh+vZvBEcSeY6dquD2BNZipVHmWW+CxFhccZJXjzYqIzlezctj/nPzO/yyf+Wuv
U5x0fUV0WGr3hd3Qdyhyxm7RqA472s1jLyTftVf6U8RYljLTIYzSw51p6Ou5cSPW
xdo/5iy3uy53cZeE2Jg1iemdRQdATQI+Q3X9TYilCgOStmDSUNzcD1BXSg8J6oU9
2E1cBpYQNFnpscxM3OOBhIMlDVZJSnuJFcFfZhviZauphyAVDZjhaAHu1iGVAqZV
D+ruqToDnGXDxz0gArExmna2mV9HD8o7tQwYlgvUpjZY9L8e/eLKz5nw+oOSPt8N
I3HTUhUaKVcoFLvHk+2egzqzexg1MO7oybhpKnIH8r/UZMB54tzEutqeQhCHft4j
rf2bsVcANHw0HyGyHAqn5vmhA+lleUrmvpsxqyHXRUFhySbJccIKd8bqV5B3T122
jzz2LiuvJSPH5OMtxQjwu5tuIvJrj21eMoLhx7fKVMY4jInHRtcjiJO8LnWbRh3E
Se6Y0vZARccKW2RU9CR1PykAzvgj2Pntns5cLwjlmM73Z3KDYznaOyLx0LVmW73z
WNAeSeIyfwOmkkNBtj5xSGSlIDnn77OF0XniUiSpVzml6uxwbcj4NcqKDSjcmotB
ZlgOFZofCNF1OtMIhi8Xe23u5vZDev/yIqqFkwZflI9DEO4ZXxE3SSvFPZ/rMuUn
TUI51gx6HUcFWFsXKpvWdhMqYcYXqSDP5Dk2FpqMn2i0a0jHF16IWh0qsNMCAqEN
I6QAV5eRzHm5jUZ7DwrwpUq+KSUHraX7e0AM0O/U/8T4+DVUcQ8KhS1DlbEromY/
oX3Wq1c5fJ2eDBqb9i0872jQX85QjYIwu5SUrlW42DOyazJ8VU08d+ft/16eYlkq
0tLFGmdnUmf0FA5sez7D1IqLlGwv8fG3BUIjiJ0zbKg6agGSZJgIRS/LRjyC3Fvx
c1FlhdH13CWoG85vWz/yAhmfChAfdW6lrmL7PhdqFKVZ8p0f25/CqnwOGvTgU9Hb
WNrQy1JudSOJ6PUI7wvODhCABRZqxZ5kOIj1nPR/vMhUGZfaUJkN4H4z4NJ/jkfd
ByzUHPhHzepm9Q+bCpxhJi45qCC/dhzAcEQzI+fFwnHb3vk55zyA/WMrZgdD3LcA
CHo63n1oI6PzE2BaGJbm2AYujYlRVWZXRpw652WC5VS6dexpSEVNREdv8T6R07Wi
sq05Q318Bujw7pUJrYkQShnkvyNVB42RcbYVzqHHVQKB5icyr3FN5em1t3Hkdvst
ftIjchChqfqRnB0s6wWECXagFJErmj9xApbldP3gRKU=
`protect END_PROTECTED

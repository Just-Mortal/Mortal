`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qag7u4Mzj6Yz+zId/Oyv9j2VReT93t2tH2bbRGi923UgBBYwLBvo18RLdrrw6T2M
nc8oiMre+wuRe8Bu/KgzQxFNt4V1upg7IId9ATRTOITq3GPbVeR3+Yu036gVtFgs
jQlBuTnxKmiJdznsqgGXQaGzqOD6N3zbpj3d6iGFch9aI2zJElEUlHH32FAW7NSV
1Y0IkRD3rIQk9pwu1Vb+Qm/NE6M1qMQcYOGXfcj8mHpkbC13IxeePqmhCTPNSnAk
PX7prCLb4Wmtt2lQ9oO+Fsl2fS55rmfqUfnPIO+vb2IGP5AtsIF3Xe+YeNvRrmBg
6h7ynDdKXtRvukflawPMfoTIqAYNV8G/OB3ya+Sj6rNs3dICjYqnse+Apk7rTueu
QaTTiJVrWKLif2eBLf+69+t7IDeSsb38TfmkvCMd0luzHrMcLWTiXOtYxztmehrE
9EdnmBD5ZVjjLqHGWlmNPFnynMiaf+HiBOe+zxSPM2/iKpPOgHyW5rv8DFqKg4ri
5WCyPVPQJ+TGSBxPpCpDLu9MXSXT6i5TZKJInnk08+JySjFiCUzhXvplkW2xmllZ
72f209i6wG6FEw5h06onOPQoB6CRRP9gA9n9L7EKbgX/5r4bnETlvd3J5Mzn+OWJ
yKLokBtt6kfaOQ/M8PL1QL4MQusz6kpKajsco+hTYBv0Mpv0aKRcPSIE5qVbMSZ3
ey1dpjfkd046mJ9GQ5VFuKnaEnPfVxRJwLzp+60GJ9AD9dPv+t/9ItaFhIjTXL2p
AjKd+Z0gvN5bpY/zZrqTTsY0+MEIVL1++EtH1Vi7V75VgDmz8E+YEFBSRYps+HYk
EuFk4hyiZnzWjRLfkaK9K07C+qYpcNiXg7UpJztY0xhvsY9fXWVtcmczP2TAe/ya
eIpgn3wvRzXVcQcShXTFArkQeEQPgvet9BTo/fZt62dvhOxrBSooMPEhpRdQdvwq
arE3hE5C77SAdu+SHBDHPi5IsMDHQPNre7deXPNe8GKhrsJeiKjNnkRnN+B5ytua
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bJlPmsYd3kpvFNzZQ1rIWVMi8jn5gS9FCvg+9jDpPHrYAaGhqiDW5D3OJImwyfF
Gw50na9H3QpAIZyZuJN0hqT3/nta9Vn5pVSNAYMUBzzrVZrN//9f9mqSVVHqWyUh
eeE35xp73lRn/iL54c/f7lOTVTMA03zktZjhD1BrVXxs+GCCvTLBAuhA+Cz89HMk
VaGae4CEQTTFZ1o41HwyozLIgxmfCtkStrknm0km4Jle54ril9Veb60HQxK7XOzC
cJAX17cVi86vzVjJA3EQCCvVpDmsqUFjzJP8CYQhzYVc4W6dldHI7qfofZy4Eqfb
ch1QRgOYrp+3GX9L8/TR4XmgEBLt7DnpfYQW2NHUpxR+BWNgXxsF4hqSlRS4cfZO
1ZypSyYF5nLaEGdevUYkqPTh8Rq0La+RmvKEsP92rPQoZzaX4SL5PeljvwUQauUj
4JCouOKg+Lf4M17FBBIuZtG07Zf8g14QQdKtdzhZvSJOLCTsq2u/BcIJgKZJ8Am6
IHNyrsFmJa04mdN7qy7UvP1KK87VGKmCzp23H6f3KckPbUB303ggSDXLATQYqm/n
VRgdiMc9vchIKI9ZaHLNyoX0xjKtkSd/z2io9PpQSQsRKXJDyAAqFRKZa6RWiUEK
XHSijhdguT3l2P1N3RPRL+M8LrqL5mhVW9Sz9oCZoRG6Nh6zJfeUgFg+Nz7QKiEz
boovZSdC9CI0Y5D0M2xPtP2OCRkttm+QZf6x+4DW2ObjoCCwMMyVRFKeVOu9oUp0
fvhsDCd5zYdkkqFnEGTq5CSxQhbv691kWxgpmDFHIORM6Uy1JakSx/xgYlfAyUoK
Z78Yphvqqfg0KFHw2/2BnYwCQ7w6AEcpl9zSPZP8YB8mevmkpoYBy+WLd50pIkEd
yiXs6JePLwRoDNXF0ug5SF5UOJF1pKHIog8bse0moq6yDXVWEGMgQZf7QcjoE+mH
aYxa9u+b4nz4ggni7fkDHoW+EMWWqSS+IYtduA6mFE/t76InU7Juo8MfWxWuDnXa
yyHMkY4zSjOinJriyQ3dF47n0FcYzRCAnRu2ORUOkHuC6GOw/TVQSalFRhLZHJwO
xf4oGfnPO2xaHjTqJYFGElFdVHx5XXLPHfcbwz0r8KZCEh3EWtQ3MvwHCSyDXpqw
+FN91gtp9gpN9iFkxLYBRWyaaofulQru9mI9anbCfZf0pz9dhYCyNdrW7W2vFA7F
N9YSavxpQQHlzSmi/ixAvirkadO3RKb8ube2ig89CVQLBrg2hLUDWK06Rp3wooxi
gsxhbjrbJji/pkHx8ntUSrwsOCOlO7KNdvJtetdKU5syj7rbc0smKcyP2x+LUkvs
hhyW4E2D9MjXVPy2m48uh/5McuACoKUnBk0ll9IDLV+mKORcKK5DR+8gCbctdjFL
AfHQmclXC10WgW3mxCRKS6SQ0k2XMv5jecQSZDvGAOqWbHYIbtFk/ZmS3FhMkqw+
DmJmTFDRGc8Zbux7uzYFtB35AmVUr6ElK6V7WfCrsToz2iy0BQ8sgqrhJdbxpoad
x7OvfmPbBiHKyXbbCAqZk1lJa2baeoYsCS3rjI5axoRpYr3EosaeZiAVwQYCtabr
J9q0xomZIT0vvGl0lUQxBSo7pxo7UTOVxkB8guIf2MCtBOSagS097ljkRTqGi2Tf
yAXckdH/FSDfPQWnEEhEYuQgKNxDILB6SEg7nLbHJ/H0NVulKL8VVYdIA8UlhE9M
PGyES1ElCJlDyzOaBPkLInnGsqA8BPsQW/3FjuAJ+0wb6bLgRenbjMy9WuVbKtNk
fcZn3zoftRioiRYx+HAF4NFdP7o507MHK1B2oBI0KS3V+eqbWINwe5tTSdHzjBVR
ylIv91DeRzkER77OnZ1jHKQeR7lkb4ea8BcbokMkFH0fhM6Rp+bNZcXpjGVfmd85
vm3QQYGXzE1+3f3M/C8nBW/rxf1zS2iNsJNuSmSnIHgX/EX2m3hbh3HpvBGQbL8P
2SH8Uykalez1+AGiHYjx9/FwDcF5Y8sBJ0kQp/QvABjFf2KISe3s4BzDBYkDAWvM
desWm/I7Rb6AuxuwD/+S2V785GHtPxo6CaL2zahmNB1exyk2T3kwX2hi9DB3WR+8
sstnTgkjPqH3rJE0GXcEGvLIHuDJd5C5647Z1bitpOZWrMvnitWRv51i991bO7EL
3xIFJS3LkneeNMvQW/8VKzTPz4fGfTEnFw7Q4+nAlAKb4hiaYPTPjcY0NH54YNQj
d/X1Yxo36fOAanMSv4ZNhco+W9YY2Rk0sBC2bxvRlktOb66cAtu5ofAyJ8Zue2sH
hMRMcV32tR/q3tYEggGra2ub5SGuxHZdN0fNGYUpekBGjNijpFSN0goTnQXqmkB8
OHI0M7TS3jZDMf98PkFM3CaXzFcEFLtXGtZRYykn8MgxAzrXYRArvwzTosmc3Fbl
thFw3nlBYVdvL7/q2yC5TfgqJAZAcorVVognSFP+2RitBCODzGzVngmGUgNr8cvM
vDWMpxEFhP/MnK+OlkJOAvxdmeqzSX5p6YnNzMjejit64wQwTru6bjJft8GERviO
/mNa0oUcw12fVIgaYLNptW0j/94anZ9QpHxYt4/t7xecnX9b9sMjOxIIECIUKcA5
kVmq6hdiO+TsrvBlRdX6CS3mrZWsrzEHcaWZJsvP8vj/Nwgu8wHYYnr7P6XQ+2HJ
qaqQw0l/WByx2Pesi7Jbdcro6XrU/xET6KygTgrZK6o/t4WRVMZXbZJYJHe0C2Kw
iA5vBUU4Ef5XvwZ4+vwNh51FbT8IEMH2QQ8qYtCFRQL+B5wzezaCbECMc5aLSvZX
P3xCk7VBWOyttK9AYzbC1hLqhy6G0VmEbQPqmr3e+abx6I03k0pd7hTC0b9WGI2U
Uh5YCCUlDXD7IuTcQFykDxffR0713n4mzJQ8RzevFqQ2HkOMbKCVIf8SEwDEwxy6
Fh97UYWUwh2wjX7hNReH2NvOL//tMRZp78ojOcNDxYjmYrIoXVt7lcqSVHlHb9pe
0B8TykQAfqGinCCIHruECSGCd6J0GSNbVsuOkX1fwrq1vmjENsVyxnI9ha1tQMvs
HWjdYk3FfU3Sk+mpzJOrf4eVkHLUQEHAr9uxpGX8O/+U1Ef8zQSZmCbosmjfiFF2
FKXAzhMUl7L0r7z64EoSLs2Udl54TAhOY+NBkgAynjImzpB+FhMBRGe5H/F+3qvA
ptOBoisbtBSaEnbrPFgrQhV2RUtCL35Xf1rw4zPiqwV/TTvwTXnwyZymKs7jRzQ2
KZecMh6iFWqIIMIlZLSpWg==
`protect END_PROTECTED

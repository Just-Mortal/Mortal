`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QQnci2z7piW2T8F+GJt5cOFJTvJZ/GuYbMgCdsMgWhhOsLcYi7ZF7dsb6afB/Bt1
kWaYBVrCRA1cE2Zser/1F8K1JohOIIDL2XCPXHQGMraiAkAgbpB9Q8qhHXhmC+/M
pvkq1aT6N7K3fAMn3YPzi6qL2mMezeZyM3t9EhLu5zDA4NrX9E7XReEJ9zw6CLao
UJhew3aaUitR4g3k6KsviL6vL/meJxTtejycbr4xH+gw57CdAVdFEZMUgLhSUa8V
B9RFPXxtgomIGDIT0L21P9J9zZFoQLLU9pYn9S9SbjTIvjE1dzvrYD8MipQeCTN+
x+sStuprcCE9q1mkFWKmtTuKOOsyyhlLiGbBbnBnnbJSbgTFCUfp1dvy4OiCj125
Qb/WPqW8m0fShtkZfTj/A2//CxBb958VPfcogaDakRZwYh5B3q7f5Fnz9GJ+Mc1W
9FBIZjwOTOR5nZzcCUzQyHn5h6aG5rqPOfD5y5HfzPcadZoQzt/AIvaidmMGdnjy
k9ydbrbn07dFmKFtOdE3vFWMR2zWC/A8hfCDst10pTpfkA+2k6+MFfcCad37oLb/
F50N7hr+g3yZ6a3tRiWK80CzDmq3WA8np51x7dP27f4pP9D1l1/k3md5svwcAF/1
0QE5E3MCYHfKEk/S5JQfUwPZQxilXV7sfvvlpQ11li3AEgCdJPRqXSVxc05S0iOn
Z3vTFIbtwFwT+l/aMXNEePuYdDzC1+B3rZYwfyHJIxdOmGH9bvx48NZxOWROx44g
jmMgHlwPA//cX1lopPCAysFPP+mRaYIQvBsvUPsyysqdPgFNahjJrQHK8L8GeLgS
BZrWqoWuS3sOx5l2I+fLY+S7qSMLsRokeLbtQGTbC8gqRNiguF9hCxq6eYb1RWXe
qklx/tdtjcKzu0m7A5J4LBKxNJTVsldGq5Ze0M6I0zTirwP8CY9uTbpaUSgwrC9x
dl962o6n1FD8MCRYK2Yjr9t+HNIUGq7+Ym20+sIKN7Ku6aBF74Fad0RvZgrJlAWr
FXe5DWZx040NSOvX1j905Uzf9vz+V4Ke4FJTRpxlE0gPoC5+RIC2aTcIqtzPxhJK
bDCiSMbXonhJOht1BJ+U05Syo3zHEcxFxRKU8IExa7TjY7U3eBLZIRGNj+QfvO0R
nniM6LgnpiW7G3DjWHuz4B5CMy/Sf43RPGPuqovDkKrIbp76Sq9ei1ubmFHRaX/o
Ano40SAjms7gGCARGyMGwEGuthrTO8uaFsry7vyLlSiAHzkTBjk2NAkJ3X/Iy8zc
yA5M7yC+mWxkPGMkDcVvBrwPdnTEVbPjcsLz8oDU6zzjrsVtnoLbODwbXyq7447G
NCp3xR44+3bOMKYTcnIJEZ2+wml/9CAdf3K1bHHJpB03Ed7h5sXd7+GlVsAS1sGJ
Ddj4YVJ80rdpZDVKhzOUMA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZuS+umLXyACeseUcxGVWqVvEdn/p1UKgIaycmOlf/5RNfFRs9FZZaSnLLyLOFTM
G2mtP5kk79nd3r8DELl0RPQN0i297ecfyTMEquDu+D/AwvwpWDG6F+2iak32jx0b
h40V+TrgqRC74JhbOMf6cJLDUAGboZ0QtdIY2ikSsO2I++mChIULDLeMn+CiPySl
9zMBfBfTSNMqjXWrqVEwYDDGcIkgOz4ZffWHACkvV087RyZX74Rec+imL7vDucfP
91MLzTUuB1+0GtjcrYIF+QqfFl6i8k+cb85+WAyY1Nm79+oxYsMrmI12AYdUB/+w
gmXeXkIL1Mm6IxUjLvvoVva8MJzlpkUKD/Qb0B/HMcP260Nx9VkqQU73q9icn5Uz
+48YJO3a9xi4MOipQGjLMJNaP9iddlGiH/KiM1k+3vlLtx0BgkMqwIr2XNTGnesA
nCVSsv0tlU2HXvnBnjUgQQ==
`protect END_PROTECTED

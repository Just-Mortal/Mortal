`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJrzTQ69NhMT9swVNECbvpzq5RAH0iYehfqC8I/7Sg8E5CzxlyKtaXVLhOXoaLcW
8nmLEBNUNlC9vmy8Zcjz1y1TZ0iJQqAXFcq6NWMcMeExuW4TEZbxCzssrd2ZLlXt
Bxldbx09EV6CUFzpkUV4pIEsL6SHhNwab5WsSsWuCTThqVr1xwZK6MPoglarAKOi
5JeeuN5QSiNUCplEhPSUXZv7otcUoB7q6Iuos/4knTT0AohlWuLapsyVB1GZUUrR
Ii8iqusZMM9RrW7OkFY//1OuNbH3/S231HCRlfmOeed1HmCa41vJwT78BCeNsbkp
ONkuKUlGxkcpIkmlyWDElJ3mnAVdSDpNyGeRULCvjKOCH70bZ5NdlvFdxAIPqeon
bCWQwPSZBD33s9hHteJ+ejTqJiTwfHP1pEojbqD2zoIuEkKkQ23mZ2jUHQG6r19r
FBJkNqStaePeQpNWATTsLmvv+kZA1bC3fuarDA+CubXv6fljCm9Pj87K8FzRasMV
/xM01a+2E2WjmBdHx8iMCUFz/BK42YdXCmlAUERSnrNyA8gVR0WOHifrb6ZRa8+q
zF3UKQmcCe+yBFFRm60QD4usLY19W8rAjjoWd9YcU3JYi5PssWoXTRA0p8CgQccm
+71uINnwIX6Np6fq+pg+w7SMRXfKgUo9EgKZal2IHZkw3YQxnWlkkKlewPUem8Ua
DFhVTcJKK/qFxpU3nf/8xwFNp+EmEyXUjT9cnn3ZkLxQ2G5InP6gjDYzyjbhH8q9
IRhgepkb2AesWBS0kmLo42Kx7yBfv6+9sugeo1mnvh1V66yUIJ6LL31p+Mz3MOgb
Y8W3dKiLW2YpV1QTrQwtcMzmPyhPzKAU4J92Ip3lVsaO3aw+lbSOPCPs9hgepnuF
03B8KWCjWvs4rHly4Reimd/3uMVuo2J5M/OcqQOFb7hkI/TdOocMhCydTLpjjUL4
`protect END_PROTECTED

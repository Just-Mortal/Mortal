`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+JuGzu1RgYCPw0CDzU4ORxic40qfnQqojnxXru6TVsIb+L/px2cfCg7ZQGy5hghP
K1pVmcrv0WY2JQri1Pk/WTWIx/BFO9FJmMHyb9MoNA+py6MDtnKFXFHidqV8/Zxc
NjW+1eiu+cYk03T5ov2l9+JRNx4TaFVzaWDYSeB0R9MMO1j+pM1XoIgwTzqK0/qA
nYWKv976CQw0zYSLjbo7FbnBTFN4zKx1vZtd0yf2y5Vtth7gTZvsTq20LYwa/Wh5
a+kFIomBc0SnzmdrSdVRzMHiD5TThzRV5dNuLV83+nTuDVc+svRBDlV3CI9aoUwC
NTd+nx/yOTGu0PQGQTaC6fVIy/Gcrd960p8JjzFd762OTAE93Mq+XeeV59QqIzCP
LI3iOk8X/PfFVr4me36LG2kpH383+70CAiPtlS9KhmK6za6dtOTQFubSaWLrLtEc
GIsY+zP5HOex8YGRSjcaH63sdx2IdGGvdsarVtc5FI/htRBpb5iugC6XSlt2jW6c
p/g/qczXLyLDK1KVlUduenkbbfyURBU+uKOVgh4qwIIrgmeFy2hErHxBbQCfyfEH
j7M9hus3Jwu0cIBKaYt6Mz8Xu9eBl2w/Jjlaz8U6PnJv8co1yKohZXBc5ewAvr3+
nPgyFEj9Z4Feq7zikF50GaZ+sM+UIJ0Fr22k/1ajMqFa39aWUN33gp3wa9zWHb1F
89siCJXVUCf43r22h9hIzvP7DwO8mb2hXNQfys7AMydaSr6lyeNre09piPWzse7/
XWUMPYwLkUoq+FQdcLFA5rWbKMSX9zWqh/lFUi5BTmq8TTdJA9sgXac9OzwjXTBw
5O1AYFm5vh2Lho4oEge55DaOyBDSgtHn5tH1KmdPfDgdUT1xt0aGaqzNOEnOBccn
8LxPLLRQQH7xx9EwCAjllDGY7suK1qYFnoylcFRrU6AeuIHs2QWjORwp/mLHf+OC
+r8umlHlpNdNNUvsjk2cv1UyqIpfp019TMD0TcePP6tl09UQ2t44agjf+J07xD+w
R8cxBMPWjv7RbuVzd3aaRCKOu+FlTjIvkt/rE49A5uqUszDdbHpEFjjEZRcXOvqi
R+I//QfP+PU5gf68NEPVdxT5YdYVgtM/v/z45T1WBVAMiDP6/lZrxvCi/KORL2iR
asvfqR4/HiQS0pnFZt5tROBo5RRLclvFH11JWy+wzhp2kaSMSazw6WupX9GGqw+2
tSmqw7zcIHCjz+p43kP0qaS8RyPQh1AKivjih5s5Bxq4ENU+of1teuv1fjhONy+W
0wDSid4gw1RgiP3z7Mtjz3UTUTkTEi0f5Wub3EConV9FIm8bqr37o1+a+lufTFdT
DuXMiyJ2bJDZbIXP9fgaaBgh/OJzhG/YbK8rNsADF1kM/NB8+k67GH8hTQhthdyj
102p8PHABT0ZDK8C5yeTh1kXEiaZtWlogTTZIbXO88LT/EbSnTObJ+cekNrav7C6
gv6eTabRANjew3EnGpigs4mJ8s4STJxw8EtX7I4dwlC1sE1h1KJc2qXprkFX3ps+
jwFnkgy0uVZGbI5cfZFLY2ijMdwSlWw5w2BTmA43Obq12w1Ot4EbqBt2dP/LOtwG
Q+T1fwiFne/W04ubkMBzERQ5sm3y21TQ5OLbprl88r4HP5eLeUudmUYSQXvlbl5i
4Zt0rKsWp94njdptH1KhEYEJOgieUCtO36qGHPmKpiSk90M3vFbEmcUqs4kFSYLk
g8pqd1jKrrQXBf/hAj4fRUqCQ/hzXz3BMgqo9dIP/H8z1hKJ2vrRRz+OH9RUbkRr
ls5Vu0iq0jvNTg+F4+6grQAJVa3UHol1KmhW4YB91mQgJb+EK6HKYYTFd6mBLQW8
bMw1q75qa7IuEcGspkJ+Iw091GzcLWBteT+DKX4YSAH8ixjRTXY7f7llMZk+w7Z/
eI0CjUxFt4G1s5LYOVj5qZ8EWTk6GVpROF4+GFCWIIRfavDrErSnmoYF/0Lh7CH/
w8FrTj36ag5v3LA3ARchymMT2oB1PpVRCvPQST8137iPjJOUFjcrlxLrMY1vNx+i
k4OWcbIHxM9jHOxHphH5pUmgfYUfsg/3QiBd8rHJyPdDlBDCuOyxcL3cvFjLmlVF
qzXoGHOlhx8uRj/zc4en8NQT3EbFpihnKdoyBHofo3UXYB6NHAgpRnGBrroeJePf
bWii7kf4hzSDnDKdY8PzD5HjV2YO+38CKlL4jWt2tHWZqAtG9on9vbHBuaIN4tFI
pPRU9Od0VEMMo+yCCBOhQkCGwM1IUX4yJuLqpgg1Cu2U3kMU9+yIlxGXP+VXfe/D
fVf6X2SRrVd0BOZTYi4dqTofUu8P9/TYu2XHCdNJrY18bXCmXf2KKfmvP1oay5EX
RznrBaMbWUcvdVAe2jh4+cN1tgJouIyd5EJP2i8DAtOAbkC8VoslzhjxUbCOqeut
/zBXuEL5B6tFy1+S2ithLFLxNHqjwS3hzO4QfigNiFc8n237PgJv2JLVXszXk6rZ
b2LiSMFflTTP+XNVIkNM+PwtfkI52uwxkNY9K23jvsTRt032NwnVE1vOKyC/UnVA
l3UkSPHT1Hj3x879KloxA8CX0ZOZpj848EZPBxCPcKTPKMFm4zh3r3i3eBpkq4nD
7aouwPg2QQ8TeV2bfmaoLns8rQCQVo9TfNv9/7iMcoe+wHS5bvRN4EmgxcWl0GhO
S6vOSAYN8sG5b+rEnPcLGde5G4qO8fUQlOLih0Cke9w3oXcgyEd+trwmb15XK1IR
5Zv69Kde7nlmfnfCj8D0eEXzJOgkpR8XwBiwnZ3UVQ2QmiE1cteWusJ/TupnsMeD
p930y4IJxRoTtynk+Z7JJ0Jfnd4r5QViteOt/LEY3UBFypeOrwjaFGq9xg58+zqg
k5u5WPs2/dX+szvDhMYzI6ZzyYEobBdvbRNgplmRC0xqe8kgm0QBTgq1DmnhhVOJ
kY49knY/4UMlyS9M5mZx7qy/n7WpnNl6V7KgRcMbtsEWDhnYyb2pWS+NVa3CSY9s
pcZJ1O1PnLkHLcTdzaF1BtqrVkdSlYG42cU91eqypZx9nIIh2q8eTBhu1MFbStfa
MZ113Y74xaK6hMM/HvEmGpEFoyOBiWakjVw7xSHililakeZUWN4Qn2mBGLVBAnYD
Jo8psnmS6yel68qin2gPg/TtdNpwFRVqXkWYVFP3LodoZx9sWM/Q3obxvBJW9nTs
g8CrN/bSEvo0yEMI312jPfjZFrxmhmBFy7rWzUJbr41aF0pwspg+43sDGwEK9FFH
HGTdk4/VrtmiTBSPXH4dgKjCwvcInhkgA7g3iBQWXs/WwTMHiC1K9YJiOjp334tu
89ZDPd6QfFDwh8axoDKpgAToSrL+hMR5Q0ks0IlO17/mWDnvmaTAfTz+D40MnsTH
`protect END_PROTECTED

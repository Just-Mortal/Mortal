`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gNw3c1215IcTzU7FuNlBAm5yUZc43DxjIHFsltAaAenKxEfyGeE6gRmKJCqfl9wM
C4QDamgYhTPTXxa178cKlv5vTR22QVJf1hh8bpRa7Fgs7NqEPPyiT30RKsNojaJY
rI+V/To2A+7qtuP1/xOjUBVZarg7uQbZN0C+4r3MCBqtDWRlSrIkHRA++uP6EHlH
uOfCF31JuKlISIH8v6UW2SGwrECiVYNzaA153dAVthSuoKH+raZBNeqTaP+0yXOY
GWGw/01EQQ8DtHE6Ed29XD6fKxSwiuhxQXxV/wDPlRC9p/bsx96Ot4HD3/6fvne1
B+EIdea0X0XgWL5m9iid25ArFFynl11o8Vyci9dv5n3jzQ/uYlzFHyPvrRHW5Wmd
BuGgPendRCJOBqomtmJtSnbTtghjVyvV3//ySUBEq9/MQrFmz7sfhexBHFijlK1o
hklnhpJoNNct0Z0LtWblT5lGFgXRwakMnyXKof+QenureYSxfAsXeCoS488miJC0
P143HUDR1uyjZd+nDHQhxL7myAqSOMQ70wbMgZEZfPTljMx9M5l9Wtf6/N0idss6
GtspeaMXAEJeN1PDIxEvWunEGVbH7WGXgEHEFH74dIhZtTZsW5VNV8vwn82xDyX7
3lflGq/bBQvcGSQZdeesDArTt2uC51aU/+qqV1AKJRLt/4HnaJNKgIgcXBD7h6oI
pmfUTsOAiYztVZl8Xt+aooV+LmDiLoeWW8yNk6n2AgvHGCYC8ngAH7rnxKznEbmx
T0M9wLMBag2/ccpQg54p2ilOt27GM/i/LbHm3zMzFGWElFfeDwK/Uflyie39xMJd
z3u0FBHj+RHf+TtyZoaAGxoOKnpPIl/kZ9+euGd6jX/SOsqRLYIVOv1g3vT3g8PD
0TR/5GdBcc0bzD2v7eR66q7qvFjEwX+hOMo16Kkwvk1T8Q/QmbFCFBpQy63HuLfr
WBd5Zufz6kqv5XHELIwTFzyWvSnogpQVwfwQl7BLqV7Z1sQ9vm5HSqZLqJT9zVeA
2mKmYLCr9cIFr6aky2DYDOMHy9x6QffTFmR/HgiwoGPM71t794rWdOquI9bI6ibx
8Y8bHBduP6ZPX6vdIPIa1q47oKzaBPVShVVIKJEGZ7HZwmw17ElDqfR4YKYSfLbx
GLbzlfKUpxWyqsaTcy5dsUKOqtg4Iz94tZKB/Z6mCGwgVIu7V7ql6SvVtr59Z9s0
UggarZvlfwbWVUAY4yL5Ua5U82z1PTKHQoDKNMdtOEyeTdGBK3ynNlg4/2rVp9tp
86L+Y8lFk8TYrAUWYjMgCT1bCaWMybXrQUWNpEzqtqDesrbZXvBES9CuVb+j3otF
ABAOjdS3ac8sh8uYASiP5peM2n0qnrLVcMSy30mYF+vBjS6DXLmWUrDx7h2NXEja
AFtGivlz4JyXCGaW4Ghg+P4lrYb9e9YNZSv8fvQIBdPW9sfkXkaAOwMQBwc4ysVg
PYB/2p5thXzpJNX2tBKJvKePVkZm3jMSzP/QLoBvBqPMtx7UImKdB67UBboPNt/+
RHhK33ukuYmwYH8oW5BLPDSe4VWOO49YB8aHsLdsYFmEowcwEjNuo/nD4Ur8kM/d
WNrldB1BIA+2EYUOAOzhk31NHYZRwAU3fRcAUqPQN+qZ8uQKM6afxD0p7yt6JKI4
4hqJcm0jlpb6Pa+/1gP3eyJSRttwOVYivJg4KZt+xCcIeDcuzIB0NrVr1hujQ9qP
5u0wIiZkQezpYTr2ZooIKF/ZeF4WU2vWfMdzLULEEeft7DgT8bI48IN/1L/md/8o
kc1IS49Albdt/g5BpUQpJwVUnke67bQYUvgvUQDzjLtE5dzHlAe21j3qJUrotLrS
L9JXxw+TRv5KXH1IMf7iLYlq4VAixca9qydDxupysK27L+hfzOMskQq/cNqrhBQ6
bvVVregsdIE/cYCrQR/e9tR1kMIECxp9Lngeab5iKoJwac9+jIJYR+DF+Nqqho0t
4LtdQxsiEUe5anoIZhzBlxI9wN4JtbYDDlEaMjmYHh1OYO7ym9YLHT3G6Gk7GDVF
vI1gCzU4f1SMDMGNoPKPlhKnFa8pa+ZHCzFuj5ZDz7iHFe+AfnCjgrfVi1IHrh1J
583kUdOwrtmjQVnlmKinSjdJMFW03rKRQO/qQ+un9TO/rBHq7N3I06YvdqHg4Xsz
mviaE3cmKK2rnONR+zoy2HvjuDVpmGkptP6RbOj4ZdQJHD5uFzPHS9/Ed56UcDdB
yZawD4dAOJZRiVPA0hwd0h6yyoggAyvPgqpruXkuqeJ0B5lnlVeUClB/ePcJ+1WP
hUUxQVfThlexSKSurQiNLYyjBPD3+V3ttuiwN2CeV15ugFspNk91fgWdIAARi4VG
wew+s0OMgoRK0wmTRwg43GoP4b8IRanD9LCOeV3q18grb5+BZhUdlmS2gAiwnwFr
HBydEX/scNLvmzQWNX7lhbRgD3vcYtw4BU0iEhd9syNvpnjI9Wa5LPripzJw7XqI
2FQQfv9MV4mL38N5FYRsqFLVEb3iYF/u+4Co21p486HDEnPUyLt3oC+E8NpHbi3i
7cGrrnzSHQFFNW/zkj+Fp0g+5tWy/25ynlI7MMD+s+uPspXzsxpAWU7FpwwsrPw8
vdC1kUTizaRWxwq0sOMAM/KbaOM13EP09NJ+TBkizxmkvq8KLP73TmM8KdBKd7K1
Lh9WY158jJqDo8iV4XgwTd2RBfd+og+W0IquugzyIATz3/14I4arIy8Qc2YDA+1l
P0V0N2GsMrjUzy4JbUNM0HnZnoggzRX/HrK5MNHSLPaVk+/jQm/rUbXMiUhVDeIP
SUZUw0dF7IRdXJhuFy5iuCbfoG4sX0w3shktqIgE4BKrtLnTEgo4Mo0VM2vNGSEU
Cx/fyjhIWlsQrXjfgEK9TogY3j6oG/ewGiZUNC9iahzjPIDlhl50FY5CjDmkYEeC
XR+bDq17ISPoIM7TOQeYHj04TV6tYAnWui0sO7LkgDecPI32LPe/xSDpuhHHF+jf
ZAp6LhVFw85SFiIhJtBVnBN2eeQF+wu8U/8noEv5uscR/iQ8d7uQ5hP7U02LLeR8
AojV3esyjPWlxZJGuRyRAvRJwNs/1w0kC7oRFvn5Z7+sIviTPoviaBEapaKjff9e
b6CB0L+z3yHoJj+8UwLMsvbH8z9jIXkoeKmFkRQ88DW+E2IovR0ibZkj2uggDszX
sZcvyBjo8M3k3ZyVzUo6ZT3f1I8IRgZpGn0/LXwXyH06a7hSvwlS6V3N5v4OwajF
bm4JVtjGBVk8pVjAgx+DDeUv1KG8LyGzwd3n6Pqd4H+pdwkT7K5bZHehCJ69kawM
yQqUtdUbJPi/vtMnoBlzGsxYlXtktNtxMCF0vWFeDFbbpdDEWGcXO8QYKM3jFX/K
NqMQ7gdKaTdXNXpZoAAykSYERCkIj0EKG3aUfLjo2dD15I9ELOuYUnzzGNg0daMu
NfJ0nBi8DutCbEOMGwmcS66oizFeNvytDLCoBUx5HT2kT0nayNrjFxGhpmcnf8v0
Q7sAR2x2CLcXuv2gDeUR6cv9fZF5ke+dN1ikhTzSGfrxR6wEIHB8Vaos8SHJi1Sf
X1cHCjDCKG2nMF7Q0/OGrBfqfir+B4QIE0XLfAwrV2yjOwE6z0TE2+ybXeCrUpso
7oNG4KsFk89BkRuTB185rGEzIU0Jh1g8sBTYLkxvJZTori1iMD0kesWtfiCE4Lch
honPhhe3d79zwdkxAMmqAiDCR+a0eN0ZiD89aLFtQ3oHjkVxjkY6aQXMRo56dxzx
d4+PVF9RZuBzMD3uHHYYvKKM+yDYsEf/bPPx+gmhhmZl3P+68QjQu3rlFhqjygpI
kBPxMB8H87O1q1MIZg6k+aNgk61huj0tVXD+Y0u12b0s6HOume9XrqCHU1U16RVJ
HNMneBiy7Vwk9C3yWhzAxRphnyliqa5lbPQ2LDl7WzKeN3vyfVrxz7fO0ZqUWOyR
/dws69CjqMkEjQdM3tvEZO5bKCh/KnssW6GpVRunrqkIzx1G9M+6fJWfUvXVDba0
IT9Ci8huwX507o2OVrEIL3a8v3iTFSxaNJ4o49Wehn/Gudi/SkYRrUqq+PWn+BMP
eqLynDTgEohgX5GeeVlRYZ3gQvrjTNW7VlqI+hgcjyvu+ILaPQf5gGRF7r0st4fM
bjvTFgGca+OzqTidTHNFNancwiWrH/MPZfPiCOD3mhRTqS+cHWktiJxC5dLBe6/T
ppkS6mReDKVDo5kXT6+du7sqfEvhFL01EudRMtiOZCXZvCYc2TpVpjdnh3PgtG0n
mcU/2luPhgik/7qLJ6WEHfjC7zqtY7EzcabcWbhd54o8PP2TDMgvfaWYK0LiD/cb
6l2zAzvhK1JEVIW7vu/WyPehm8bhT/dJF1RkXJt0O7sj7Kxpf9q4Lo34V0zyl04T
SK8gdCNkmYFgkrXKH8TCagtegTckFAC2lZEVTIaTwBIByo16zeLLX3rEEER9FaOW
1u6Ggo7xUT61+x6AyvxqyTRGPsfjxqr3HgT2QCatAUL3JsPvJ4TO+J5twz8udzLf
uIb8LwZ7Y7JWPM/UmrUgXCqGtH9smvNwbAm68VGvyRw7a9HP3GUE+KB0iRveINbF
AcTBMGLs1mzPVmYd4G26WQ+lqloP++Ut/JbvjW7Uo9bmNL/u/us9AA5lJ07pNtVM
CwqgnUjk17SO8psf1LCms/TiwyCaYHRnKKHmXXj9ogtPElzYTyD88UevT6EPy5yV
pPNhMa4gEZ/PVjJv22oqaHTtVf78dxDteCTaXxnoWnXoD3JCkRVU5yuAYLODjfjl
2ymLMZIAF7sjaYzT9s1ICFv50upiSl0HyNgm6kiOWzAih+YgylYncS8Gt3T+807p
B2gQYeQJ3tEFGApHLvBicKMYLCLkw4L2GK9ewy/QE/nIv1zDnuxORjCLS4JwsthD
lMFxIQO5uZpEOm0BlPY+NW9j14LEvG0/k3FTp+KF6zTcJTxNZmqWLvo0f14fTZOI
Gc6Tsj//ZQNvpQwSWkxwVTbrW8WK98XDwGWTXmwI4CgColcPn+1K/icNV8eB3ino
c2Nmf8aB5hKWTZ3yzl2hhNOEmFbS6qFNygAqzvYTGNwzz3y/h7SS9phwmZoao3gZ
X+Wi4UAn9sFoKukasDJ4jfNVSVOE3u8+xwmiAg9GozrB3oLWTfk0/bL/t/G1nJ3B
FK5Lw/AHZOypyCmDTtmWngL6z0CiOgPvWE9glzwinXHVgJhCR0SU8+CfYnNS/ZkP
D6dF4yMwXi1CeaqHKMihydGXgBM55HrVTSdw9HMUgHyY8eute95wMQ73S2FpCvTi
IEFUDgFuLMgGp+pg9TCStPFOuKjF3M40lFuXr/VNn29UDGYDOk+RagAVZqNWgAnq
7fXPw2Psz8gW+C7WPwatre8a2ykL1HOCjUtVA3LV7+kNwLv3WyfC8nBRvNi47zY/
g4IlvImYOU+Zf4EWgTdVZ2sPLpG0oUjF6lNZ/biVEoE/fP3fIa401ePRFKJm+8Zk
bNq/LirPRkOJaxlRj1RocudoiNwTEoPi9FVUnWo5IxAySJN92bttsZTpeDVW8FuG
xYgc6iBcd4vQaEw4WbJN1YXNNG6Z3tQ8BYhoJYOFuTottL/CFnQh3ycWPFYLLUCo
c8uea6cYHEr46pl0lp7VpSHDSc4fGWmEvxVd7efR3RRTdEBH1/R5TCDtlMgp3aif
pqshazpDGTYOmVejv/LbrWctDdGnLQl5rmSckWZgWuGT6uA2T/o/5ARp9z6zYtc6
QVZOiSiICC0S3jOaVVUCORj33FVQFuNPQcb4JKgpEGwaY4YggMUPVSLvWYtu1LNo
183EbYcBgHDHoLKkljcAFgY9MIHg72c72rsQ5EIh1ReLXwaS4MECMFL5srCkzhmx
tU58C2hm/mRSrvealaoxKi+RsKdk315NnWeI+DCFrvd7q6VYHSUTSXScoLbYM4hq
9NYWZtTtrsOtYzC/XzjzgIX6WyDYMZlqVWQnRdVKMit22gxUjILIsRZI0R/Vufjm
uhUsYfWFBvx7zie/d7YCI4GZEdzxtZEh/t+5xsM8khS88bJVkujLEJPkMMZKb+MV
dlZTkP2sRh5qWPO+yYv4AL0cScDAT/5pPMNNLQzZxyfK2dEw1MADfGJmQ2oPoz7B
B/XEVnnaUPy9+hDqoihOmQ1TLm/hZfAvnOuUBxr+0Zhr3wZ47cLIz0+uWbWpJiox
JEj/PFyBe/05oJ1aONW9DNtfF6+oT6XUHGBcf8f6uXu+h4L4X2E34+iejOhUYE1O
m1Dro2am3GGI+cvdYxF1pyj5cd6SO8aztlxrRqTShR7DB1bmpnBh7sTFjjtZkrSE
yXo2tJYsK+9JV68z1OqNxlWVh/H7IcFZhzUuJvhIYWQ9+d22SHmOuRfj72vwkX5T
TvCcGaffNTNpZR5lklxgo9O/tmE7UQ1QZYM6ZXumG/IBccD7REZ1NvpUjeCZ/6RW
g2zA+DymmGs90V47EVqMESQsXYa4sXMEvF5G+YqXEyb2oSs0Ic3SzuLua6MSzxay
tFwOerJyXWEPYG1PLZWUO95GChQsE9NNSe3mID2RmHzw+tIoDwWxodM53OEFZYXz
dEqFcdBko6ahxDu/K3ax/5euHZ3LXuDS0ADQXgv5n1kYX7pGOXteGbzqQ3r1ymHh
g1VDKZ5X+VCEY+Q2IomEDubcmJJ0ZRTAW7QPQS59IqP/9oT8xLyPlYiD0fnatQ5p
l6L+W0PA1GqBlmjYz5hIuEuc+ZAvdhj+Ex7Vkdi7R9pErnhMLdpgiZJCehdd0s4I
fSKifqgyewJp8dKePyJnqbli4aRd3RmuoVSbHDW2mjMTCnKxOlnP1We09adeBzzm
iqLzQycX/42YPPAsjq5n/KUzk5OIzKxHgkhXdiac25lRT73McGu9hYPtzH2OlyDd
LNI1RbBqC+LSIsnOb2KSHUGMeLG51FJrkxbHFbfOO5T/OgQF30twC2kdXU9wme60
Q/5W2RI/ABjVSgCNjmLOBO7GDmvNUXKQHo8P4fkjyx5mrh5hCpA3+/3t8Q25EPyp
0yt7zYb88PAgbwJDGAhwouGzlhVKVcP8Q3Hfjk57nBIjK/NrTQ4O1js+kZEBUNvV
53S+CZsH2Ggs/sIPGh7IbS0mWvdZ1M8+yMKh/9O2eS2HNzZjjJ3QmmgvqOOm0ilV
lWsh91W4Dee7Q+KgFc/xilHuDMwr1keCrs3o4M0dX125Lndj6y+R+DIWwGFGCySc
UdP3hOnhZCG31IZAu9xaBnsgQIHXtJKgnID58CpcGWBeEla30mH+KN+LG3MZn1z6
xKVzO0e0Wq7HpTUUwq1o82SrV6jcmZqtmQ1pHY5cnjAxe9DqU2PBwhIZJGPDYSqb
gofiav7WN8ReeA/eQTKQL2eGpB0L3XGgts7H01mcX4/4/07fLngqizZoDJWHoJbt
hnOKPk/JqnokuoR0CnCcbEzJFHstAODJf/Qk/RdSgB3HcHYi8rFh0neOQ37zZKOh
qna1LIATefIWKTn9q+l7l1cGAOCO8zftXIUjKdGySbo5Q1ApwQdeXBudikCFCZT7
6CiklsModkUpPLbNKucDdV4bxtpwQF69JZHVDynuXgAy6E/A27i37HXnblAqtPsL
gVagKh3GEj14Ju1+QeHAzKEXuEuOX4bvp+ldXoJhEZOMc18J10P64CRJFVz+O9ei
kcXMog+1pCmExcYFiTbSteWi3O2X/aKEykgqAyOwqCXcPI/sWhpNxZt8A3mr0T6G
AGPQNo9qB8zbKu1+cUIglDn7Tkh39omD1iRvsN4spJZQH9mS6wEp94wQVXGmqpkV
MiaT7UQigwpN60pNWUynKl3ILOtpewdBZIcJd/0BXIeyUEsVcMG9bWPxoiqxlBYv
v9nLBjsn/kgr5PRhXyQHIy/HfhS6GS4saivbiex9588oJVtggt66qed7gArUQoVZ
umKxBboCPpNJdu5PK3IkDdoUsG4dPvQeQfyWtJGYCEHpdV0WOwzWeRTiwe3lJvgI
C49iCH2t67EbxciltTb6Mgof3YZaHLsox3y7TRtInAwvizSd6vOLFLyNk8LmdMkN
T+KSlDn0eHYiKdKjWE3h2zIx3G6X4e5IM1cm+GolBx8qZ+gCjxV6Vit4hHqGSYa7
8MhKHODUxqknLFRcRUodTOwLcsxxIVnM2MIFhEaWRMfXeRHhCtHXPD1R4TunywKT
Hka5OIBnXjiE1hvVUnfk/o0L90/BmUZmswPhUklnNjiRCNdiXpzMEoJnXRI/2SqQ
jWW/IJUy3/+2c8yP16RHHRj5tISCrPLZXj0gPg6Aof8hiufQoHHSmboxcCCjgV7/
TTu7Nfw6rLyVn/O+wktQtbdTlUbRt6HDX9VKVdEJmrEBaO8PIo/Nbzx7AsRr44f4
zlBCHLFnOwQQRqhLJDqmMMwPp4K3UEO9iz4yCB8NMqIfVr5pLzgMyi87s1bdLgtL
VNmHCEdA8vS4E3ilzvLUZZl4POlaemrrdFb4Wf+2ydJhBuBoFXwPEixLyDoQeQlw
3BFNbtcNA0K1IahtCasGRitSgw1qo05JP8l8IWWhDliv5QFyqr0xGrQjMy2NGNPy
pY8xYWzUhaSlAMFeFQD/OiKHuI0eeOnMVHwirdrvpc2GwJhDRHAyK2dIDS8vvHjA
HkE2kRxUN+6H4tYSP+iS9cCo7g8v0mafhhsRnhcqY9G4Hw6fQpbkBMMvAANmYB3J
li5NdnbMZvSrVB7+qMVe+/cTVkaAlnKu7Sk+plTyZ6fRsclh/woaJAz8bAsOErRH
bDsOdhStETWkRXLgqdiOO4DSXi4naq4nVU36ify0V1cUe6HRKhGldLiDkkp/027K
miLsEQ0uXvaG/YRLOasuhcQYNlzQ+4fCahH0ZHLDmD2buo01RmjgDysUbJdziaKz
MbIP5RRCZN6Sj9ftPWcMQXwYJMXhrLK71zcYYcAu2un+iNOMrsmT+C40LvWFa8gQ
el4y+QGs82s9x9ilIft+rQ3jAI1zGy3gMNDFPcJ9eepBn0mWUmrTH0N/eQkxH54X
xgHvx3VMOoUG4eb6sYM87SJQPmIxhVODa10NxPQqE5ckR381T2ZcncYxw67oPckc
DWzG9yiY6SOkwHZPQivrsJM2XUi83afcUJyvVH8RlBpex8GGGWD04VM64QeaCqc/
3f7vJcdb8pC/VcFtm6zT/7ChqNEXmOKOfeeg+jeNWw2EDO9jxBho1Jf7lHrRXjS6
M4P7A7FvimRdgXEkP7nASTXp0UHqPdubet/upyt/1yUACSiX+MrO2lRagWNkv0F9
vzsv2jKoS+t6jopyuHliXNEbSfi6qv04lyAdmkDip3j6J0Z3i+hB4C8N4SGepzeU
T73kwAQRd9aGvOWbcJyQcmnWz63TZzKqXAMrANiWh4mVzfpdW9VrU/0E/ywEkFl1
xGB03yibfRUkg4HfgCDAd90NspViySW66tqpMljth/BD7AmKae5cHsPieCOjbIs5
e+aYo4hAkLIPa/MMqy6IcD6FCZtCuwuiFbbYtd5FiRse84CdbTdGHcl0eQ2ZgHqO
IhGVURFtnrLD8Pyb6M4nGv9LmeFTnb2KbmAVB5W4UnmHaf300Yv9KMlZZhN7sReE
ZZYFU63sqPQOO0xvWY3vfurA6XoWWibFp97+sNdbM81+8ndx/H86djpINLfqyyvU
7ENBhUokmjz7i6rORogbnfrM+RpA3j4Lan4WJc+tmkZl+HgOv7Sam9XkYzil3v6p
rW/lCuhvqyuBvLPBvmBZk/xJ5Sb4qU2qnFLe3IvuvdZm5mZD8tNyyXNOkwIsahSe
vq1AO5woWxzfExN1zDqf4n6uUyJXR40E+indTjbq1oqqoH5Cid+wBBmEXSVEVLTC
orULtMUBDemiiVeAVaWuXEAAs2FuIDGZdcXZWwuP8P+acI39O9j3e1vZsRscWS54
YwtZtzR36dpYFnLepGUkmvb1cn33M+wVMGG5YwhWIl+6xNNGQjb3YykxTlSXi+6n
2A2z0IR57n7g3uZV5armz/98d98ZJH2tloP9NzpBOU5Fx2lF/tnVIy0fuB/Qa2Fx
x0GKaGJPa029x+hUx1mSAjiOWIA92qjTQI7tl97nCaRUoEQ4/TTCQvZQWNyoLu6u
jfurM2vHDxd/+RWetC8weejLuy2eGqHc1rMuls9snIB1ymVuwh0hOgt/bRWqMYD+
yfu1qjlGrQWTkqsZwToJXKbGMw2Ew+q7N5w2cv9H5DpSL281k2Ty4AkgbFUB6BWo
vmjf0mjxPR8yFnP2Lh+X7K5/oMaJUwyaGx+a0KTSp1GOfY985ecydZ8LEP80hpV8
wwYwRKurdmJ8bqZxRbkMp8zzkVhu6CKafpLtO27Sc0RjWKq1N4vD9Xxs7KDFa1RS
rXfiuyz1ia68Z+/V39RNG4qdjbA7CSs0mVCv+P8c7bx0DpDAq57cISwrCnih+/QG
ROpDZFurWxFQoGBa5G90X82Tza44oaSeZeWLgkyKs2a223DJFQr9JjQNjysoC27q
sEGHS0Miwp0m0SQmguFY0+Fvab3/yplEP/gUb9RsGENA3d1byEl1v1PEQmNiiFQa
1MceyOBLn4918BMJdQWF92uTbY4un+PQXz+1eGTo1CvqNNDpeYdnwBjW7qlGpuFx
k/DCYjzLGLfePxxm0N/KcydeoKJ8GEbMsslWSjtvI037YTVflHou3TueKrFpc7Dj
+aObz+7VC2hJgKZaPfVKD9TZyMky7V5eAvZO/vkxbvsPgaHbKBXTmOk1J7QCLITj
HGpZ3N0FhsH65ywKIV3U4JXopus6S92idy87ONGUP3ZAyXay9Dofjv1PcrVOlEY3
tZHA0B7TW2tWxaIo3/hEI8KXDvQh6RN2iQXwuKdwdxo5zcGoFxRXX5RkEj6m2ecP
vr6nEblC4WPqEtqjuWqi+9okQA5RBBjMBIh8FW8mNwdFK4y2OexuAEoR9vUJ+5mF
NEecrWzoPj/7+nDS8wHr25f3GgppuINOylupPTlwtKNrbrVbzoBEoHchkDWbJvsu
zsy9svMEgpeLxjbkxLo3UGHEVTCtoutaX0pn3i4LqjWKZyFnvT7hZgivWhoiZdhW
rB2ehiu96acp55BU1PkVZRZ44rr+leL+alZvSccxettNvzqKYsS2e01lC+S1lz3Q
ySZzYohpa9ok8Zxo0a3cFehkWf58niEwKzqbuKhDT13sINqzCYn5QJ0PLvFzqABp
8NQqos63k4yU0yWHnZxRfPkVdmIF1I4xyqZ8jwUgA374kcxrSzV/4IRmbsY14zGC
3917WLCU05Z3ZS2nNfq8EdBlwZ5az2tRhOmmIwBBeZE5IcW2+ngsJkFJ6deyBh6F
+U2t4Ufp+mkkSU2uDFlVL8fQNjCJ7LJWZrxzDhEeF3I5aU4wefh/h6gOGhy04HtA
bGaws2FUL/dobvFeSh8fRZzobRIZBT55DCdT2xZzwGqUXVgbXa6WOk6WHqNx+9Yz
x7+Gj5gK/yXtfZKFIQLy5vPA0R1Mm13cHRH56NgjqFzs+IONGK/VgmtnHB+YL+Hs
L3Btt/oBSFBjUArJ4evDIDlrJ1K1W1PbguuwxENRcui97H+PAgK7zyxKr1VQznFA
edkOwKxR6CdCHTqIfmIi9fMMPwazDUmiBPeLxRafCPG/LvJOmS8c3Hx4DGLMt/D+
eusBNUS/UspE0qdmVbmATu/MZ97FpS9oU6EfzWt4NQA2iL4uZhQZqOwWsHKfDgj8
yYZMOAlZl9ow/5+sMixHDTcqJmki17DlN0BxUuiPc9uHdwCSXpBNDLsUOV7pgOqR
4Z1DcxBidntPif5ngTyFEN+zqFAx1I9bT2Len0a3Ghblcb3l0mGPTldPOomIOnpJ
5NPmeMCIcgq3sONdV5u7hdUD3ueuobcCBBPpzTkml9oYLj+5b1i5EGAbEeXHzvhR
F6o0avmGMAzRSnFfPsuM3eDEGyQTJJMCJTNt9wbboRJfUJ5gZM+KahhmsiP2VThb
ItkMfHxV9XXO9K//5fGfixJ+IWx32kZw2KKcNQRcnvsh9OhuO8yQQQMZWLY8un+C
Ib9jjwdBhYobRIXLnUN4qN2KPDdjxrY80ZRKBjNCyaM6ETHYNlNJdU2NwA4W+tKj
bxl5xinlJXAl4hv357AW227XAftGCa8cougL6wvM4Vp26/48T1jFbTJhWxxkUerQ
BotmWHDSCghHjcTotN87v2Ghj6/5MxjzZRUmTkA0dbUyg8NPOh8+8EuY45a3lf9W
JDRTyKeb+uCdobNZz6brfVdPVRqHzQ8uGKzOS5FtgQzLQL3Os+Zp0jXcJXjDwwrN
d+WpL/WADpzLvrcFndL4WsB3b72d8rnpTxldOJX4N0gf2g5Qzio1Bet8GLUIEvO4
FmRFoupAeyzAGrJrygiN9IdxQCQYoLz2k736ac1FRcZOz4TeF+TkJ+xQjqHm2BrQ
RGLf5Nfza57mfa1XGRG5gKSktjws+Enlf2OmZJFMbF+gTudOphn1uwMWX3mHHVpZ
0xnyS7vcuD82yeH9H5v19nzUFR9QHKLp0eftoqema9+/rH7pcsk17DTCflRoJoC4
VoJCQ42PYDtnbYsabf29N0Iiouj3KIAysjbFWXC4y69FgYf1/B3lOxDNQ1vXUrC9
XPh6OYG2a3ytaAzG+crAZ/WPw63Z1qnHCoqR1Tha+Wbbf51la8dSweKjV2t8BrP0
nIsUp03nEcnoRb/0JE0ssei20vdC9Q4w4mIReP+Gdig11YwYiRsO1ETeOK8ossAp
jAwJnyl9BH5xz0pNdsUxXO78zkMuqDLFgJO2vsZzPzha1wuEgmumXgJbJiKjBlGt
HJJ339wrzOapmP9Kjg59soI5v65JDjLiUnmi+62zLDSf5P8+KO1FJn9vXmG0aA2u
8TlXduPjCF72QmDexsaVFteksljhbxAl50UXLc2YeWd8VIrKVJZErqEuJ1BNrovH
QkAOOc4ottUxqo7u4vso9Lt8HR0yR3DTeZoVjok7yw1S/YaEKPXMvnb7vm2vgIbp
DLqVZChRd5NBQHkSzuzSNIpMLjjS92akvSc1/B6ZtuYEdsg+OpVJFK84ZjyuE8zX
EtEfmBeHagWqNE/RI3+39ZZJU5dqJVX0gIXteTdx/eGMlo+JnaXMfuqe727yqzCR
JNGgP0vS09zErEW5sEM9Rz4byWPA9vN5JslZ8aU92zwAr72nIq0z1B8z0iVS7YiB
Q8w7y3EoVnVbVJsA46MBE2rCNlRU3bVyjSEiHKthRs1C+2HvvLi6Oh2oPIbquaRK
wvyPFLRGlQEBBZhiTdLFAXIJvvMBVjomjO7L5WkNUZP6Bjerop5SXoQLo0K5Cu+h
qfF9MWeHNsXOFo7xFmU5TevyI7OZiNmxES/CE8KicEM3ciFMU9MtXu0NrbM1uzqD
zUUP75efXfMdKQhr0mbSsutyTCLorXgaJIHqyrQyJj0LJLk/VCLw4NV8zUL9nAaL
c5AJ+9zDNarP00BMfXfwa9OXQlmGpwAQecHGyn4KyCYfFmG3ViAIG0FDB3rT4n4c
DEH8XgsbCK2XxrxI5o/MteCTvLa+eaf2XtQYRURb0wOScABAEVoJN65gpGvc/64N
CUJ4MUveN5SXvmdu/hUMvTwxkFRNJiHJKNysvhmVj0Rdxp9MUEoF1NdGGPePQVO9
E0zAFUK50BytPZGHU9jna9XtXG58FtmKon0cUFhup8UiGW7edVI0WnwgYhSMtbNr
G22AaLa0iMg4/dwGzEgu3020IiO10Uxgb/3rl92LjoG9zHnPrdEi3eIsphP4ny7b
i6pNUIP6++peR8Sp+CvvxrukMaBEGF8yvncpmZL5Eax3cafPes6UVWOIFvGpolKc
JKokmo5LSi9Bdk+OH3j2r5UMqXkQY21jT8t8IK1ARnvfWesE5LstwYPITeh4+U7K
CBKmbl7nKYeOYzxndUnqp63ji1FNDkozy0snSBpCWyFzRJyqJs/OLoYieAbYekvE
4L78uQ0SadmZZVy4Y9VSD6ly1KRikWRlFpgFMD6W4hhssdw9G28C2rcl61XE5HTl
y86b0uC1pVmv1iVdHSGin1gD/wdRE9cKNPcpQ4S6aPi89VZUi9wuqh/KFV0rUifT
zvnVhv919zmRdnCdZI6weBdjKFNSV6jlBS6cklCMYHbt2KXXRknxz9DPIfIUU5u2
4eUkjdG5ciQxvzYtzU+fW3q0Vrep+bnNH01ShxpWLIuVWFGYMLuKMRKgYLiy/SjC
xrqsa/4MGohxKN0WH6M+Wj+jZN3/KRqWXPnaI8Oh4aketa8vtYuvVu8F2meFPQ5X
Bcl0Nxr/x3ly6s7NmL9YBA7THAx2lUqjwrQP7Z3NWr3fQr06KDK9xLILONqLkak0
vBLuHq4JQMvpyZmsbEFrOvdSYJHY02lLJdCWS52PxXjsXc2r2awG8VD7jJldAgeV
qk0t5/fuOLByCtjgvfHSZHQVa/KPXgAP+J29PvF/cATQ+ivWxAI7rAsfwaUrlwVw
WNbbCh5MQN35BIQgvhOiv8gPeL4bZpI2a2gZNY0cpGBOmlHgacQlWjB/mh7xlikF
+bZRL2XYdehJo5ELUVsuqNoxT/kfvYoeSIfScuaQ4VcX1x52q0vWb4lJYMoleQHz
jtLHQ8n7ALlqYg9/KzGaHz3v3sKD2KhV7bLujYPutwzS1hTYyghz52vgqrcFr/nu
ijtu34mFNeHKBRFQKvk7PZFg9VPFSO6G08J6Ts5XJn8yoyoart+IywEua4DBmxpy
TBIVjudAx2oEj630YUzhoHgauz5hst9nIFZNhD8/ITEi0a1vNl4krkxGkNvgz8GR
SIuPZa7fxKZzvqt0BYEUwuADtZUKKmt/qfU5cg5VLJPGlQ2a1SSy4pyNIPcITcnf
xxC5dQW/VbtgoJ4dvB0QqKIUsPwO5Nf9fUNVUm0Zn88+t1BDy8hx2NWGr4zof6v+
qp5/z1974JCXRcELLMmXWwZU8sO0fytj0U//3GOjiqfeeW0rStns1GI/AH80e3v2
bp6Bpb2UqHfloxtjdgX0w9cr+Gx4UNBhZfKfEjNdgoSt1ySjVkszcJIVXVuh/Pnm
Acflni/Zud92vCJeYkelWlggJAKwBBL4e/Dvt8dh7bxnJmdkn/y8ULbuNNlwwkd/
N1YcWAX4MAtITVaWV9WxRmX4XCw6N18dAxIKu9FOfSnIIpuRrOW6It8FlKLUPhrZ
3dLSriepcMicJXqz/vEcHO0S2s7dD6HfpQGubpz+/KmDdXZflFVtIomXYvwdRrBk
wkuu1A/rZArz6ANL39LJ994HdarccY6acBKfMJxv7p46XOVw2HcpCPBlSk0VPJTp
liiAYGDk7g7uBjB2/tc1I4greKxCNnxSXD1vLbdrkPgm+f+7XRBY26rJ2d7saFRi
eLPQ9wOjL55FqQoTlvOf7B2mdOU/yEnOsLkNRyhSBsfaLQ2m+XAhYFfX7bdwBM6/
gqE+giL/ED5BJg7tsXRg0fMS/pSCMH5qlx/ZqXP86hu9owXAyc0KyK5tWjSyoxpY
nkctgGv2L5nG6vg6Y3lLAdQVfMQsUCy+ngG9NuThQYw=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d/HawL/5DzCdFJhNp1l1/nTO05C5FAOi2/g2t9iopBOLBKlNeP7eBg0KpR7fePw9
HNxWouE7TsHr8zo8/zTm2W3nmNen1EQRBjbxVmqt5+z7DbRQFuy/jIZ7xOJLH+rS
t1JqyQxUNoanwXv2jLnDA0A71noMGGXm8H9a9G3FPzQdSFJi9+pLOFHhipdDKlg8
/abxDQgw68iLm0LuV+3AreO3AjuCOhO6F3z2VlVHtX3HYBpa6m7k5Ale25DoTmtT
hniU+uMMcCrt1x1qXKiFNWwtEOjPfM/c3g8BDNCLrSJ15i/J9WtblaaZXM2DQxtb
nEBHQDndY9+WD5l5hSTXy9gukwHOUp8u7lWyqQYlZNmjsmEVA0GHl9xadR4OsXco
SvkeUv3OIbJLePPHBd8YQ/MZPSj9BdgegYyFpY+/GMa7oMfcgbxzg2LO0uiq9Kfo
oUk+Aek7Vh5tbSnNA2c74eBIh80JKCxxB83T5Gab4eNGTsbCHpz7ukN68uW0+Q72
seuU7TeBGaSaQIxIKGM+SXFwVaaLB/mNJFaqRCCw2vOUYOyz3bovr3/OJz/jlxk9
iAJoAVUFxO6UWHb4vb/HbD2DfcG2idmVA6qojk/hhIvNlshm+5+/6okbqX03Is5q
fquzXQOXCoVq8C9s7lsztpnb9xKLUX9rhYn72+yKXc9kr0gn8nH/KIjZkeDkkFao
WGuqaid/k961zInnp2RMtVyO6qlXJamNIIEhy6OdwK3+tGFYyrY8Baev4xE7lTKt
uk0+ZfA5oSEjQuudG96cokvsioE44QmYmJK2m9XsPrx1JSpDJNII9wEJkv3EdjXu
+sUodoA7dVihq6gB7u4F9fkzPu02Go77RHdPl6sryL+Im0LvYFMKKulHl/vsVHO1
iV6QchltUVKGWJNw1V3cOQ8xKbmBs1aCbPHNTVfnFjyIj1KNl+tF2GqDa8PfKtIX
aM3W0PfH7PRjzuHewDpaj6McyJpwB+BgHOzpx230dW8t82+K5/RZias2S/TM99IY
nqC+UT9imsOgJCd+kv2W53BKiM+uLf2rkiFd/QiayqS8K9cJZefXa9kegWp8b71S
J+sVywSxYOrmN0EMktsk+6wwY14hKHG3RbauHY+tu9d0k+7blQt8uxascwhpmTtR
w1hGK2CDSQ0oYwmGpMBQVWqRzXARzyguF0x2Kq11ZwZMqxcr+CZTAcjhl9vN7jZH
UNSVmdDOBKl3hGekdSVO7SZOXHmuCRsTRtnajZjfazItgqhnljUC61bzqfTBd0hq
PcdhDDxRKMRaRNnk/rXYA6z1GRlPBJs//kJL3kNKQigvnB5mAqe2QarRSJvJGELk
oXmPwHNRjqJ2J+wLif9EVknDUi2wEW/8u5OnzFV2BzsYn7ieGPzqwnDzhilPdg+I
BxqMiv2+Y7f3kIG2/8xCEHuouLuh/ZtCI7ABL403J6n1qgUfyh/ZNme2L0ubQKJg
fwVYY1iejzfN9UyrGJWOiVsEhKSZ0WF24ROLlahY+PW7vBkYQcgfQlLiukrBNhEl
XNEPkZV5A0pcjMvefvB8YEXKeGZbEjk/UEPjSVgXJnlbclUDWMvyM/SYGJ4b1ZTx
kddZRZhWkCGwYzkMmlQO2c8iNzF+JYNx/0oxG+hPkcUPl2ovfo/mPsgVqNSmLdD1
8/xDhRmH6RbdAXXxLxGh9wtu85+kRKdH2OJTQ5QRPjWOeLlSFqV5ykRvqsjU4Dpl
Q1UKfIUJcIZ1eeyKoDnKZp1KDbs7BY9wRVQHZAnpnf9bZdlEgAi4LWXtH98oCVDr
QEVOvwuXAdwWEYsl3owmUZ09gsRHYZNp3bDo0MG5RZI2Xt+5hbjf9AemTxhbMlXV
ySp6BeY/Rf0NhlM5O8Ry7hX07vuIyG/3lrtHbe2hnJdJaARLBdRzgfZKPEkiXcSD
DE5LpNmgy0C8TpcSgO+3ozR3N4p4et6g/qcxul+r46QdZ2Glqile6G5hkFW7Lbh9
evCHNn91oxts6tfzZEGnBI0/SSGeW/1id6lb0z8dK3b/KbNquHp2tj/FlAL59XO2
rwKq4kWZuglVk82ACWxp1H/WD2UpM1M8w+JkccopxjfipdL+fQQU0Au9YkhtRyfM
gJ6oJc4w5vIDr+PwQB4ReVTmk/S+Bmvn4gepm0pKv2WrTeu4KB6r22nuLj1KAVCD
ZtrHga1yHKB6uWdGr4Bwzeh9N8szRWoMd9td1QfDlCwveT6pYKGhrUnteJgD3yU1
K2CSBdAItR8YUwwW+RcFwvKGDTijwtFfgc5XXlupa8gU1uOtQs0ZqVdox72OeKSj
vYGAm7f0iOFna3jVKO+aZIZA/0hKhdWtn1AFe44v8bM7cY8RFqoWG9+SkxU0r6Jh
EZ5UeaFw8BZecS1lZcHPhD1Bc45XI+rIDYHugwq9xp3L4YDMjPlg8PT1+Sjn1aEK
lwxTcTGWjK8D1Ppeq+ESAR/qAap6imEvUx2iwLi8KguB1Hw1WdXkbvObZTxc/24x
Te6/pd2mNr67maz8Ze/Uc/AeT0y5jPOxfBqAOjztstJjTpjtfsxzKzSge5/VfPiR
89UhZ92jcC9ajn/5SZIO1vdpK0uUrNZAhVEce/cOJdHmfnUaYjXqL8/wYblOF6Wr
J6Zmb+7+YsCsnQFv8xIBsw==
`protect END_PROTECTED

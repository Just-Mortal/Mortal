`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
92SlEUutia78RwLexeKu1LSyp5to1fgIpyzTxQozJn0pF76QvqM7aR+s78XC4JXb
liv89j0JNepsBzfnxSb0xw2Ccuxvlls8eMPsF81RSZAEkd5ow90PHDuWtj8+EeA2
62QTC+a8CFwFvaFLGGCCX59IgJhlAvbPLmxJXhes8I+KhPqVRqPlPlXQp03sek8D
55BqYpNQ53XCwooU5isSo0yvIqehzEtu3qrRCq6nfqTXcn3WwOfEm//wg9RRcX1j
Zf+slQpSuhy3FUsuLGUGO1L3t6pXdkrFu0tPhWHbZom1O73AjvdnBU8RlDMnlqKQ
P2YWpSOX5RA1KCoydf0Vpnhxnid0M+GJqxD8D87Trk+6mKrZmB+R5/ThQQB0S11x
OjA6Rv9KYpY5x/NKKfjNLmrAj6b9vFbb1oWlPIS6+VBecUZ4RR7IOjJFYZzpNQ7A
V15x3biflLyksFCJ3Vm8+sAsislwd5TLTF2wKEkcPbHanKePtFX58YwNJT3oBDUt
rQXHEiA+zESSRy9oLTkvVoCVSLSsIX4t2V4qZfMAleZFnXq63HXavMW28Pqaed3I
18LE2Clqh2rkMjAfz92ua7OAqrr0l04wm+pPD+E+/rRLse5+PpQub9SwCDtSiR3W
My/vL7NvwA9EiEGZ/5YUa7Aoxk5ffB+obdVwRxVFyid3mNrPWU/UiJtpCgx7VvWn
IqxuZB42fByHM5AP6j0mAiatIC61UoD5Nbt2V0GDEZIND4o9/yvVHVyCdj+ceot/
alZMygYlJdzuvfUPmZtW1sQToamPeuQr1SEHJjg49gJEIZ4uZLYHzzC08FsEs+aa
fcHQIQRh1WamUf0bGGoaHoOcHOnAkvBvjUDqpgnSHZDGhPAO0bQdSFNpEUI1cwb/
AvVx98eKwArd6uycd0YbCLHeKJ0YXrW/0o3JcUrG0LQXTBeDAxafhjx22rnH+DHx
TzgUc4JS5G/T2BJcTTZoaGMcRVKei861DB4OXDg6C7Sv1wHUAB8vyVrhTEbWGoyT
/hqiqTxvvdcwDI+8ypyZPhcOggDJ2ASfirosW3/sE44R/mu5eLN1xl8xuXfSIdP/
OYXVKztI+fWxXxJjjFSq/GQ5MvO+230FIwr1OFszLo6UjhbDr7+k0riSXXLqFrem
3si4jWdBKh8lXQ4X0yLuSWyB5GvXfi7cASbV1UVDTTgk14R7oOs2whi1q/LRovzR
SWNzMWESyu5NHq2iYYUB4ATk692ZsNWTgQdQ9Tjudcb3JxtHBxwbUW5QdFrRrTbN
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SdDPmGOXbjHy16Vavf0p1MV6Y3YwC39xlDSBk8th+9NvhPhQfmjw4/lfDwmqn2IJ
NPOdXFSWyAbH99RjmdUTa9nGMYRLW/Gyw9L6Ox7FzTv9rfHJij5T36SFRL0Spsr0
4vbE5t0LuuSsMAaf55c6McsSFUgY2u07mAJTSZZmPLIXzznqG3T/rgJmdGLiFE+b
oEBuUbJcddGBhEj7xfjFJWAG1/YfEdfLA3tyFj11lnaFYXp/cXIMKOeprPRFveWb
fbpy0VTR9l/BNg1SNbVIkGl7f5ZMjKUrdh3QfsXQU8m56HXIHDkUN+akLZvjjiBP
sN3VcqcOwZ1jpLE7xMKEY65xnCqANXaRqWpGbO0fNB4c7ywwHv4aoZI9NjJGfE8K
lDdiiFnG2kMflHovfBWhEobTSDLlkxo2q9kzomrr/W7MH/nmDbSRZ9T1YckZEY+c
Z7GNCFjjgHlxn9f8MyPFjkBkO7smQ/JUxVmr566xfIRjLR+YjTMOJ2qznDtY022f
BIY81Th7eFEyLewClqt2ITMjfNLO5N1atQGnHJMcjZVW9zE9wAdCH1v8yhOM4I5b
F1mJ1qVKfzfE5RTes1mBzD0fWNRF2Urvb6Myg0s5+xQeGjcqdBYaSLJP/Kh8552b
7jUDuMFKRYOvGtuLmnvxItJbAdGnYaw+PfP8/aOmu1iRB1DP4wQt2iDVYNqkdgZg
JvZWCibF3RmcWTifLx7wBEWHQz41vI5lFl+XtbHHneiko5U563b/XotBjg6uBau/
6T3NMwgs0F/PXkTKUpDrvXaf4LvGmNXuMCHuCJlqYbKQvgr1g/+cZCVE6MnNGlC1
f8R4JI5jSLLol6iPOY9+Basczqy2FtV6uZDCtWiJQ9+oCyr66RdfzShwO0Hu/Kyy
YUdX7YlKjL7nxElZEgAeCGX4B6LlYO0+wiFgYj+5GCGm5E6/PCHKFxVXIvGCgnl6
Jn4FxfH+af9jzpYEBUZzN7InmN7k/1SCOYw+1Z4gYCxLybnmuVbxMSO4od8TIDon
XBgxiwema9+Zkw3RIsOUWcXNSzr8ADft7EMVXFHU+VSwjxBtiE85Xlu40VmWZB1l
a2Joe6yMkB80fGJBSeDX2gWHFX/QH8n6wYkMdMF5Fu1SXrec7HrV3KbrfXuJ86UT
Ibif94OUeocyMhAirAO346EhQ+mYY/aCQu4oTmaaXalbpHCNcM34gGvXg96XIRjQ
e2Ok0ARxHOQ2QsIhJAuSMWnszKDX2Ai9+X1FKyVYTjVvr3ykkWbtTsbuJMQZt0jH
dc76OnBJ+8xpNkb16SYZQkBww7KwTx5hNE/Fk76TywetTIfLs+DTxrcUmUtfZJ5B
cjDtcvECaWpFjNY3utVZaHeyxIZtSBwVlMTaywmPTtTd+Mp/NkaWzotqJBFvIQqj
JoN4oXOY9AJEYoPELjvUR+LeiMyVevWBp+5fQf4MT0QWXeAGfIVuwnF1a4+t3+ue
PwBIo1EzwKsvdHAGXgvR5c5WXx+QkuwrdAc1pyavnyIF/+CwIHvClO6yx5kKKD66
+N9qI6z1QCVux/S+Pz2Awfx/43oKvfAJBdOL2CuS8KnZrjFM5Cr+r14l617qowLz
+8UAEf4vLlkU4n+VlKC2/QR4XNBH/KtejEkE+wu7xPimhPrj4YZLRZmCmFMy+DcE
VvQD2auSjHEcZr3rWQUtTuBUqd2xNZ9pbaYt7bjyfpjmaa1EnvotGcfDofecMQB5
s4lTrTF6s+YcIxPCYW+htjVjui2Zbo0kKa2oIEKSro8iTSUXpweoZWwe26PzZw1/
LIR2bjpadI0jiAYPgkQ6vvfFm+jOUnzo06YUdyxS84M3fx+N/0paY83qMLnXMGAE
DMpAUjK7wyWOm9RkIk5NAopUJNMQ/GXrAiTZ8UcHSe0u4JYxKkQKOM3LiS7aGOOw
rqZPV4JBY5J14F8TNXzfwmpjq/508/5IU7hkMQnIy/j6FKUD+jrqP4hB2M16oFAn
eJDNKoA+8xiaXSxyrOmcgJsxahlpyOx7i+nY/F8xCLFa41U1j+C1blyAnv9k9jbL
pZA1Ai5mFFY1IEEqX13C3P5r0QQfAWf5L2oQEt2VuL5STxcZuU12BwUL5CqWcXnB
Pffh0R74KFR/oAC7irFl9qjgpSSWK04oV2edBztcPYPraPz/4Tl5QlT/kVzrU0vL
+5don3Mvfxi5nEhBlEpeE3Y+5ydjTxnF5t+caJURqZLei27zdkHsjkgOAjSGyNgz
kAN3b67M/Ur/PzQVQyzESUsEUtq2in39W0TxD9tOw/DYKVXZ9K1Hm1+NraoP1biH
5iyGo6sEzp01xP0HT72GBpPTvaWscj09oMIDwVn3KKg+WKR88a80gHmSlY6HMSHq
ygEzYYZW6kyoSf5NGs/duitk1odjZRenDCFpS+LO9nRI6RMEQv4rqFPew8ioLlNj
cw5g6wEYlClcDv2gpnNaxObkc734pQHfnd/Io9E7FOibaa7wCcne3oNqSgxX76t2
Fq4RHHocZP7mjybV8HVznTruLJUibC1aqotX4rJyvGZS4xMIdxqf0EP2M8CM18Gy
hAWvBNvrymEJYe/iIlA5DIp6nNqXwC8pK2skA1O/MNAJLQ9G0BR9z6gYwDJPCIRk
juhhYPeYmnlgrIw+wN9uyvzMvaEE8ts4Nb3yXBQCtnT07A4K9FhA6K4WgLDK9+/w
RP0coa+OU2MVrdsFZ1SF0xTSkF1M8yBxs/MelylQVWlJKN/Ql/jfzMdUz1fE6WtI
2dYLhEB1bqKTuYHSqBLxJJ4oaRwkPrRWiOIJOWWxByOiO8aeu+NnWI+ZTulkA2gI
sRGDgSWk44Hr6rJ4WQIgw2q6dV8jkbqizJ34ZKW/JsP/TKN8G1AZibOEHk4kkc7S
jo+qeMeYWCRm5/QZy9foOD2QtuPRgEEpULG15wIVNV3ZeIAlxpfs6NYi2yphJNZz
SpIOCqmCKe/f53ByuU9B0vrGDGczH8rai1fGdlvgCWVpzbJy4rjbeQjUP+dZPyIT
FS4IbQZcWTPUrSRKtaTpFmbQfVre5UvZdd+Zt3fg8xFYKZk2kfVjAVhDCkTDP7VP
YVhimlsxNDq3ROnfgz66jPdsnB5nNpOZTy8orRyBdmRTjgd+G8eOWhhrCaJeTEIB
bG2aJkyGOCNuWValP9OfrU6vnTXFdQMJeYiLLx9OLm1c+RRp9G6SG+IXlGqaYUes
LUwNY1ysvDJIJ9i43mU+Uu8fB6/X6kbFkDVsPiLtTzghuiqpkLHz5Cj7ApOrlI30
2TZlduuhFnGo6eBlvF5ruraEGP5eNcGWRme/woxt02KDbCsGvGvVi91R10plOASo
xihRj4D4AcN+swvpYkKBMedVX9wOC8kkweutSkEB98Ei8X0nc/pmZkq8FPknlMBC
7987lEfofGvZr8EXJ24zo8gl+jx6NkNPN4RXAXT4BBth6KKWyO/rOHCl/ix63OLj
XZOiGT2pMvgkwZVlsPVv+G6QtHjjgU98rU1258PhOdmOTXXSXqwgiAiwKVZSA8FC
hRPDbIh0tSm5OLhbw/tdsrR3zNi4rT98+IEb4u/qKaDJuplEkgfPyAkPGymydL73
H0DtnMntkKlJp4OcupTi++wCqO3J9kqEqoB3ENINXvQwMO3iIDK4hXvRLG3k9TZK
U0XTR8rOMvUcMFdupWevibdkOyizicmKahu46DAz41l6QcfvavP/jiaILC/IP4qG
K3KGuwNdJmMBTX1kJN1oZrORRLLmmnOv5Iri5yIL5yGAiWmLduzze0QlXOTwxU46
XKQOuo8V8qZmNHfPsAVrrjVJZxKPI4dwU+1w5gA6AcoAN0uuTw3BwvXuayMs4wFm
5HWD9hM5lmwzf9yB43D7FbhJiTOdNBSlYsDUvRV9MjOvKJbIlT47ZOeJUJHgizsf
YsvaJukyxE23+b4d/Km/qKNwyFE5troHkVeYnKf6UrxX5RvR1DEufWg/96Ke1unc
SzOV38Th4ZiLe5dUV6bSdLOcmUn9CiwZBWAdB7p2vlVOZ0NlRM/hfWkt1LRRpiDM
hPFTqopM7TtsBKa2mndrLrwi1IaDAMFevOupGF81UTMVZqFKsvJejVpsOyFf/0/E
8iDx3y5SX7E8QaRrcqxnwv27HTY9dLQkHs59rvfOmxNU92ONMCWR/tNQzDK7eUYS
PtbmznvqAgz14BFGRj5ttOJGbDgyFW7Za+U7sBlHsYV4smCBjR40Kzh8mZ15+cRC
Nqrmyu1Pk3rg5++6TbJc+08Xl0+RPE4xC1B7ZdaWjpvN3X9lHGHJex054mvx1Teo
V1hLRsyqawSc0P6LKP6SEFqYMVTQ0votqSUylW74Iyc7rs/c4RheTAARF9M8L9Fu
ydrkFBzW6VNQ8ek863PWjTZGBUS4TumOPkXZ1xrIM4zOgXnPAva5SeLIbsZUkjUV
MlkIqGFP0tOkoHWrI07IETabXhUJ2XGquBKuYrm4N7bcaEbZ4T81KLwmOwO+YthG
/sclafZ96cIRQk9ZY48MWF3IEp0mG/QAVX58b+PgA1xTZVvbvVY/mOznoHxNEfZh
pv7IcH1giBYwNdCSnyartQhH1+1GvBcLuIshH1sDEBtMEOHsNFZmyurSYptaf1Vs
LuR76URCbfiUNBgB/NJwivYzN9qR+/LoNHfjY/yjVVEReOavFS1WLTw/7X1ftQul
UmziJ6YeMzT/fEoXhsnh70OTwX014b4BPz4EXQYa88RsXyiYto1maiiBA6ka505R
LnVE9Oj2kLQGGkqunU+vH5IDWdxX1Ts9dF14YjOyCmd0kIxUF++Aog5wV47OuR3E
3c9y3bjq+MW9zEIsvmtXjIc5jbcIBTxhTtnN2Bojn1FGUIU21GCl0/ng+EAiZCII
AP5wAApFkfeS7gA3ebuVLWKjmP0vfLfql2AxxB8zpfzerLu/+MqRIfbDB1EIDu9G
xulKjqAVeqamxXC15AkmOZrl/cRNzkpuQ8wYqvl8JfY54m1ymoemolHiZwCVOLsy
QWDIA91BO/pLmQxVMFtSGw0bKJs8OZKFLu8tPyiz0o8lhEWifG50Vv0vP5gQpSZi
QabZZz03KonjRdybBOKl1nAwlapXijLyKWIVlfRIWhTKbR7pJNNfssfe/NkehEBB
weRySz9CpaLy3xaBa5LK8ldx6aew6yc7I4Q6NqjLaW8dewN+Ltny5UGxMdTC0OAS
wmIHzHDvHRyUTlJea9k2Tfv3OqHgjQ7itEZihf7mT+6x9GeCtpfIodiqyyZ0ELzo
DVXo/LDjm/YkeVMFQLiJ/+9FBVjaQm3Btvku+ygb9MfFlpT1ZEE2+s6ns9mG9Ymc
qtEkPLcLjQlbKeFfziWAcmksx9eTQMXx2uq2g/SahqMkAH3oR3yiJzD3+Zz0mMQl
UtxkOinjA+RjI0rMw3opXPY3uiA3fTAtfEPfs/EWtyS7vLUALQ/NyEmfXhaJa2Rr
a9Vlq0HGILuFdMerxa30XO4ZJgcA9EOZ5Zkb893z6qIprM1BdmnIRekJ+9G+jmle
oOURWbRZe2OdSkn6BYkdgJlLHQIpmEaj+feeJ+h3yz1pUhPYrc4BL7biurnZUU+1
OcKnA8kY6KsXHviIg75giuWMtKbcYVp6sH2ZXE2GazOY9+qH4IerqhPBNp7TRXHR
qlkqkDxJ+4uFa8aocPRWBo4xHyG/X8cLXIiVq7AqfEn5jPOETMzOtk949sZIDF5H
WD2/cqcJh3scYK8jm364NGh4mWKRCrr7QpmCaV3qhpgCXon/t6UdS8m1b4Lu85Sa
W2CebMSnut3kySReSmcjugWQtjMQXlOSxGVCsQaPaoo1XDGvdyJijZLM8KBTZWhY
7hItyLcHl7sbpKywYR/WoDU/3zmdVtL4FlNdI+IxuVvJ1nJbR2zRLeeBvah/aSnP
pj09gog9PPcEKdHTLEhEQKMXb0zpYBsXVYMi3oPCoKdkT5XyE0G6sYZPk1fw5I/l
1yx91plxmjxFspxQ2ucerygl3V5XzScYhzMaVyxrjp5gZw/AiIuI5E4dUsKFkWc2
S3ZYLgCXMf5gUXTPf6wkNVC4fllTO81vS3JdtNWxj5zwUnFGhrCpF2WF2gNmNwMH
Zly62G7vQWehvgvefPRL4bYkhkT1swuXV/Av+OR7Sakf/l4MeUDqpIV27+PwF35J
/ad/rqh8MBP+dWaHbya4KrZY8BZq0F3nD7ZEBx5Jy/xBRl+/n8OwUZaSuRLyin2T
RafQbMLObm9Ao5z+rB0i3PzNVrTmZ3BX/loU+v1IjzwxUXsWd2WGt05AekW+MlNV
lKwWl0YvW0O9TGNDxozHEA1rDpo8CNllZZczORpe0BYO9BbFEBg8RlZTqPnrY9Xs
Pf0JJ7ZqvK44UPEJDr/bqxUMrrrgIt0CqWP/PkCuhN0GsAR3VhSQDLGZcZ1+wTMW
mcWRzZOAcEL6FPSnknsjnhzfCVUmSILkiZD+X82yaw4uTNSIuJUWFHIz2HhN17mo
ekGfpEc1pL83ZCV57PTdCB1s115DYjMk9qLxa0rstUpklRQyoGI2JcCgW8ldhY1q
IumQPdLoRM0r+Z8cbQco/1Z2++4uhCKXfTfHDAB+gj4I34nLsUe4/Mt51DW0gLyD
xXmnjh7d0FQyeEItC1goEuFrkDmL65ySON+k/L3fMH6Oo5WvVg+VreMm/dYD3ZGx
siF4GjeBlmWg6my6ud+1mnbsoORS3UxtfX/2fQ7tGDeYT1c6ol88YlfURtdh8rxs
Yb/d10OJYwL+akOPqEihFWAepC6Pt0F+jOqfK57Ua5P794U/Xj4zPM71NkXOLsvU
pCKzU5+dOV0PhM4k7uK4WB0hUYxTcZBnME6kC8YWcsHHHTbcR8/HZmfKJA8dyFph
Wjz//t2h5L6uSqgqA4YJmX4f1vgT96c6S69+sCFI3ErwT/+JQyMXYg6by44yu8qy
DJXeb1qSkgeeeYSQogYZn95qxYpXs9z0WcChsB/NQ+xTZNzvYwnP2/4Djskj/GVK
1upF8WRWs4MNFSJKwpNspkiOOLBMsWKJpmD7ic8agB2bK6NOFdlxE/5dkbiB5Ebk
v27euxgvygMZXEwcYPSiOPjCyP6rL6Icdz5zHedLiY/vBcBVEoPnoiQvOVxMXgb4
KsWDWY3YmVSh4nAyDr9zlDn0j77SG/2qUXlnKEhY2ElUr8C/DMlAKbXbhTScfv/v
8u+UFfAad9ORO+gcy/s7i1vqsFRD+/cWfkhnxVeT/3Ck22dhOKJYd4+Bd5uEM+7x
uk9BLliBlY4vATZl9aQV4NXbuVVDGY0pyZbW+zSQowHRwX7r/kWiVob5r+k5tLsj
tf/2NS1k7vmYFhumZmi54RsD0waMD6ecn2EPLfer/QyvQ5aUKUNaPcW61/vOwvLC
9U3nIf2h8j8pxG39ycjEJnPAYpjVYw9SYH14rWfhdgeVuX/8Zc/tzqrX4fVdm7MC
vf9daMt2xW8LP1z20Ye2l6sa25v7uxCRbztRNWWY1ZLUUwnOQMNnwob3fFnehQf7
UBmJdGHEr4SQSa6Mad7m8sLXM7kNZWWKQgmxUjKOdmBwocl6f4MdJA/Y5iuBX90c
aP9IEgic4ZEGFEE6OEOhN3YeX4dtFtpfUeqXsOGMVBlHke5AXULv56Fm1ks9M/dy
pUHYktlmOJcDw1YrEuRbbQhYvPs/kU3Ncpo5kaz26RPlcaPGk520B2k/USpG2luz
EcQEiRwrw9C4cC9e9Ja/JtrxGX+Q+ucZKinIWiO57TRl/Tq2eyTdplb0jIFocAtc
cwxW7ivcYQYTV3vfrO3kMqYsSMcZkwyvJa50vRzZayGSsp2qdunvlCQEMmtGcWhS
bk9RXoTg4wpj3qPI8DDs+XsUl9izPox8/2+20PmRuwlcQMFIE07GznHZoHDcMl38
6DA560vJw9RmJL68z+1fbI9VbMHYElKSC+XJUF4bk2ecE9wj3UTJEfxD3XT+Himq
KcxFi8MdAPS69/lN0sfzp3h9WNq6SNJsxHT5Z30uYVu7CG5fUklJ5DsMDG1XNOeU
g4fI+OPy9MMv91zxjXtALx87mVEQ9uAhGClwYutq5aOdsq64sCpVdF3Ai1A6BW7R
UsT2CWNx4/hidKba5u87EoxY2DWZ6l43v+icOy2xcF6Q5fsjPi32wK7487XxJTq8
id7gS+qeenzp9gwTa0baXRlpDTNZbUrhRAE4EM2SHadpvHaWKr0YRFXhkHYICN+/
YfDD/BaCJ7FjJND2P3C/BhnOuKeTNK71bPCTswYZaBtR8ZIza5frdC2e01dvIRgj
tamvT+bK+ufcAz3oxPoW1H/e3t2tcb0TB/pXMtf2P64ERrK5iCOFRZ3jTnHBH0oF
OSIyCfBs/eXkKXqyaYgmDv02klZG1HiEMxsjKDnS++ju51ePYlvFOff7FZOgSvv7
4Fslc5lk0YiAUo/1PDCysrd5+Eiwd8IC95j3AkWqWjPurYQuAHsaoWCc3TM1kobA
+W3fWP76bEwcsIEFEklUtzFqb1+kIM47e4Jj01IcTwIMSIA/0Zs+Y1+kxS/4bS3k
qlF/obbR8X05tukQ0iV9EJECI/NFcTuelVt9izN/2MaMbeHeQulPBmN1RAfw/dAD
Ptri3EkdoMERhHfp/5oTa6bYwZWAnXoVPl+cCqU+uDutG7o5mX8fI2e09vCXzbIq
SEeslPoSjCXyaJ3/WHNRu7bUBhbIRiOCMwEmb3vPsbzRkjVQRnSSVkstIQBAfByl
VKseDEFJMx0OInAhEF4Tz4q08TVxUpf8Ga91cbhkNGWiFyMDcVP2LhB6n+YkmnXm
5+mm8OG46eQf0puFQz/gJHorwO97OWejpSyWkuc2ANcO215/eGHPbsXt5ZipysGE
i5yuUxzIpOMkJSJXxIuzcdQ0FiwSFKqs3rVC2xy2NVK2+h2+zXq+qIHNESvlrd1R
0PQ4FFsg9q8sy1QUuDDWVH69Ssrg5bAETvdaDi+Q/ZJMsWiLFGQu/U5LYI0OV+29
9oomQF3z/eyvbnfcrsSHxcBFiUyxqzcfeBgcwm2eYFC774nd7bs7obOhjLylF3Fl
gKMXoyQ+4j8lA6o8MPZKKQEbSxuHNx4uJxhPMwqo1iMmNSF8LjjBH+Y/8epyFcEw
wjeVl0lesstffpbZq81RjgNqmWtG07UUrd4m+jogYqCKcrJfgW4ceF+4XcACrPip
RHJVfKc+VVff2cTgLaG8fLHFuhBw/FANSgJMXbXmvk1egheQvVVepnXj1ObXyE7a
G8pddABJgmr9KrwJ2nTFjyOpQK94Lt95FkB6hHULSqAdFPriEg0wEEOZ3mnkTJZD
Vd6AvTl3s/GGINcMZ6ti79t77zhaGsO0ZkfAsTYGFDfrObFQB1cPJ/R58qTC3DsQ
bcDxURHECLJb7IeC+mKZTd9yP/UgeCvMPADDKiYDxE4hfQn+JJTJQs8uQGSycnFR
s59yB+zDbWcDLgSXMpVJ1YIazXwkWvbxPXDzYOXHwxrvj7jYnMJfzVCBtlBV4gQC
xKcMkvBKzzWyMaLZo+h0ihLCLc7COtMNcCWaL5VrLh7u3yvRHuCIYXqxYVyxMovx
Ce1tHO2frVlFhbWmnuBBgIA65jr9ocRsmvMNtZvrRfAGHNP+HKDZyyVKXyx/IhR3
r13JcSvGcOhJaOsC5N3NM9bd+ihp5+1D13iaURCMjlCA0baXSPvJ4trQhTF+fEyk
CFkd6A8/Wyi41irn5+C1cJzSTrwuUWiuOkgIgJcvCE2zhNAKTBROrWYx1nvNANHD
NVG0YLIJjKSoNZPYzbbDmCCNFd9w6V2I98xSVP/EcqTuXLzpkQU2F560zAmpta+p
sJCw0bsySXXPS7kkp5AaJ4gnz1BO9Dta1Bi1iTlbuJ8pW8h9nTh5yBcZWv8+sWIz
rjQ16jiod9jrCsWx4a3ciwF8QTx+u0tNASybw0W/GmTb9eVYLFoT65cEq+OlF3Go
MyvB6vTDidnCNnPPQLeqWeDIDHnZr2/StvnGijDhXkmDqXFjPfrxkUdVnVfFFxFE
7GTEqBRGlgjs/mPfqTAMeMkFSyp3h0OcWPRfHxf0mZiVT44j+PN+Eu2Sj+okgIG+
ZhRJf07fctQz7cZIn1beu3p28/n4OYf6NDqBWWUFCLczRgpEoTFwLaIGbwdOvNMN
6q8QiUGLVbmrqMQ6Hl711Hsoyzh94szpqrjfcGoB4dXDY8UNzyaDVVC8XtJjtqw7
LBX0yeXadR6BZ+MQNpnZoFlVh5PyXLXuTjjBwerd8Rt7blW5bmX3RSupnB1lkagI
qmhNrswQydfvGASwaVuVI2nz4KtPkS0ELB6s+JdJhpOHPEorU/eFtn5C1YojNyuL
KMZl14eAZrz+mz359hZdXzOI57HSvvT/b+CRi0+xKDFnx8AtZcAb2oxUYMmG1Tg8
wvUU3oXN4Cw/DL0IvJ1mc8Rly3sJl19FP+jDBusJ34wcMYCIm4jrmoWh7ckJEskx
1tQlP2TNZhHH0j9SJletuDxPdsgp7SWR3l0wOWRUZhkSBm6I9kB7oVAgN4M6PjnC
wFiM7I7sRapEzKEao6Yn3fAGZDZfmIKvIq7lcXfX2JDrLq+U2IDP1O6vvM352QwA
KvBlXiaQZtPWaXjPLPZPPWM/79ufXFV+ECpdhLzUTH8hhZX/+VkAdK/hLPOicVQf
O67ShrQT+XZQTB61UkacIkqYTmwjYt+mh2lRl7ANDHJ3oU6fhboiKzepsGbiHO/+
pJQSW8RchOyoCVVWXOFSHVWjszSGMOff97jqK/zs+d/iKnWFWlhLRj8ogrrCQmda
AoqLnBXoMtsbtPc0fz0u2Q==
`protect END_PROTECTED

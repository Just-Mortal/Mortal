`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tVbH3TD3dFR39nSuYWAB+Uq9tk4GBxghM1dCIk4k7OylZJphkQsXcRCtFXVpvwE
0dqy/6IJsL8CE1/S7pCtS87m1DG+c7beL6O+YrDuLwN+MztkulhkA+nFkeDRjmgE
NG0b7H4oJjx/vOBzYi7wwu7qrbI5YDfvmKU7MJ6UWQ+etJ2WZFLds8b0fgS6HCSQ
Mwj9iZpu89xwR52A7aIbr4n9RWdMA4nrlA1jxYY0DYnzdWxtqqISzuaXDoXzx1y5
2SuP3yYb0g6w9MJyvH1X5kbcVCIbbKx/n6iXIJpLn4P+MhD/5rQgxI/SH8BdKRl+
eGoD4GOivpNlrMnnhNf0kaY06n+8LybJXvQZzNbXRLBXkqFP2VJjtC9d6I0Uo3cp
wfp7K5O5w27XErJ7dXhPuzzhaojFnncNZgNYi5GznkDsSIHUoGEVEnd2YH57SNcD
Wq+O40I+ginq1w+rjjrxF69YPPzfSJVG3o+DRcKocRvSCR4D5v+fo19icaHzF6bE
IB0KqMxXOOKL4hr/9Adpp008gIBPkc7/Z+RwkGfCNvYetSPBM7bNNOr+IeWnmaCQ
/T03G+hiQv379MJyNql44qKEzUD8A7W8DEdSy0XHEtZi7rtngIZv3/yeolLKoEy2
Llk4fXs1YsL2DkNF2pQix6eqtHtupeysqkXmn/o6JxgNKNYKFaHHJ4AiCLjhB3sR
LGnOVtR7lun5YgSmaGM4wZVUuEdjj3SsZlYcRlQE2VvhNG78icPOqwbNNsxJ75LL
tkqva1DYRGo6Nap6XoeVVf4NJsPiraYbWh5nZbRPgUmv3DdFStYDMkEYieSx59WG
1UqtoiCDgd5G0T7ByV5ih3lIZFyehJeA5VMh/4ZX8r8sngUhy/5W3qrBEVOWPDS0
id07kEVpNq1KEPPNjc41ILe57icu63CZLgZus3/DtplN8nESKb5KxZYckuOTtHzC
yUVoL+trHTDr7LwLvCa7yxY7ICnATv6X8kgmdqlNGG/b3zsayOL0OrLhRe1sVfXs
+DgNvR0QQreg9oze03gdR314wfCthoAJDxDEhvGxLML0NjegIF6neXdYqpxESsYX
ss21J//0HgxE5kYOWTZLuXzomKibmSDq1tYB1/Z4RwDyhNT0LJuhgnp0hMOt+Exp
7sM5usBni6iQHgbGvoe/lUARkA4ZY6cTpbA9rjll/snHdW14VvxGXPGT+0IpvmBr
xcScceBLhWNjtQuVYe91zGgsIVSjcBRd5c8LJ/07ob57rrPz7RT34X5jIzAQUN2S
V1BnIyHXpDM2vvQHEs1rctxAmF+xkXqDo8fcB123ymiBBVqin5gq7aP3SOxClnE4
Qg8tOTMUQuos6E2mGftf/91gKICCeyO2PGXd1JswXUmOKO3ayvAO34Y5TBSTE4FG
RPdvhESbU2DXV9R7Tig4SYcZviNkIhdT4JZuyGj0zMNYOwzgBjILFRqkHNZlZd7T
qnirNKcOG6l+WTE2fzO892haBDEOusuyVhOTRcvctM9afgp9CcURbZxYxnKer1x4
BCuf0yzRlDDXm+dJ0s6sUoqpLDnsWq+XTNQMcF6BztDFkOXW75ayjO3dFBjeX/7R
s7qUogEKgG0P/ITQCJI+i8LsVDREZ5FYtvDFobHBjJ0WgCXVqTxd1eP+xRhffUSB
SZEKslowU2aohA5osWQDnMI3pSljvJGYoQgAq7SiPCSKajMjnCuSTwXQHoy8lBZd
xQ2cDgN/N2k6cwZXNyWO5t3oesx//z2gJfocSUC3eipNSV5sPPSIf5S2pZQwHsMT
kHV8aNA6J6BHPALAeGpK+ZkZUgoF41M/TpUjN7Wv4ui88/Qe2DMzjLTR3+paz9rE
`protect END_PROTECTED

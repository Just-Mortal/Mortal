`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sg4CH8R9Mr7iM37H52u4mnKgcQs9m6ZMj8YMHFJL4E8Ke3QS0BKKi8MMTQpg6JxS
DhXRu7qc0tsaLwg1QU2/BdzFge9oEXnfwFzGxF7VaMIbLJHnzCukzITmVhHByHiU
RkZ80L2mMJTIQ5+MiTlZOX+9EF0NxxMCrd3N/ds0l57ZYenq23BAGmj8Lo6CjTAq
83bOR+KoYRZmJRDjPWTX6nMMyAWvs6vTSl8Q84bLbaTj822pKNrSzC8JlERtYxTC
DGMsp93Oauv6R3o1Cc/FteKGKCEHh0IBTb8RlEeqycENBEQdjrb9GC9zQy5csYkg
eAnr9bmc2WxhixhZ5IsGIfKT9GMKW6jBzrwdiGVzc9632cNU3zSf6Cl6j5SCvZrv
CfhYct70OGTzLfUAH5V57E0kDpJhGVC+Aats1R2wVOGXdQTcx/m33TmT+Xi5cCBN
aJPB6PzIzVc8cHvkDpn6A6SKM0YcjyLvuZhoSmBk6hMsEMi5FSxwZKn8NScCGf94
AxrrhDWa936bKmmD2mkY0TS4C2Uejzpb+Ly4+FEq4/Yx9MtwwpRht1LYgFA/QHCu
Zyu4SnelRygmJI+5LOEnlnvK8eBz9+TDxQSSUQcdlhaPHhaDtdXvXM9qMtfr6BmO
D6Fb2pzpZFOZt4cgheejHx/WkHYe2hG1w5z/wKblqQn6jx+3Cpo/n+/cIYTiuUvM
MnC4ABre4zm5dHAQ1k4Hlwr4zekurxoyHUOU3S5KziCq/ue648/vSCeTmI8R4rxi
/FePO3bBCA835H7yuvyb0R1bInDkO0bbkwuRKiBs9E/Nf9dUmtygsMeo0yLjv2Rw
4sPz7aw+dLmSVZLfO1b6dH9lxpqCLzuxdhVhLLRgrXgW39bM7S94tlsmPPMq77u9
XTb8CFRdkzUr7E98K7ZPJZ7ZAi5PfOkYYErGXAsPCItMpm2zYBesCjHFxuIz53ld
Ih7Q50itSacMcCwNFw0+S8Jc6qh5xHb33joZKwHrdLAAOpMmkmDiL6ij8NhmWjiO
wIfRzU72b9nE51RuqpjngULacxXbulqmA6d7v2OkYFRbua0kyrZBIb5h5IIqC3rD
RngSAHYAj9fTVKsgprs2qnABjPo2xmtPMm7z9rpdJfzlsktf4RZKpZRlBfaLbOmB
DaXdM+MCCREAljHOvzV3RVO0CVMcv6yqCIxVP/Q37QeRMF3zTqH68XiptFswCf6N
Zt055uS4mSGi9h73R0JhfA+nzwlHqy2zEmXNTd1bSvbYADNMRKONZmrVDDKseQrz
Xg3rsglMGyWeb9sLlK+Z3zQQIOSK+Vq5shod2R/znIkZpldgQ8Q8zwkTgez1f6yH
Mx3UmcoYK0AFaIejxt/ZogkkvlORjuS/7G1VVsU34Myp3kDe5gEC0joVDdCkZ6SB
HfLWxN6X0uBukLQJohP53Xf4Feb4T65BdFS/Jq0soI1GWD/1YIKQQfrHkVwWefP7
hYdxUeRVDsPhsDGTi71Eh6EdQOxDRiji8JYbGhVsVZRxjgZHeYz2RhgxxeyxSB6W
TApvcgAKYSAcI6L5PfxhSOJjkYlwt+O4pkS+MgJOrJ3MEdamrCTORnE2bF7Ne4Rg
+ht85SzSTI2ES8CWBdsxV9GDjc6ddeR2WXPe0/wvgOlnUdhbsvC5AyblmjSP4fIq
FnZOUuTmGMsx27sNkyLXUZpCALLR38KV2yKrlDpawBdSsRRPyF2uR6tXjzt01Erk
H7dvjEQD3+xBi57PY/+GN4LVXZCr926h7KftJB3H8SA05mKlSQFf39hmwko2OMYJ
Kml7xrSxpnRc9dDXT4hC2OYnoOhbI2FPQxRokY/4ylHPB/rM2QMJUCGFQrn5haKM
+UEELBGeqI8wWKYtA/lF7NpwYQMFvqgMb1tKkoqxmJwClqMnHJRE/gCsOgH1AQJo
zrnbtxEcv5AL9QiCCBdu75nROvlwk9WFkIgD/2Umzhld4GZ8kVbQbfmFk4Ns+BRA
GvKG8DNtiCsfqzhmzkhsMcgvqZKSog2g5tHzL6IEMdra4rZkc4mM0xt1nemq0AQX
C9ITum580w7gsW+hHf2/l+MqTFpiMp9O6Adbw9pmExJsO9XHTAsd23V4o0lGn0lE
1N9KY5rwL7pU+ZW+9dWm8OYULx/iN9SPPiqfhiLl1g9Ivhi5gQ6NrD3e+HAbuLVv
WplIIcCn7XangG28qJHndKETij/yt45gbajd3Ekn1nm+fT2MzFc/2HOAaDuT5V3Y
LA6TK5r/DeyYTnfiwo/g/akRRXu/pzWE4WDCCSDCQe5X+5vpgx3J/WMXM7BGUt5B
ghMqW9RVjzw0lLe3bmWLFqTFVVCm8T/XKVxGwnqZj1WL1MeCnjR6O4WCelmgDo5w
rz3f0JXz1gu7DtmZQ/MHouO1cR0omPQWNGraXXFSco7WCJSAb91ozUnUZGR4LKbd
20Y0JXkVW8ZZdoBOYCDWscrmloqD59vR5VfmWDJiXfWNbSZFXhotlXGW9jhJVp27
LizE0K8CY+9I9eahndFiHi6fGkWgT0hYAx/OWMlftTkEE5Xv1CvMH2yGthFluyeH
nUeHI934Yyc2UUcA8QF0dOpsBiuJxPJLWSFThRKaBjnaXdhuvxhrOVrIHeOaN8GQ
nJh/2O9zIXJht98ud2FmU+bXoZKOo4pHLAF3N/A7lQ1kDgAastNbaSGeW+GvH0HN
bMG+e8XttElhsuqT3EHmFyOsfILodlkAPDMfKob8ic477d9Mbz51QUsox1oz4BYI
U0QxZl7MZoe5z2RhWzKlp51rXZ01St7CtQRZmBevxNs7/5wWV9pjmgfSXh6dDafL
Sh0YJM0+k7AbNxfN/N+HfdxBFh5Q78EitrB3Ul7OHwHyhOZZ8Zb0kaGZCtiGW0z3
Gir7+LUdg2AplmcvArR1xAVj/zJhnEd57bHBbEPcqarf+wSOEkrDml2y4AY3SMfy
o0an2FaDGi8FSTSx2zDDyoLxqeArd5aq23fdrlHMgHbF1F83F7lZcEvFehCXKsif
r2db0NDKdOHIwTtaq/MyPBt39eGdyVfwUxz0xmNWJ4PvPyuTDViZb06tt7C5pl/j
DABeiFJikiXKNdGoNHUB8c8DAPhUzFl66235QZRxs9OQqIj2myVr7ttGdawW/Huz
FeGqyRz6xxtmipzQEBlHBWSbmU2qetTk+9HaFbZZckqR4V0ozxB//Hn/TgMVr6vo
wWrIUHiPE9cg/YvK+LPTp1lmWaC6lvS7q9SOi7rW1m24qLvXrA2GLw6Cc8jBtJtJ
fMfmivMu5rv+dtp0ldyz7s8IJ3fEU73UL+JToASJg0YIrWEXZkuFeiV9sx+KVJ7U
Fzzw27k3J9GczfZAaowy3+SQJ/Wt8NTdYapuwKGyDEnn2/cbCeDJcWemM9hPuK3/
ntFh8bf1tQsUpfMjYWIMVfO7hORgu9edbS4ZXePhYjRmRAEAw2drs8ombBImDj5a
YorcTVeqQsv/veiFH385wG/4G76f1mK6LZXkSJa58Ng0zP+7GkWrQKgPCkOJH5P6
snrnonoofQBv8K5p4aIJVjzvSjuK42ODAURnYrgMnV8dDpT32Nj8g0sKdCHa6XYw
Ko7xPuyR43vA3gR35yWEaQ7AVg+/5Awm6HhaYrvmfVtf3dZ2Rii1tCd0bTt6Vz2t
2J+EGsCWQNDzCwlw33FSUT2PkqGkkSPe2rDarUfI/Ou38/i7pkcKSJSkKVG9LIs2
1Y0OtSJl5x81u/QQeBdYVcjkVWAi8hD0C3Y4FexdG31kgjJ2T4BCDIVRxgc+bkqX
m+90nnaU5tiKjX02PGhCf/6QdbMwTsGNZvSedH2Cu4kg++BIyTQ4aSRsq/vxek8a
tUau8RW5EoYSekqu0ao3cWXUEHr4LugY/8sUKFMmk6TMbN1ceaBrpv0oe4ep6bqm
wJ20yax8N2/oRWUK7imd/yRf+Ph8SNvW+F3jE7iFfcAeCu7hYgIiIQWqLV55sa0f
TQWPpKOoOGgfIuxBhMyhb033xY4WbWubesspWzDaLxTw1A7BScNOX/oyIxhZcGN2
N8H0wEPIiD4M61hbHzzH7AM4/Fd8/q7KSDX+OVAL+1l5eOqoiQsp7oh5TD4GIzXB
yU4Sw/4RljbVDsRhtphbJNOqJIvVfuQvbppAU6PhfTjGBue47J6SVp5SfDYUd8KM
0D2j0pYZsgLaYFvoUOcK8QJ68Kx9jTYlyqQPRgCh9AZlzGtkg4tkg+igRyktXn9c
lUn1f2kfKOxWRiAIH67MJyUgS4g2rQdrl8lJHQ64UnGDROfKhpPB2nuDgfz1Fbeo
Uj1ZPTYzQGydtQaO43ZLYQUVQdfVIN9Us/2FmGCoJA5Unrc0ahspGnnKgSHHV1vz
sXbsgRF7ajG3+Sf4QHJA+4qvSiJEHAQwJ9JCxPmMwWBx9X/7yNLadA7vLpoQtCWt
mFkJquPfL17Q2qkCsHhruA9Fbp8dYiXAhDQ6MaSEa+ufCBPwfb2zi/uYslI2Yjuj
RVlWcxebUzlvqVpgazT3qqqcfkMAZidFRMhdNoixMaqldohMSMEifhhc/6vcM2kL
0EQNyJKXp0DgyvEVTl1TY0KzqRSkbuGCSFf9VBHfKdlhTvHDeASFCXcXLs9s0T9+
eK/wQ8YOuinIv1WD6kpG6R9vw8rA40py8NRzP4rduKDJ0t7nwxSWsNcg0Ms1XmB1
5eQDCnEZoVXEqgRmfKyNCFn+l9u19LAPgx2DZkvHqIhxmIGshT+XhOiLQw3K1X03
XgAMT/UakqKUEa/LqPMujumJiCijGrGFv0i+2C533KV+vTGv2EZ9QNfJsLyIElMk
YlU6UYcaYXmlBuUjANLKtZflspafBioEFLYk6VS5iEeuWyjgwkne3fen6xFunggJ
Yvx4h3OtdDr3xZgN4jqeKToxU1ryB/gvxYzeBRCSyKVdRmj2gkLcxMDDWYvqu1UW
EiEVgiIE9CU2UBiG0gxE31KR2g19sQ6wztP0cN6UibDM/g3JYIofxpqeWsEP5S0l
AGZ9ziMdgY8pKwmbMktvTD28OuROUk5jPPOvTGsTHueAc3d9jvcsfGUvqE84otwS
f9uJHwtqIESkut8UT1bmyTPy1Z100BOWNuUc7dMOXHJZ8dkkKa5AgHHwNL+qoZmB
I9KYl/IRQofoeyWsJIUBLdGMoRkW63LmTJE2dJUu6ZFPL7DOrO6JzPvkdMasLlZ2
0aWvoBie66gDVHcoN+lAT0I6nOO6WMOE8HbPwi5r3xX/XfmWRcz8YEi4q7LFSewa
2NoD6TaBrg4cKBiD6dg8riaK1aBfgloeHO/iyX4zhK0/nO69ILIzWXL6zRvCQNlH
BGOEoMQgt4gmESa4gvrzW65xpAuNtOUrcSpKliaIq66XttPhA2nGoJVDZynFj57m
gc8hMSQmSUl8rWxwhrbApXYqs3eMAt3smDg8SKmEyVc3v659Jr9tHs3W2Sktp3jz
X5l2q327aBCfzaKx7xNwTpFRNlOD8+frnGBl0vpFBHXPNkqN1Yu5E1zWAl51O8UA
iOd2VYzfiRaFlvPNLtRMK2NUAQrmDm0jz3gGy103JPPVM727Fhp/p8N9ZrTccVQw
EHz2RoFWkbqRA1+beS8Pd50XlZ1Xpsuw5ZSwd/z/VXB6llDLBL5dU+oVoxR6wb7R
Su7xe28fWGCHXU9Fl3BVJFKCTjSTwXoMBWTQW7Fp+S2XsQqqpAdbMcuyf0U0H/5V
c0ay4tbWCg9JreO9EZcNAMD8VvXNvs65DhOCdMfPNuXXaEgMpECgD4Ww6mkZiWd5
QZVx2P+RTF7LpfaTX2PuAaHv1xkLj6pUHsO67xV3tUw=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbWAHFpjJHdAHp7mLFOKK2UO45SykDEv+bKy7mfFBKorYVtgWmdlsfbcwYesC3lF
DqMkm2SVgSeQgzc1iblP33O+fCULkYz0xule53VsG3G3gzF8sLyJrB8hdZ52Qt9y
COB/LFUd7iDprf1kNC2BTSPHMucxLg9oXD6ZO75ShZf8TujQzzjZRJDLiy+q09pO
J+lpX1d8FM8cWKTLXKCYmPuFe5YuPlpIScSqh7k0JJ7SC0O1ymjz9/G+HSZVRtxl
yO6yB7omZivJts7R47T4bB8dz07b5IrLcnP/lqtMcbD6y7YYVqbcLjioELI8X2EX
m6sxzYbFt4RAl/jymWv9sGcOwV+BFn5yIcrXXQGXVRT/ifEl9hsQRgA6VmVQ8vcY
j4lP7v0bvnWYVmUNU3KFC+3UdredwGz9Yfx1YFtvLChjj1NiJqosIXMzqsX2M6lw
VG+zz1sc3prqn6vpVWjp5XLZMA7Eg1Kwn2Zt73Ez9A/kQPIuZzfR4aQ2bCUe+tON
jGJOk1vxOgbRwnNzyZvpMh9w/I42byv2p7dnC793YKUI9/y9q0/vXzteQfbTWlnc
hdtMuObH/aCiNSgKkES9GXxjzFi/acGgOvE1N1rnQRM+ERxmn14Jw9IelC6pczHK
Yd8QB8yR9gUkk9+IJpfhS3hRraCZImGpJWh7s2UCwUau3BiOt5SmtzhTgAT9byVa
yQRy1PXOK/zjteNMF6dtB3SxmFoqwo5g2pyo4XLYN+0w1+o5K1/pfFa4vUnc/9FN
/T54aROz8eemhzs5eQ8gAL8AFNSWEUsHGnAJqqvbgg3rE2V3jOaFX++ehdJ3kkaQ
Myayq8zpssKSDuiRHOJUFPSs+fFafygspSIn2LdxhTD6zC6OavEw29dj2h9iNlS5
iSSOtU4QSDIsw1PtUC2vXRbxE+1G9PqzYqWDrJx3IPvkzQGKEPg2fv9JnzKoGczx
Uuct2SnsU2JkjcXteYEqREaE8meUoJbghEVnBf4l6XEqOB3veHHxuOyi4R/WPmbo
ceO4oSPHJufsuYdSe1x2JHm2Ocz+ik+hAvvPEhOcAPTEU1LacyjIgFNzOR/KQs1Z
Wi7aGLbXglzxbzQEUFT02/Da+DSACdYfgBD0TwegWtpCRty/PffJf7+Xe3gyud6C
buoifquDEdyE00x6Zp2fYncSh1+Irw4qJ5wMjWY+NPLrnNUAtfxjGKs5Wz1Z+4GH
ilw0cY1lcrZ4YU3iHw5p2YfogEqESYQCSxLjXq7dYJgV9HBV7sWtuqL54JpZLpYB
2wiR+yQnqEW+OmO4n8LQg6/0RJhxsCdmyUu71jctmWqrqGZ4V3Y0qUXjji+ZuRIM
pU6L40T2Fwe+w3SxwNmJKImPFzbbktwN/e5SFm9tvmDCz2XWgiM8jEPwn33F2o7n
8tC2EZ/boiOUG849NgIv7ZO4l4prFX8KsBFz2Elaybq+MKg/hoE+BtS6rsqq3kqq
PRHiLDO/FpchVRglIWLniEH3FQ7+EkzaGmAoEbxVOC++IqaMq77t05C975geN3kh
fw373xfhqlsN61C5PSsOgXeuUQhKbCFzKOqhi+NG2kFuqLybgM9RhuwI2552/LhP
I9Pk4kcKpc2t9gHKLO1nt6T6m6jXUr3i47UbGpVsYldFTdbMpm0FvIHOL7LhbJXh
C/IqwHft/4kWtMtzd+yXBfPCVDnZ28hxTlVJ419BB5eBitXLSrHU3f9V1V0NyAQL
VRXYHD7K7u9XjLyhoVAt6MlsaePOyo3rumctsj22iw2uc+V5cRPU7Gg+gJ9zvDOf
nw2iGdL3sqfF75yqQKiivpW+kDljpjhrf8BG6BIRPivWNorZfLRIAguKzKEjRf11
NYaIFvAtobRaxbWHpadP0Jw0YBwypGRnfHNgQBsAP7QWYju41QUTUyCEhtBxfwN5
/5N7KxyghdLP/Az2cPz3cutz6d9PETRk8y8em2dCAhWtpYjXFiu6kgcE9EgwdZwY
ZxOFJyLgrdDA+Ucz9YFvZkgaLJ28xbKuGN8dPKo7Izl0BrxLH0LOrob44QEGmGgN
mVNILtwd8xb8OUrdHSbLfGJ93mHsF/BOK+Q1wMQ7vcHRij+R6rDFg0gCTPGG5Zix
PA7Wzh/74ZkyhOi4QYVGXNGcMMcIuNl63UY7xpCxei6js4gsDiV7a2q+g2cMtXMq
+udSx6NvKNbkHhBjn6jS6aCRCFlYysGJklJNu3n/+Lz6Z8eKyCJFeuUZpLVRY6W2
wtBwJnZj6bVPmtu6zNKzu2jzak6dMmg5i3fz0CATFEJMMRE7oDwuK2Qs6LD8NMHp
89hnjOAmhjyxmr6gSmLUSlbHWxYaW+O2VOm4YOANpCTvwt0CNUtoMCJ/PSQpkiGW
1QqviBuwSvey9iYKyrXais5LyUgdAje+drk6oj+stS6VS9kZVxb6mWIBX597o8gW
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+NLJxepHC5U1LCfm7tuLw4u0uwDbnRY2U1OCJ+gQUycjd+FKmn2lQtt0ydvOMhYQ
C5SY09pj7RXr3KFaNIySyrGBLqoUZeUE+G06/mWoVzGBi10ywbbBkFXXX6VPqwfZ
IMhqZuelfFXZyI/aWqOwetypXBgEuDp2836ciHJTxA/b4iyGj1mZeMPPqs4LIz8R
//lPN3Mzf8ffWCmpbjBliNDqsEj+HnVtZs3/P9sEVg44fl+9X6ihFxQJYeb0T1QU
+WXlUTZ0MJyMznwxNQpbL91Xy3p8XLjU8zDMEhHKoyjSe9hLnyuFjGEVzeRuitOJ
JPamqZjA4PyThk3Cby159TUyQpZ5xr2VwmWC1W85GHjhViZ48Ti1lU+lDD0qYzzx
/5iElw6RQUKWNQfXP86iXPeB99uwkVcv4FEikKDNNA86CpMOfan8rHpvZUC+Ca+o
fT4CNNFTyGgGuYX67Ugp98jKMBMbWe7HbMCSoZzJv14Js0yzk/FXQ+tcQX0qMg3g
AE+0/Cz0yW/OO/e1Xv1qSG2nJkWYzFqyjlNyDmjyya8NyRQAN2/7uxNSuvhLeIcJ
hTLj2qAnPP9ETYtwfiCFCXhcC1Pyqo8KzCh2UnMt4VI=
`protect END_PROTECTED

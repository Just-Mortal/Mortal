`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+qQprhlDv7n/zviEJ/oTkDAJTRrr4ZyU1YSQjgSahd0JT5lvQyCxkLhJbhDKcDQ
PKglRQT8hd6miwQ3d0gQhazjtSfUWDDN3nO0fLv4JK/ZSQYbS6Zt92PHh8H/+8jN
5yjuA6Mn2CTCWyBEWgYeePHN/q5Ak1eMi//kiAO3oj6J9aoQCQD3iJF728gOrBK8
0ZqfO0oXfX7WVvl3AEc+c8xM59n5sLlHtgSxbsbk5swxKc0UhuV/fdmCh3Jo8z9G
+19jzb3oEoNnSOGiksuM+PvsfAWNCBxJajenNK9WnlWkX8RQCx8WaqHecW4GSnd9
OYYrBAjLU4kJ0m41QNACJv+jrv9A9IW4TKGF5NfGiYtrhNU4624jJ8xf86N+zMX2
kIIUnxH+73Rspki/xDZFu4wru5DTfJYInHd2SwkdAljITEb3XRTBQIE2OXNbkGhy
JRS38giOdGxPhPNaUmRiaamHPC2Q1C5lRfeWCGVwWRh8WCqyBmCWzK+eT9hdEpoe
0YY8U4wAUVoinZSAQA6zU3iBMte5iVIc1uuk6NfZVdmwmopaSfB5N4/+yDtol+vb
qOWSklJOMlY1ZIXB6rhVxsV82MApkXxngWPjc0Nl/09XJEAgF4T9ddugGikRNKYW
Nv99pokaI2XZq2kF9xH2+S8Fp4+xA7/3xMTJBeY+/Dt5JbCh+ENtAAMQITFlQlz4
whacc1hdMjx2FkiplZV7k6MTklIyjGEQ7kSU3swIXjY/VEwuY3E8g/Cd+AMDTno8
qSYxYL59gm1xwgD0M9F6QmxD61cMkfnrb+5FKT0hUDTW0eBjaqk75B2P3PtAOsrQ
h66wp+Cn3GsWZ8p+QIl2hObqxdqafWbA3mUV9xHqBVlNlcC7vj0bBQDPampdopNE
FmQvSafRrq0Js2KFo1z1LJNg9jCBwwb2Pi7SF7al+bPUCsmtqrX0kAKYxpzZIEhB
zmG4w7z7PMr/ScbMCUSc0ldNQX24NlU89KS42xOuzg1/L44xvxdv6Mg++jJWhX63
oLqpK6EFmEYdLHm+P7tWZYkm/OwQhZh9onpB7nQGtvKmnljf0+i2gZC1W0nl28Gs
duDsC3u/HEgSq7x7mRfsNVNUrKbAbJmsi3fgVKW4AgYo/rJqI21hOddDdU6ZzraK
4D27uIrANsKyXyhkRaE5DAS5bfY7iSai7ASyHVIAimahtTRgPJ8W9dF46JctjuYO
qk4cUfeMABJOwQebKatD1KIaC5rrj/8v3V1vFgKNbXJciXc6P6u+rK7HVT8Xz3El
iEHjmH8OM7hsdTnWKxJVzbjTNcS8WL9QDyUUfpnu8eLbYi2TqFQfyncsR4tS4f5R
/e6/ClI2rM/2424xneNmqLqafhuDVv1iOaD00SpHKcamvjFGxybQWSbqNnAfE941
+1AbNfpx3D2sOQH9moxOBLIjj4gbUn3pntHLBoDrYkZMR+ssrJCYdC2Ipv57/Idn
PleuVBHCZdLSTv4jn+19Gb5WpcUpe+nXH7+OWU3mK8Niw7AdU0eMCgGPbY3xRck/
o2vfqIq0zLzlFabB5E0l1cVF+IsLo/h0togVqgXKTjGAlDU+29s2VSIx/lIwHwVY
liZjQqF1IX+d9GRv7uaAk9tgr/BCr9Tjs5JzPEvBnwc8qU8q72p/DoyDgzI+ZS7B
+KzS1GaraaGPHV7Z+/1KnwM+4+sfhasccswxPiJSeGMAarcy/Rgvxopk9m9BwCcJ
xFAPdmQcXEMBrTP2EzaIJ3yV+dZGqmMzLbbQjwphdDd3hS2tU4tlAl9PUETpcPDg
40BbBfX5MDs0JmxVybUxpdNuFgkWV3hdCUL2Ec5Tk0AsyCnOreJOdetrKJQOuzVb
fuflGnRtTvY3Q6bu538a7OQE4KCUlaQoe6q5OWrzGBuK17YNVqxH7N5X+BzwibI5
7F8ZIpsHzptzBbtHyraI4a6mxlEfi0fn1p9USPwIsIkAMmf1dkF1SV6C670Mc+CW
1rzw90Z5E6ALDVGAomL9eM5tdTM99x1gk1poDc2nZAbMoavM8mNmP48pYqdkdXfJ
+8XAA1ifLfhWoW09q7OURFdWgXzMWuTvPBYkTnpGko4so2m2KQFIEqWoIXkkthGR
JrUQuGDEYL0Nck2MzueLppLqzDvKtlzJdFtNpGMBkC6LJNE7sK4oMuPXFXNhxnOf
u+e69YBISw1ggZJSZfZTP5jDgX8XLmghI2mWVkRq5uy4uyLY6/N7JFUVCMwCCXiU
syciQLrMx+IERNN9LMd9oKXVjc9VFunpTpIx2hqylgaQBYaQZeWTes+JFXHqxPnS
2ziMJMnmcbETVpoK2yrMQGjMPnJ6vmhRDnRQko4bHUIpa50HrD0wnjYjs6YU9rfQ
vUtbCp3aYxpx9Sl1Nkj2lgJbbr21n6itWpg4e+cDSQHikfkFYQcgbluQKbOZrMTT
KV7NHrqedJFt6k0CHAgolhDYxzjJFPegwwYt5OqhfetwQSw2QDZE2yQ1Ts4xeYpf
9HAFd34Jrh6RKTgJySBEOD5U4RbQHhs+x9tR8iaSccY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgqucpKcpNl699VwlTDfg1qyeNQ8qk4oTnwkxF1FSJ6Az05ocd9upElgtSc1bRgn
DEnxkiN+R4eVOB03Zi8OKsRXbuqJl7RTaQQQIjv59Sqf4jlKcTo9LS0fXecIKGd6
fuW9buz0ZzMnRymgtGUJYxCtrFnFwaVJCnslYDlPKZd3A7u23TCbs3bVbZFI59oY
YWYn+Tw7ixYqwuFiMih9qBSiD6e+69h4jbg0IkRd5EExAV/Ecvm0gx98YZaGpcCX
7NaV/OPnYbBMKAQsmDfSGcozWa1qZPNxdh8BKThGARuwX/28117Kbeu4y0H2x6Cw
JMHND6ilpc6tuK6A3NLZ6SvusXpgNkt6TYNJbCqQdD5e6rwEQ7A7qCF5284TLUvN
nFd0yks7qB1jNVVuQplRXgFROCXhOuAS4kdJofW34BqosTdEqGrtBIDdAqQkS4Qh
LB6OFH8MeyxXp8V94qzcdBzIS2tem5UR0akhT+OhfiwY0ofPu1T2+RQ65cLlgXoQ
4/4izNtQ2z2MnLymB1oh/TeljkRnwrtanvjuQYp/4a3/MIyrYS7G2iq0MN+slz6W
lzOI6sZIVpM2KlkdfYeZLri7/Ol4s8Ywz8KHDGfq1C35pn1R0ZAzTNK7LQhgfx03
yAZRaamO44txD+dOGEsCGb0uwFEXgnSVY3C44hmHJ7AfDFLoj6PsHOMIaase+f0N
PXNfVSSHdUhYSETzqhKA+PvzVhsyuOa2BUvw3vFE2iat5MZTjqwCWTChjNvBULKX
3BNQKJRJ5NGiKkHhDqf2ADIaAE+erJqW2pkf9nSjZ5G8ev0oVh0x5XqyUrIH/iLC
XKpBy1C7NLuquolM9nOpiRRkn5aQHJRT7cROXWqpMoSmtlfC5KWZ0bnDucphfLnB
++8psbdirBnziS/4GJpiQZQgx/o8SRqP3SAvGK7DOvd6DQfAmaJlrFEas3HVeylY
MUt8ouW7qkux5VGG2u0uubdswIwK7ZXQyEmY+5E3LbDtdjXFDOEQWacBRHTHJqEj
12EnaQRgabNrBlP0eBltPgbZcHJtI4Rdbatm38bYiTyiH7G6+Mxr6dxzsaPp1bFD
auOTMJ+TBCtMj0DVK7yvrhQw95YzImW5BQH3Emx+kGwO9twFZT9VcLUr9WHSRUW8
`protect END_PROTECTED

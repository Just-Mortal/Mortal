`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9lBrmpyqpsNKSh8F/nlKffC/HBLEM4XMO/qs8U6WIMTOof+QHTiZtjzoZFBhWSEu
JRzyRzYkdqE5rcyU++2vngOW/dZbYpTBbp+GM0TgIQ4k03eV/NUAffOWQh5DgHDo
5boXX8cebJudGGUwajqgBhaz65ix3gD6htVUZbtrOCe1xQMiBwzSjhLM2lRPmAnS
A4LXRInCMnR3AA3Z9Oz2iNl44jck9ebNenlWWiDanVmdRFM16N3nUUVrz7QX4FXg
tQXOJdNshLX5u331rD9dg3A4Qigxi5ZLqgHD3z1fOSSrnGd3CCY3P6oTqo/BgTmF
0csAfUP/zi1Uz5Gxk6UYa+GTUCQ/KIVOol2rIejt81Gh1ULwI71y1bLI3xj2sWJ5
13Rhmw6hxs4lwdxWf2OI9Ueudu/yuGP7t5xxDdr0XNSPNzvUn2q8Ytyc6XR+laJg
TbUZ2dJADABuhwbnW+YiifHsiLlhmquWkCJHP+GVKG5nEOwPo7A+gVVBQrwlUbK/
0Hq9ZuQlqNDU77SJVKFpxi/DG1Pu0aJtKGzwYYmAsTX7h1klxo4vvVkY2iO6SEBD
KEr3mIik+xpJPWk1tP2r9A==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9Btjuq/NnzqHgKlqWzu6+bL4j/LMIzp2n97JmhjB2tMiX/qmZ6UIo+C7YryzYoG
XpHVj8LuDqN4QbgcjK3Jy6ZuFgBEo5BAUyq1K/n/edpsnBl+D89OuBOf0YZPlNv9
/b0woNWrWevl29PU+WEMxp58hZTpdxzcjdY1jzVRB/misVuIhU11LNkluHi1UFUa
1KjOl3uAsHcXmukrkBFcGmMZ7DfgEx3QVO8AMH8MX+EqCb2gReBidahLOct5NW6+
NJPXD7/s+tb7+KwHGuBDMcLwMEhJWT6RRSiPNfUyHBX/oribKiB9C6l3Q0EaaLmR
Dzoq43Le6QSwPkmaNSK4VbD0Bby06byykBGRRVILirmCnQ/F6/aQBhDExSlS5mxT
/JJqf7tzqbxNTg7Ue5lX5zvI13aiSz0XRG6stNZErGR5YAOLjvCWyfnGjfd5oonM
YH3ZAMhAEv/X2imV2RPBUO9pD6YFLhHkjl/KXYjRVjQjAoVcAIgksOSHCKf/6lWo
X7EXc6TeK7wiHMLJ0xZXWtJ8fkFtk3FZ6+cE93tw3mTnBevIRUmwjJVA+D4/eZfg
8JnMfxc/xVl2s7MpIAahWZ0nTURJi8nGzZknQCKwqrHY2d0N+hknaxRg7HCMM43B
+8DA6WvIsIHd9nCrKOYnwYzT5P6VFUVQvQh89hpTewELaznD+0CLXrHb46jkpGNk
2+/jLWXi80JiIdp0U6X5QOAe8gFirytTvH/NRnpwIyBal+HHyYeLQKYAZDLIAuFR
IeScwMxEtXL5HaijZYWa3JZg/vJwoXPvdp1xdS0oFOuV+mv9GRGnMqTqgcT8hRWp
d1cgqlHwi1UEIhIErRJb109S947OokPXP0n1Z91L2dwJx3EcxSv1Q/vPBTLMJPqY
XG/GEDXvMHU8cJy3DUofG1/bU/YKIOSnDaupJhfUUqtlxnYrvDomDtR9D85OHRlf
CfOhY5dpHX4m8TjZut8NnHicc4fjm2pi+7lnQQmTrpxaOjPA6ICXVk5D+NkJo9MD
/NBFSHtTBDMyWFPqOHM2jHuUAAVEW8CSedh+Zw7HVZHzbShjx26f+OkF1kGAlw9l
RN7e3Bt7VX4VYZQhAdImMg4jLeMvm9rBWQD0cQdkWN6MmOaEkuAEUYi31RObDlB9
50rA1OKPfFYqGTef60p86j0L7S9SStRE/wHB9t3QqjlBKZfa8gLlkB+5H1ZDGnw0
3KtGPE14EQrSKjZdVerJjYkEGmms3mFPd9bulmle9D25+kb6qtomisi/KB9LU4fJ
ZOqqgaU2NTPXkA2tNgrWZLYhO8Ym8lN9elt1jnjKFUTwhyz1Zi5ORT7IWR1IZ8XE
IK6tZjninGktED12jZNCdWswH93rE3RXAZI0RmocwFQUPsKZMyviFanRctnhtTE4
+WtVNi0oLOervEHA1/5q4OEFBOEPGG1OOWCPWV9nO+8eEkgKTtlDjrH3wYDCsAOR
Gt719+JJ/anHGuQ/vCP5YHwM87V0DrjB9dRyIQMvVAHpthoLo7O6HVZyk1lRmg5i
H1EYKcLHAmxA/XOSDM/leqPgKzL5TRnvgH+JrN27v5FoZU1ntYUGHLwI78pl9IaM
MhJEizJ+I7MXhEqVnTPuQr1iPV8AkaKnFu/1hr6rPdufQC8SYMkoaz5iHmsrkJIF
tFso3t/FZk/OwMix0Ge/USb1d3RraEOisVuXhtHBG3VDWSwHQ6rUyk5Iv7Z3GIxx
M5OQOxxd0kQryKfkmvsrlhHVhzB0H2Mi/zmHFeDsi9ns4cPDie2U/q/KphpUhCu+
WiPgQKgfp86sy+fR+aBDEeuM1unch2tAsJJhtpIDfvXVx5yyobpvBSvIVDYNLh67
Y5ftqtmFtbrY6YbccYhBhrtVeSRTFxSY/mRGHNQZ/j3ndJa0cgFRUtd9+RMVgHvB
OZxPCxJPfOr5HsN9twyp0lUZVz/tfFZ8s2QGUX6fMyVWmDnuQ+98amvWBirRakX4
heZ49fR0WE19e653dm4xmWP7371AYuItp5JxXXAGvtYm9WKOt0/4oZheq2w7ElzH
8X/LnlLfTwsbil2UkxBvTjBysJVFS+p/QRxHllzPBsRFYNbR5tBesfvHyomL7zQR
O5sRm5ZzCjJtB6+QhwomZu5W2L6VHRClWs2PZFPI+uknYLZnsm1DjTM9dAqGq+qH
/PDof4sLKUAnQkX0WiszyMkwAQ9lSK2gGKvmAA/5wd2frvYwrohyqbJR74uDEXek
mvlOdRQDkC2V4Cj0UMp5Exdv09Lrz0rt+b8++EwPK1Z8UEkEMxubZU7ifc2xOtg2
lUSvJLlIHGfPOGweCKQDwzt4yM9oSWjeNya515oANGwwHm/6igS+ad4sbdMN2wK3
tw1vWSZN36aIyZRTwGboM/C17wGbUj3Iaavv0akZA6un5OYvLvyU+hs55chY4cUD
wQJ8CXAaD8+BIWv1xtA+4Ia0TjgdM6BMvhOAQtg1NhMcBwH01CDOtfARWSg6jboU
puICi0v1FTOTNTlXg2uhCVPK/KXReCd8nX2yKQNq1iAmi78oqIFXfgYmia0Jlds2
tkAQF6dTC2BToZzMKeU6qgBd6OEVD7AaFt/glf1ujkgTFlEWiKbmbRWW4aO1sG7Z
Y57RinxuaTtJ9WhG+wDRFa5ocfu6HO9RM/C+jwof3PV+UTyUjiYS2UbPCOEDHJqE
02uYxkxHDTj2AplyfvKQGIRsBKRnEZeGoVMrvUoob9bRZ7mSES7B0yWMMChB7/Qt
UyHCcTdp1bkMK5QB/+cz/BIqaXtehWyGJz8fhoEFvvZJVgOgwgnILYKZYYGqYV/E
jW/uQAz2DyBhajA2lFnKmpaKjwWsKASv7SE56Xt+7wT/PbP2ixTL1f78LPFZPcUU
r+bmspiEQ5RpCBR5mq5+WezzA47/11tb8kHKIA16WJgn9DOYUM7pjJM33uIy9O5g
d/DhlF0BAeeNi2VyMzTSc828YgjCEzMwQImnkdBcK4K/WMqrrcpPmXIKyaVwoPr3
KFzgBbFihh3G0+O1L5bjDIH4QoepDjiHxGhp7FjZsSVvwB8zx/qI2j4eLprVyhKh
62uqHdFzG+8qBKpbtlbSHQMdjfXnXu+/LoxIQxYp/zMwfWgAr91N2Ci0Oh0rfMhm
4CyL02MYnUmvScjBhAfBrPmmPrlmuFI7mHPlxl3CL+Nsc8KrAuYXk7ITrjWaAzjk
O68lIST2Rz3MumTWs9zW2mPzDOlT/ESeNlowrQKro0w0EFVkfL8Op4A9KGJUUvYa
NpWmfskPFqM2J/oc5QtqRXvO5Uy/VySg8cxpTe9m+a7w6VfzgT07en/RjTmhL/Mw
KWwOv/JJg6ar03/Ag8FpHQ==
`protect END_PROTECTED

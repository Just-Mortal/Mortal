`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fAz7+qC+mkE6wvnvJKRWH5no+kgAyccZPQmu4h+tBh8nmRw39NmeKNkrgiBvx2LA
c1V99oCEn05AwH0MLhGfmwQBl54AnSYGOU7lEYKAP395ccxyIGdv33jVPzlj68Fi
sGdqiWJ3CLQB0xPi4f5zEJeoZRkXWCRadxcNNzjF/ZJIi0NPyweb+Mjx0hNLbVds
rBlYFq6B+jUhULK8oK+tIhSEqhxd5/XMjVqB35tkc6qwJPyXGzgYrXI28/zhbxGp
NNd2ryjcSEUiIct+XQJ77VsNv85nivrSxX/uqr2ZNtG2Ypq+iBIPB4lZguyf7gDc
HR/wDH6kD/4CGTmxvAopJT3tGfzoOuCDK+x+mg4g0NerSAvhn/ji0JXvGOQ05ns4
+550/wGiiP0FmoifU5PLekuFUL+0E94oIqblJVMcSj1SuGyhZZqvyCGbrRsQGIA/
2VE1QIJ16COLV8uKfJRp7zBhvtQmlD6wOe1UdGD/3EwL5TOtM6NRDDLHjmRanGVD
XUUrzenzMvtJ/PeN0XfcO4a2U6jErWrK/O6Dlvu/7vrUIQ7ICsv01ST4SQYTdGmq
QCyGSR2maIbaFJgnuIkr90DNpF7CfrxucNY7g+AsaZZHPwpYk08Eci72/WBjFDx1
MnHdy9xvH4Rcgg4OzFRy6q2vF0HmQFXkJbLI2gcybZmRIBCLFSB1/tEW1rugP0wn
7b6u/ivEawCJBwvCwD2Cc9RMDLhQXp1bR/zypJlsG1FvcV83MSNRWJh6zz+qLien
Qs2jwdkYk//2DAhzW0/Em6K5r7+DSlMYqtdf+pa/UcF3+oRc9ov0Ywrt1C6mAaEe
H0t3TPcOEk3QsQuCeeqnvQGTZa1ojbfRIoLQvHp8j8ZoNCSf/HwoO0Emt0LHth99
lWSwPyxsRAzvXtpMLqeMDQ1OWdJKEYp5+i0zg9TpAkv+hA+0sp6+Isw00sl1sEDP
DGNcao7hSVANOpEbbHQb1xiPq3b/wg9gT6LaXJhW9M1mhQby3J6GmBN95tMN5sq6
0rgTk1+a2uniBcNz4kB7/y+TjxK2VFdQFZR3VqpxtBXV+YPPAmuHAYjnCn1hIb5/
akWeAueEFXxSeQQHQRArFu/9N+fzWznRUNx/iz2Pwes308Q1hRygMA+ZdHvhiAci
LrswHK5sLk/xXNCvd2SYEVkBD1nbaDBfgiR3mlI2iUC1tj3j+o7joGk/hpSd7IU5
/dCp8Ik1xiUNLKLmdLTtBG33bXmV23OveXSe6fbc7gw2pCCfrUzg50dH33+r/UgX
6RKQbIOZa+b30rPySJsv6p09bXbtQ2mKGZWqQeoA6uvRVrL7SnwFnOPTNN9/s3kY
sRnHvsr9jFyQHg1KMsIpzvlaYiLiUo6sj+b37iwViAhITvreklFpkBIppzXqFwoT
+8/ca4Ps7c9F35I0a+QP2zaIF8fSNk2UYymW29ymXsVx/8LYbWYLKqEw1hhrAMoF
A+oyMp1Capb5WZUyszhvnYqexKAaqobYE+jUOVesjgJ0HZTAldTAa+Ekdq0Psx43
akNj7FrY072ctQ4tAargCm+f/63a2k1Ug0wf/n3AWYyYOAwilOz49infyGxd4GFU
H8yJW/qIWMNZ5DhUrBzLK+vzt5av5ZOJMQelGUADCxmp0ljrpVLJn+HZMM7u1ecp
ZuI2K6TcQxikDEc1KRmCJromw84pq+JdYo7QffutbnwtLKWQgz2MDeXi4Hs0yF15
jBq+UzsGUvFKXbwO2sbPwK7JZP8t0TVAzounRLpD4LFe7JYv9WLApgAzoMUJwor8
gyJ2iBiOTdipEJu15D5Qr+JgJHCoUZ+1zktwlcjb+MFqsumaNNb3f04vB8rGcMB4
Mn4Di/CW0lb7BxTi/GGkofWRBI5HA/fGWR7Gi5b8CuIAekkL8uW3crfzu3gyoSfw
Ls5qIRGNZtXZUGuXi6hJ26uwgI9tOEWTZ6Wdvb49SBIM55AgkraKnY4wlc2IBPAQ
YqAIhTQ0vLJxTCUZ8Q0hAeKsrLM2RozKHnhW+AcZDlx/yHmYpJ2OCubixSBBtFLT
gE865xADPrH7bVHrSs7WiATbVYAI0hLAJR2klUZQbCFl/yXsNbl9lejelqEBASPV
l7QXsRttpK4oN32UhZxxS0ZSTUQJ0j+zKTjcAq8Y6ryzLsA4jB0f3FnzdxsxntlB
cc/EvieWzWl7ciln/1su/wZlgq82RgCXx3MxonHKK7anW44R6GGIRNE0iwm9xRkx
o38+aZFoiXLgQin2DWgCkMN2Y4is2AR6WdT/LPy2iwax9jLwXFenwtZ0c10q6Ilb
fCtJ/1WDp/Kd3uiiPsxv+dCPLFs+b1/NAudXzAfelGd2bYs0tvGg0yAeSQD4Zvxk
fWTST8xj/gLHWVloslQUmRNZUKOmwgJHXHjUgxtWCwEWGyipidvJ91JiIdCnLg9/
8jIfHllNrA9AZYzsHIluHUxTFxWfdz0532n++emX+LUU3o3zzC+GBtipezhXWhL7
lnQyLl0A3pSQNoIUYcAtW0g31jiUL4ZjYdR84MJmeRQ=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJ+K5X/RPNCrce8VYLhy6/PdJLkzmulEchqPOoFAcBNd/n4wS1kdOGsBVPkEDwkm
4SLQk+CXl0sqhZtU9m8J9XW4hri7iysw7xaZXYT/p69ShCWqpgE2wCmi6Css3CO0
AYUxi5j9ifj6LlgHyIaqvDjZvhzj7NJX8IdO1HJO7307T+8abE2kQmJHJ01KVn5U
izra6za/ae1RJOeIp+w4O5lMddrMVhjyfEna+W3YFFK42RNDIxRL3oMWJCKVHmHI
aY1eCj0fa89tLDKMAZf4/D+826o8iQxJe4nrAyCzRlycQORNWYrvk80FxX+2BbUR
KksbvysLMOZ2sE9nw+Is6OAl14j1UCoseQvymonmHN/cdt9iyym8GnQrPoQ9Cn2b
4U30RFwv/pa/zpH1Y6C0YARwYZ5n/bkfK26lmUbfYos+mTblvGJ9GOhYZ4WEkNAZ
mfWH9y8XyiA4d+Nq5dk/hu8QMd8xWwEKZNpAMuYSH2zWym1kpv9gwGgYwbRN4WA4
k/B+3EnoNAz6LKRbsZ9iJ1iFUGEqj7YdnnQcyG+15mGGcg2lBhEuMgn1UF4+FiPp
RKZR8MHG2jHhAnb1S4lZ83deTVn8OcWqc8Y3h/UWtKQ3u6yCticgGCz9ltvi4xWB
pdCt4HAHDhTtBQztqh+cHYQsipp7ZaKjIO9zLMkxjJLDRFQEfnVwvIJTnxYeEx9o
`protect END_PROTECTED

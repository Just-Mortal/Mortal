`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HE0xGE2QoP3DRgk2jfJif6jJIsq6o6u10gQ9IboNSz4OjQObFZCwsZZIMiUpeAX+
nYoRkLs5jefENvdCA1Gis+IDQ8ocbFwS4fzv29Acv4o7izc9t+qldevI3Q0oQxOu
xiMxQD0A54DDoX4lSrPCW6/b3AO2OC8NAR08sgGyBA7S0dJdufsgvUXXF17+4uuq
C7zwy22InxITc58NEvM5os3K4yniHpZh2Ei0CB9FdaI8fJGu/mp1ypTdcSfkpj2a
Rpz8zj2xeRuXsXjgV89DTaf77kymijJjnSn/V7/9HveShFSX2VlOFF7gzY9PjCY5
zY1ZyyuajjvEz2ssapbzDwW74LgVjFJZH6UUaUJ2PsOFappD1XbbYIsysCVeeoqD
Qn/8Xk9Xhh4dqT1oQaDJFAol1W9ByyADhJGygPz0EKJqewb7smLI5sPYxse2+LLV
Q9fZXqlysvRntcGm1ymcFPdJ62ZLPi71knhqbj5p+q/k3PCT/WaEFAHhdUqM546Z
ey3Y7E9OkkR0X+HlV32E5cyoRspMu1G+V2NM32oopezxY0C9F8MmM5HstLKQsqKc
3G/fCaKWE4Ip5FiBxgcplQ/QXEnrR92o1Zlae/FXW27qwrrbPZw09Vv/pBS9l8yx
IKp8OYN7qR/B6kdI0ucexhHLREqnAAwHHwIxaWhUAtI6e0QxcQk5gKzyWyvipETs
fO0XxFAanXWKEGfTNwj1fgFJfYm99+RvPUJlwV7jqOdB222NdpOc4AXLbVbNKW5q
tTmRjb3cqaQeLE8XMdoqeFPTwObBpYAO9cKvnzTYe4rrAjDKtANx9IRPLMdYs0M0
zMGeHKdD3GVYRp8p9ncMXPSDB/5kfOKSrgJkSlYkH5vxRb8vbLCn6bFxnupIhHEB
Qj8P/nLRT3uBhyTl+ARNYUE+G2xBYaL6Lk7wvG3oOPitJRAfW2MMIonDvY2mQLtA
kGkAXdb+8hVxR0IUuD1X9+pREDSQNJJlXBgVUTZDg1GEy4dGkd8I3wE78LYL9vGa
wOGH8azsy6YXtFbcnAItOuqdrlgsfNd/sg6JmWnfRofjWxOsditpwiFlOqolhllX
HzXY6d+V5tbPEfBLkOgbiE2MfInuKv/7qe18QP2rvcuryh8IP/6DLNay7TEhYtHI
xIRLoZAIwG1807kF1XH+tSM0Zf+wxWfkAQOyujC0HLv1TRKv5F/F8aMFb4bBk/XR
j1PU4bNZDzVKYaG6o6GM1ptBPsxa00y/KMA1zRmtyy7RpjP0Kngd3w8Gq+UJGl8r
3w026pSSk7+vz5Dzaf+TAMH2WJ+IDebjbtMcu/DgLWmx1z4U+BAyvKD/uh3M3XAb
7LSl17DsLoWuBeYd+u8Af3NTpgRpGbC44a7dAD/B0s4BtowvvIQDO+uyR7SOjMoW
GFvo4x/TH6DJM5Iz3PEvkxB7+ZlyClGUcDxkD8HwFv2rzM4in7k3qzVV19+H3eGr
mCUDberFqsRBaHXLMUCP6y6sCnFa/hJ8NAmkZlvV8VwIhYOGpCM1Uqr0sIU3AQ1s
dCmzph2LPg+0tQmYnlY/C1aopqGkJWOJTUMtywObB8v7gA448j9YbNPQ6UNks3g4
Y8eZHgM+UH/a8u0EXoCqEX/ft4dRu4B7XicLVbbxEHdoNY2EY/wKxHfH5Q2c1ygv
R+e3ej8IahPYbkQrqBuqF2mrMuBO5B/z35vy1E59hj4yVDOo+yK5FRPcZR0D9Pob
NV4wbg92cDW+T2CKILxVeSq1VCHqGimmi/D4cOBHi2Y+WCGNvY/uXjAWtPWah17Z
0zipssLixp5oUtznHIWLikXcKvRqXGJSEly5Om8o+8iGcmhwQs9S0nmS3l9GtwI7
0oAIAyVSJDMyaJP3Ph11uVu9XDouANy3h7FNMdsVEkVZfCjpW1lz9Lo+3GDJ/9RJ
WocUYD5FkU7oM1p3nkiOfz3L2z6jhpTkknqStGqUFjp776X4137VQadXEU01Vkg5
eHwZkpc/SHnHfO1cRVSgIQ==
`protect END_PROTECTED

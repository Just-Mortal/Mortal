`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E6vqYj2sbBaZS8YKzroWVYhA5vXcW03VXyBcK6zks/1j04z120wGlhMgRVw7gRTL
VpP35rj4TslLn+o4M2HbwfLFAZlFHBzro3iLdykrl7RRa7TorQOwJlRNPQAkitKA
TgeCJWVSaMxmCeVlGBe+9s8zOGJl9sWSlt8WJHjhzTEqWI9T37HpcKJ0VXWyEiO7
dvrws9QIWJhTZo4rFg7tJ8alLB5rkbm5LW7AE2n7nZ2m2EA6qT4d3Vsy2ENJWijv
k2C59v2NaNtLSOTjRKnKS0tPqn6tZwi3zc/azWBs2kuzwvR8gDP6PQxFphC43daE
8TzlrkXRaska26zfhhdb2I0xBvQuBvG4F+QD1N16tWXShEFQFQZhjHhqdlrkHTK+
/HYY7mtEwuMDCmjUVHI2UJnGQOr8Uh/PfJBhAy48yZGsWbKmEStYvhwOOn78CVdR
yONaDrL/fW9eVR5vGaIhLXINgMVxN1gyY+caDLcv3oGWqnj+YL+9Mu+vs25L1low
gt07bcWt+ykdEBoIrnteosAK1peQUomn2r4hsfJ/A3KC9WwhSVVT8q4L/YrJ6Fbk
yjJ5NjSwk9guQTa5tfAnaDAV0y0eUupZb/UBXOxhiUmtbcLy1EbYC6mAt229/Ngv
XcVVJlEAvywc8FEKB/OO+Q5xRvULKNIzp4vo00OOwqvUWaobpDKXKsNcw/dSFe6Q
8YosR5CaPSc9u7GEua5dcPAPw9LuMDw93sYx//flPMDGnUx3lqyb74XRMRXhZxdF
i8m9gHXMR9OYzMfBT7dXYg54Bck+jVBmE0ptZXByCFltomclf40WHmDTu88QzDBV
2YD3ZPvh+wH81skdKwCjC5omIUv2s58Uy4acm29q+FIbAuqibjqWWhlSL2e3Q5Nu
CzfgIUNKWsdoE9jbAi6UBxG5k5iOo9Fl2/dHxLH33KKvUXuScmhbfrBnY9BnDlnF
TY9x2TlyEoe4CTT7KlB9Oy819ADkgJRCW6LFewtSLt45eXPc+mEPo+H4WLHJWAd9
5ww0YHXXQ4QYLZuzr4hNOwrRsumFOBvutQaPsu+2z6iyh3lesqqJPVrvwiptbRWX
aFJt68x3YdlKsC56SrFEBhwQEqvPfr5CGWmsWsjLz8vifyrhVvuD1XArb23P83yI
3+CBbX11LypOcu9/jsMGKsQ8QPc7bgoOauSmF0Qys+sUDDDFKJNjaVmlrH4JJmGA
eHUq0XHmzFxNkIPNiQvInWo3/TH0yA6lgfBeLEtnls+zEYkoW1fwQ0FzSxAIvG8y
mz7dn93izAmRipOgWYjd5Q7nfFb8ffkLRuAhvVH4337BLEOrnUT9VogDTa3k9HUl
farE3RQAwb7S8eUdEdj1tlt0JadYwkjjFhGv7D+oeInu0GfAli6uuXKRHrXacitt
0qpyD3c3MMW1omZebwvU++s5X1EOLzjZJxg+jDIS9CfUtQVCy1jzN6asRBsn3Xrq
8LVffrnZ5JT/nagRaTFarAv4Po82YLCZ6Shikmrcv5eEoJr4VhkevmcVvQORBpP6
KxwwMegfQc57W9csy12ZkDBOUf7iXvpWqHfYMc2jz/NqVdFQA4bG0vJchKRycWME
pfoIy5cl6+s2WdqhI6vSXwyWTPGLnvIiXN7291H1ax5pTf7r2M5wQ346sZ0mitKc
wLLBlcdw0ojI+e7hxDX2ksXEUudTDZcJO6ANwgDk+ehGbtcdx7c7w7rLZr9JZhbF
d56OS9TOXgVrvCLEI6T2rIscLFgpggob/tDMbMMzGtJQnyKaeMZVdpOFrVpseqUS
CK3rXfYXckY1L9iW2C9qgYFm1PNzjvoSqj1twnQTfdGtJWMa8qBug20/6DTviC8O
pb/QH4w/k6T+dxsjr0+eMMGkj39Zb7bxfkxws77mY4hRWP9HYNtbYTOvtDR9o7Wv
0KQIM5Uhino0VnzBmAH4TECX8xlVHGVjRdAQn/cKVywymuUt8XA7JRuczSZaLT4e
6WMTHZ97Y3YpbxMeJJlcXC7ZvIm9ChkhVtvbcxGOfnWpFpssFFwdoL0ChunXMLPa
0+OaMF6MyBYC4jJhD7VfwTz732XGMv3/bkVufbXp08MGYB33OvWX3pyIdOv8lu1G
OuHQfXXnUfoYWdY/4bakz+rGVZb54+7WpJWQvA6mZCCxG8XSZEUS3DyHGpyb8Ajb
+XAsiwvhkx+LSYs87qpmQ5ZgWhn33HTRdJ2lwhVAaaIAsz5MAZHSgeSv3DKmHvny
PCBQu0AkRH5H58KJkl2pEeOXWvLCsVee512N4htjQGmwhcqQeKXW2YTGppL+ueEq
172HYY2SqH90CcDUFSSfDrIZxOw3fiI5ufl4dTnqQtNoD6dbmh/TevZDHPT51QrR
jZxHpcRoad4f9IVeXUkin4jrwuU1Um5COzkPUmitB7zXGMyZu1eanl9eTTyuaASb
/iFqf3TSu8sfDwvwB19ivR4CVbijnBUyvOdH5G7Ur291sb+cnLE7qpk9fIqYCPz8
Ot6zLEjA7Srl5Kze7/W5HBWR4YgJsM22QhTZY/qonslg/noExMH12n8SOHfpsFnB
1AN3IlGpElYoeQ4Jq5SxRYxKjiZ/FxFTwoWi+2a8/V9J5MPfhFkGBLqZpGEXN7WM
IFbltqSN+4EtqO6ozsS5kQuzrIIxyWNK2z0Q8cYAiJDfObkLkzc4uObBckN6R4An
U8vYBWCQq9zEsdPtOQoHVhfgFftDXjb6k0QCPI4VOVBeXS2pkOFga5bZVyINcbF3
nkMJCOsUrK+MwCCEJkdoafvV0yzbH3HsFJPD7A5SKM8pHS6BDrknmv/LjB5X4KDe
RLOwV1Q/RAIjh8PplPV6qdiTWwAnpBj8gplmezibimovYVDG987hSgbRxCuwxrY7
lcA3ZVJPlpnbv75wwRtO+ld6W4aUDGO0ldbElcXHF5Map/sQXZ5Sxcl/sGc479Lo
zJtI3NcSKaNEa4Q9NuTuv5FKM3urUb2K4k4qo6dPzUyRsQKLoOfGQjEuJzBTDE6w
5bRqqTzCNQyGjV08wHIYIPXUI3z10MWLSlGwmcQ0haprAh6Z1F6cT0y+OohOv/9Z
dUHa7QU2s4osH4YMjtpU5vajz1sy5IAJfJbXmh5awjq8HZO9ZjICoC6WlXytSBQj
zt1HzXvjaRARPue2ct5TC2gtkOe1mZsXHqkUzNGWMJapVVYXwrYrYPysG0iyTZEV
eEOfAfbAbjjpQANDf4WvsZTjDZ5Bpi9b3I5M60fKBEKjEPlk5ML0VhwJVpsPwWkO
74b9QLXe1DCn58n3oR8+UmF/IDeQqJU8Oo+cP0PI7csXStd4BfhmbojDJ/yhHH0+
pbr0BiyHjth4nPkkmJ6ZMqWPQd7f+Wn1l2IENgy3gEOlAxUVG/Q82RliOQMSeP+5
dCv7TZfGhLyxVWpYAhIYAnVxyRDRa2PEax1paXgdLRgHPuTvvqsnJQyI7F/Qw/3W
ershecftbuQrk1i80KmbHe6HGFzPt97FLhmr8rHlSnVYc+fqURB9WsNIomKc6XfD
5CrdNiJn7bHD0kjlU6U6AR6gqRmPahsHDqoDTfZmgnhxliFyMwqKGKB6zwim6CqQ
2A4D4kkxn/t5Wo/SAUfjkegoMhXCkW8aQN4hCTZP7iuiUgeBiHR78xjxljGr/OfR
j7jiDp0aGpyNWkzTOGkatUf7ZA8wEW6Ve4L2z2Xx+PJbhvsSsjZ2CQVEBSZPqoxZ
NDlPh9OldzRsMoEIzDO2J84y3YnxkCR49SxDL2MWdp+ZZKIat0/0z4e8n+dDTU/f
Kf4Kt2J6Dlk81TnL4ElHGkLH3vex5KvsMsJfSGYXbMqJ/la6it433is8hf9iBuC9
+gi3kPMj/OjPwUvFGWLjWwCsYncHWUFKQX7UQ3GtTAsBaU23S+DYNcxfMG57DrTC
qZnIcGltc47EgKoKHvPS8YvaapgDpFzzRwgeWbwACRY4cZMspEDNKSzzl6ANuISm
mTjqUOXrE/04AybOPT7R9oRTVFKAj6rMnS78bcVcmwu8yg0DNqPHVcBsTylNwq9I
GSYfGiNA1R4sZW+TkZFCIvrP2nkIIW2miWAvq4S6fMeOiX5VIkU7LmPb12J2OWB/
jIvg0sQeNbSBmdfRc3tYq1J4MxDq944oFYjuT/lb+N0D9BQluy7vgTk263QJqOm8
qknuw+DZf1fO5VVJ1JMssWkzB3nrNdvk7gooxR6lyYC2rYugUKLzrIgtBVS0xEEq
goM7M3NesohKSa2n+oU+lwrucXIdY2mKg1pTeFnXS7E=
`protect END_PROTECTED

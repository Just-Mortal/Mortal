`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SLaMUt8LjkKJiOhA6yqujw6+8rZZUGIiB7vMye6YTaa/qhrsK0aIY7xZc1KjDmz6
OvET/Nno4blOdED+3Ab7MWR4jHgIHqitXqEu20/ZTya+sx7S1151NRwaRvUwr4uI
G+xZAuW6f4DnUwkQV5Eh++sStHYm6uzmH6EFhXCBsVKMIGdxN69eciUCIOo+wI0i
3HnQJdScs4hubaYQr/7IhtxOB/BQTyn9BQxteqlmouPrF+OqmSrmfSHg6FXUfb8j
9IbPwDY5ooPYZZEH0VEeyr1u/Pix8Ke8TX1awgC+DjcQEKx0aM4RKNCsVjtoDMCk
5VE74Kd/Fy28QB4IBZhaeDYNKzs9+GEpkUYGv8o+mxJVc/l3D5m6yfPsuclaXSRn
g0SYdnHIBlzB4md9+O+xa8PAfqMSSRt75/A2H6ht41r7LDAw4BWvG7fw0E/yZRT3
M8+pgiHmwTglh8Rhla2Tpn9WLZOaGqH7Q9ydCX+8LjkqtE/m7+GjoghGCy6Dqz/0
k0OfaVL2kK1p+RCMQuBUDDspTVFqT6l1EqsuXYsEfsbVJrVXrwYdP1Ci0GF1sJI/
uhB86zCRHFYaHV8IkeadeUA9ntV3vcypMY0Sqw48j3v3LkLemq3MV8xXCYSDxbxJ
qFMl8bAfG1vZSkiqQwTaHUXltO0m8J6m1cVlBPLUlEFtg3lmS48dFZdQtjJbmtge
GH+595+NCOHdrmSdudhmllQA4QKfhIrwKhZ9yMWFow8HWUlv+awy5ak+KLCCxs4Y
63Rn0MwukQc3mrHU8qR/UA2L06/F63UEsYC6KsO8y0Xo32QAtHsmrtVSOunrpGTS
aaR2MyzYsai11akCw6UStoIfouXIbY+d8BCwlnahahnnD/0JbUNy8kEpFylvKwne
6/oe3tdts1uDfy5ic42xzAsQVKqHvr7B3ByjnbifRoFeWdTfTXDqW+SudbyQXdhu
R9WFaYy0auBQsJdIgebeAOpN3XYOqth5s4+MKy3fwYYgbZueKCPOObxvy2SDcexj
+pDunJv/QKZLqccGbvNURbdZ0AFQ2pLCaRbqcUF01RwPn1NvuSJG7bisBf7fyLp0
a9b38bOsSnlfMLUw0lxUezCuGXeTQe2kX5hvZk7dmn3pbC0xz65iLuvvcrW2B90d
EmpbQ99zbydwWx+3rOQCov/gf7/lLd3hjNWkd6NwkEppXNXWgp9LuP8tqOKPpCxn
4FZsC2eUnGPhZQF+6tcEpWmB5OAkKtNMTChKYClP70lVhE4ITmf/Modvz1zuVTrm
JH075nC2ROiHKWRU+ckegjneEYoCizytsacAYJcqjtACI0PCMSeqacmeAMm1mCmH
v+7N8Rejimbu12zoiD/qX26q89RBMfP5bk2jLOdAdEA9q9dVtq+zcEZuzNlYHOin
ZDxn6PaOGTDtg5zRUHsJ3nYFTJQe5FhlQaqdVEzOdFc6F4e6AQnRj4+MMGMJor11
z2IJXcnWZhVRw+WpO2PS+lfe8bWfDnxXkUWsOKaW6JEbkaA0V9iE6erqAtnzzkmo
YshSrMm+XC5ZYPOfq9LR/oArV1PPOVL6SLeyOxrfY7BzdVq+fOn4UOh+n6GEu0bd
9x2DLC5xJ3KmwQ1lYShi+G5VQSq06QbE0wx8TJ6hJY8HwpMOnIgKLwVN6yjRJUH3
wh4hBoWJ44b+RNBydmjxCkyhzCHnGQOX8pIYlGrf92ATEgN0DVq6zWYt4En23dng
eB/BPeGntZCZBFtNzPLtfuegmOQBROOJ/By6Rt+NiBedr9wBRW6uo2Zv62vtl1NJ
LskSY3eXe3SJoywiFl/VTtzNl1EJHKolP3Gm6pDDEMC2axN3zJYPLjSov3q45UKK
3m5cysPdxrlXGPee37th6aIFcUx0U3z124PXCBO0iL+jQRRd41tHdpCm5DH60KQr
Ph56oocY9n1hh+wLXlCtETATkJuNShNhjg/TV+amZPPN6tGtt4aw24Lq3cyEoPIx
AohRfBnYgBqG2byeW1ZTdrwvUGeCOMmUFFJnbIM8NpPO20g316B2IqSn8z0pdAyO
ZZ9QfBzySNrvfEoA/i2Ct55b1DNiWJRWu/J+UCyoXSRFKK6olwFmQDQ3/PdO/vMO
eBOwaDREqFWbHWW7XK+rd2PVuYo5pDnhLz4SqRmfkDj4hrwudxKIFt1yHFT+nG0E
ZtIOZ5DNt5c+uiih7sFRs03BRCLIf4KBbNonFrhG0RDGgU8FDADm7g1aLH2msmL0
Kv57hadLq6M4D1DPIVV8oGZ2wgAFDDuSH28bC2LjbrPg3j/SKECgiRVbF/7KAos9
bCNJYknuGv4nqQi0lMfviFu1n5OnlWgYEOdHeGBsi1/OCsTwqmJh/lSlh+uR0BtI
y2E/9Nz7dJzohAEqZLutr53y1ILERjsDkvVOHLrzfsiGVjtiohRpsWjuGE5DPsAW
xWVZB8oqBnz/tuAN4kWtkN74lMXm4tXHUCsxN4aRzEFjfu8RtM4dgRseuDhXjML5
GRCJw9ZKxijKcfwOY3Jkdd6xBGaSe87Em3i5oLiUq+zRbZP/OhWzeslQEzjlLFsM
9+5cY9QrWTXTfZ2JvBk84TmMBpVKd62diLmKMZ4cUOo8zmt/6bpSHjfPBrjiuLmq
/QHkS4TWp9100NBSDSianWfijSocAKTo3YbMaRJiY6p9dJpRfFeD/4QRdMFw4Yl1
CerEHe7iL5+m5N/2Rni5Xs6kDLjBhicqraDTSeW4zT+xnEyWRdCc6J5VKRoWHsmE
R1tmEYnP0BMav23Ai8JC2h2OSzFKZs7Joms/CUmcCe97yUrjfK+ONORoSym0F6Eb
mL+Wd+N61O9UPjCvya5KgFXC5nvmcxRBTEENg++ksj2zzsNfj/r917QL67+lSe2C
VJfgThZTOWktOyv9V4ncdDyPlxnjaGEIUgtJ41g0GlC2poLz9/zcI7/ELQ4S7OGN
GWxu2ccrq8qb5Kbn59f/33Fn8eWrf2GkZYDpG8MyIEtf/i9GvrowWvCxF8gFcB7n
TbI9D3fDthrh/TGpEBUekHFXUErzUCjFe7eZiwo/hozgoeX5x2JrkSQfxK1NheCJ
1711eLfMUgmQ7sf2IA+DZ2GUg/WJ51Zd8K64HzwQo/kAhoTL4nDyT5WRoQD3SSaX
0iGb1SKNI5XlJTX9tqq9FUsJvQHVf+RsntRD6gn6y0zu+aybfhi7EeAz1+7QMt+z
D8rLaAezj5Lrc4lDMU/9gCqdoMNV1RDpvtKjPRxHEK/DqkGdckBQSMkXg5IlqrK0
ZNBWJ9N9e0CGGUmNiUxWDURGl07BbT+vlo+eWnxObuhN76C2uvpLwBRDaU7/u2CT
HJTpESkwzjkYbKVIfmHtB/tkcgWfeI1h4pcic2D1B8WPQ24T2JamaetUKpFGOmyL
tddz5hWNNdTnwftizG1YX5mf3LdzJNXhZTkUEh4xspw=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIomZHL6/s1ogJf/Sd9o8MA14m6rHdsP9evbxadFrwyiQI0p1I9nEVIcZzWvylrU
92ZAJS8gpe03nacw1DJe3o/8JCaewYsX97LOtruihHH9mmrAybr1Y59K4zoh+ep9
7o41h2m9EDYbcSjmhb0+C3JApbH4vKjuZyY8bihg3E00nW7grYzaD2zaEW/78+mI
ux1/GlxRnZHmRo6d4x7Vfrrqw+Nbpomh1X0z6Xcj20W4vCUKgW6uV5Zf0PY4gpCI
tM1GT6n3kj83VBaSjBHtZQ4kHIkWO17QQTryK3zfcKWJGgLNa1NjxcQ5HtdVhJGv
Qo1GU5+Dvlxoc3+1YSbD9C11S7Lodzy5C+auGAuCY0nkK5v1Q0uaLSzRP0TJTAgW
MlN35Aq0V5cg71iWh2OwVIW+LwwwKeWnlfThtQNgBq+4rQyYZn2tidQwkQEP5hky
b8ExUSenF90odncOoPuVxJJdwwyYlNfhAPSvuEPLVoRG3CHvPVYHTddexZReKPq0
DeZylnUGI1PANHTUX61XmgwmPKkgt8WzyEuUWjutAB91SttIkWdrs3D0GztdO/6R
n3+t/ovnxhsy3J4W77UHHypXZEZJo9nd3RuCmKHcOo9Sblao7OgSes9IEGgxm5a+
HL1AVti2uiZoAGf2wXsVom3d1O5V/LiVYkdL2bXltsSqKYcD2VndnQoJHC1HLZgT
ZCSVcHM01lOplVJXKq2SJm6nVnWm5jKpIKSU+Yv62yH46G2a+QAAFwSfoBgdOJbb
qUl1ym3hJXedR8jhIlyJwSFBrnV6B4PvkVT8hKxktSO5cDoN75QnnnAjUAvQ4PhC
b0uSKBHe0eyVewMS73lh1CNA9EHFyFTbwLPR+Rqo14FhaQQd//d2sqz5iTsfojFl
9JPzh+H6Tp/tRMDPV6qe64MnGsC5mWPb6KCw2abCXFJTqPo7d4a5MFIX1el+vscC
rTKPXr7lBPNRWWHYvvqX4Ud5EtggtdMSCgmEQJ6rwWy4oXXjZP1V3/BqL1m05XHD
4QiNG/c9C5w+32lA0vd+mFpRdpwlcROBbZO/Z22IzCOxxRODpRZBSkTFS3aaH+wq
SuQucKVKXnR3xACWwq/PN3C/fDUriaWDAV2ZXFOcKrP97sGvdMjGr9GylzwRAOWR
tBO1e8pNpmhA2DXASV2YtjG928ipIrse57NLkt4QoMSyY2y37T38LQbrHQWC01kG
sm4k0DSLvVuwABQLp3kkm4+cRrum7bhsKrwOfpu9Ffzrc2CV9sDYPSFtz3bUsxrj
nh5CWIsRKH9mL9UWLXCBEFSUzof5LUSZ9zPzUEv/bXtdrJs45b/0ySuKsSJ98kun
70gRK8e3euzTV8uyagx313p4K/y7PXM30WcK+lsbVEZUWlM95Ara4y1Ds82Y/Vsx
BIEPOKayYcF00hty2nJvU9tBlVh+ThCHo1IqwEejR4lSICJdYXMmqc+220x5s0uV
3ZFPp4UYW6k491KqfJ6M0OhhIPp22/ATvUFWJjSn1rSq+WwBCD2ZBxt706XBRuAI
ar88JpGACAxa+7E+p5k0Rt9knqeR5mAAFv1gDWuWIS5I8gsBrILrUPo4ksAXURgo
ino6X4lR0KJbcr5CR2MV4LpHZu8WhThGCE5TfVyESaBBBRuXR23lgOm6pFKNyaMk
4oxDAp4/1Bu3XbmurxFLhIOGH9cByeilvLv0SSzij3isphI73nLFAjhqDK6HE2TQ
`protect END_PROTECTED

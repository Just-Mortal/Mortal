`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IqM2VlzKDnMaJzfOgP3muouOCKuMH8+2srnFxOvuAwACB7WPQLUuXIeHXgr7Sjy3
7gR9G/i/09mialeMqEDa78curO14cYo1b4L57o2p5eCDU3UFZsZDGYp604cV6FaN
7XbQToJL/mRF0KDcUIa83S2LLNU50p+KzpUDX7Evymfr4FU2u8SByS6xo2YhS8aI
L+d4s0qtzfyJR4okcaDDiVOV8FmovwK3ej83TUiwzLhIFHcwToxwKQh0XZmET6jF
5Vy35Bt3IL/IG9ZnDcP/i1oxJqlCwLomIxz3LGbhYb0RVdY5tqQkw1L/7CDaC9tP
jXHQdRiQQcB3WSyXWSG1c7YVByxGl4zsE6EWT39iiypNZGjBXUr1tSe75VxkW/hD
zFfnn14NS/d0UMTe3kBqkIkjpw/tksWYEYj4TChFCL/d0gKptvZOaTD0mFlx9ZAp
ALmPOag1jvCCmW3V2+yUWoHFWkzNozSb0aqZojJWEu2ku75hcoR6EEn8+e+9CTeg
FSblghT/5P72p4Xz4rgqlKY9IskKDRapd6IgOSTmpsLaqmPcqyCYknSZmBolK5Or
cFtq6YjqQC8eKUy8E+Zr6sHRsx6C77x0/spG85S9T2Saue+Pqk2AhAvItSrud0CH
OKRzZ3RuY9zeM4vwnoztjNf2EUpbUWU0J6xh1x2NbB7RW0EXDO+H+D8bK03FExru
9/OZ7mUsFiXBaVUdMllyFRXdZTYytTatTvxcJdpe91Br/AMuJwv5vwxcon0Wi5Ua
ju2hFiFv7MnEu/D4Xwmv03AkL5ciBThec0So1xvCiS9ijYO5Cy+RXKsnz4Wvk3fD
SmSG+X51QrOViEfYnHlwa8EgPt7Mmq259p0h8Y23wHA=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txwRmCt4jA2ut8GMMRTTU/GVurras825rbKCDWI+vao1d5J1UVXe+UngW8oI+ktx
RLLLxV4qjhjDXuRKI+5f7Bnue5Lfyj/BqTMkmKXm2PXCN35ups8E1eSGcbnRGSHr
7VZ7f8q2KYm4o6EaS9GDns2hvxGqdjm88gUndWM4I+Knq/Q9X4rT02kYveyfKEle
p+uMxqNYZ3cZB3jS5JkFxufSBnpuQAs8L+yjEvIAE6Riifkl0LYSImJn5eX93TFu
EOXwVj3wvt+9+wqJ9Y0za8WDpA9ePtC7W9T+Hbnr7l7RK20uvXVP2PMFAAHZKE3J
wdxhA+IKEBJ+yPz4TccGrbUAApJu+2TP4Pz6FiIEZsmp+y2s78wfcs/jVjC2sL4e
`protect END_PROTECTED

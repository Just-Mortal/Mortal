`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/GOaXyFiWEy/qfgR12jS0kOzkySMtp09YAspbvpqMnM11xC/4ric0QUQr38wuKK
VhxXgn+oPcku/R4T9QCXLs3khL3kP9MkZ7aGV897OhMbv7yhVUg6LrtEboXFlfKV
6m9U1Z7mjEGi6Mmu6PaoaiUg39ErV4OcC4B09cr76q7rhckFpITkVnz/lSQagAY9
icS5KMb+b3jjU9MlPDC1cP+rZxu0Ev8iYWN7DoH6U/YCyVIuebej2YqNhTZLOxbL
R3TCH4bdQELbP3+oZTUPgIMu12zNISSprO3lUX6pk3W/DTsvCbbmp2HWO7SIqLx5
Wmg9omKexPJnZFpZuZYNPkXFeKrfeSAhQyoB05AiVuJCP8utSNiW8cJZqHytnFVy
1+Gtt4FWPJ6gQ3xtXE5gR1oCtOCXPb6rKnLAfyUCW6EH1Gcs3WOB6+dcs51FS8/c
Db3ktSlyJlFqJXfm9MavtJJIz1lKhfDj2g9ntPjLxrHs0S9WHSUz/51Ia8vL51oT
A67XN5Fi7ll3PPxs7FM5/mfEq29OL23UV41S9OcHK/za+rKSbNHO9k5CFT562eIi
42/FyY/wTSLWHq1BbwJP5XAQClkF4i0Op6MFhbUpWAVFr/VqdHoaCBGqU8FRAGjB
lxOfaQbyNQmk0SA/zEL4Vce0BpT3lzDPgxDK4q3fIBDOjypTAQcmOuB3pacFSrV0
R8z2OnJ97mhedmsAxRP2Qk8osFaRu5IrScHM6Me7vtjO/ka88Nu/NRQJ39/6jYTM
wt13CY7l/07swxWB75Saik7YFFkluJSx9S05SIhQYMOIiLQxDIkld5SNFqcu8/hQ
DJj4To5m94b4PZYweLrJuI0bKIAymHwfE2iyV7f1Ka1rMvNIbH4cq9lxSlX1sxXR
UrnEgVx1IdIvVe0RxfDRiO1Zi6SFa+V/A0RA0R52U0ptPLqv1fOGe3tbKhn09KY+
zXyAqenXG1ZlyRm/Z9SLredYEcdrm8BvXO8lYMLuikt1LQMu1U+0eeYpUiUWuuun
NeESUkzDe153v0fXwzKj0Vuue2Xn6xOIyaRzlBhaE1k32IB+S9L4vHemh1zhLc7w
waMBlH+11ANB3MAsFIEA25bicdQ/NlZNulYKnoxC9YkU3qoSZKW5xbTNaR6WZxcd
j/9BnylKZE7KvjNDIFj0yRvKFGVT2HWhSep/7u62UybJbHZL02mMu+iSP5cQ7N3Z
dDuNEhhWkyZ7mCU9Iyl4u/zA3EB5rJyqZ/PXJ4GKA7ewIA1TlIrhI9akcawhckLg
QHdkm6swn++Lc/nL/sYgTZ79h+1xsknERb4dNxgCz2wwcXt1kOubgHYKi0p8dlHr
A2y6i4zbeYEMl726mLtGYMRh30TB75dnyOAdmQQMqgbNJEk0LzkAvcjJavVFRAzH
0+5oiPlDkv5ho0vcahjVeACc7NeR4trmohKAX2d3J99zm6ZkOgl6K8CpkqoePv+V
QCUIU2CED0TIXdw9uUG6MMu9+n1fLXotoSuIxsMOsoPtgPC08LD7kiAXN1SYwODd
FeHzUm1NNzIJl/a7Jx2Nm8pgv/WsgHHUJS9pAA2d3MpjAbQ9wDcui8gmy1dZFAOU
po14M4x740C11EPxZnDNL1tI/Wt4di6J0aBCmw+Q08rN6ekn/pw9yTQp/k67B7wZ
wmOWwBpYZYheFUl4o6e4sxF50nd14dvu+547VyKWJ8nJFVuRPNv4pvlDUt8I0cKE
k52zsmKcsqDnPA+ztrM+zA1m+Dx6LTakHC1v5WZ1OrdF/jKxGFm13yMskB0k8Bg0
GgLLY9eRKxQrfL5sOIWbtanNbi9s9MHzKBypfviy4UHTWFLoifM+RKeE0jBdgafF
zRqbun08NOqJn7INKCLI3RP8Yj5L3pC+nN3Zu1m4BWdiLavrxprNRukaAX5MFl5g
KCvobX6id4dmdTgwsTdffA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
89x/bfHF5UQAspL8e0hL2PzGPs3U29/UE92bRYS6lzzvjj5dSpAdcBkeYSMEgc+s
0gVKJfM2E/GmVv8uhfcedaQPXkGHm3QuB0MtLlWz59VhTF/8xmkl9cC28q9MWngD
k+qHPZdkRM3HOk1MGfSz7zAUouiFv4pVfLPMOBTTV+kB8zH2fA9NoCRP/sXftMoh
ld4T0KdRMBZshr4OHRM/62moIzc+zd1cbiZxL/RC9PzEENy7ML2LWCtnymvUziL6
6erYEBmT+h1ftUKdSnqP3xVCJ5u6ldsslL1tBNMb/bVlmUX+nfcGDZQwuZMMsrsr
Hijg573hlAYPVMkaq2gS0v5BmbedDeVei1a2D/9bn4lb1EEUAE2huMEexURcEo5z
gCSUvKVH+qTsOM8wGofbY+YWG1GuCnIm0yZD7LbHiy50SskHOiigBRDnmJpv35VH
`protect END_PROTECTED

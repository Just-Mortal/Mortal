`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dSlbzDFsSIPwu2zUi0ZesosvDLeSApjQX3UPgF+Q9/dhFrGE7A0Eu/H0G4zNJk24
+WKgIAcApeMdI4gYW5rhdWA//OdkaxBOXJ3RDoXaih0Tyc2V0J459E5TYdyYd7in
wq4+A2AaP6Si7sX+W6h8ZNF305LSGWHRiYeMsH3fI8CNlhHUsULcQ3j007+zhn8q
jP9ztllDQP7bRnftob2B3OSerbL0kMUdeHQe0G5R5Zgr+EpYK97mzK8Bf43xEpEK
kMhSKx0vXzXyEWPYfujGvvXzw6eyzzOZyzcFN/zy/13KA6k/Q/7xRqvDDxwEh9v3
St7oKO5xJXIo/IXc5GYJ9vyHqEz7Y+GbYcvUZZ9w0BpqPY5kFL/D3sqoS8u0acPW
FiqlzsA4x5cshdcuWRtpMbhXO8rvsrq4ryNomEM2h4fGTIWGSilkiaLoQhNDp3l3
ayvJijkzmJKV7p4fqCSDsFD4pnN3swynaVvaVPBfsDTWSOA8zzRZD8X241ruqoXh
3Biy2gVdyFd1NZ5PbvgBcTI+8Uaq4ctaANl/4VJoAHLoeefZkAT2SW2HM3/Pe5ja
3FZl0RKaVzxtEk4yosOGbnSCFZ+nf72OdX3gUDQOwc7X5Swpqcg+mX0YztqMPAAn
0WpfWd931oRrgEm6XWFh/kRAWa9NBRU/bQTh1k51g82KYPTpn9BeEH1DTOd+3j+S
Ngrh0IxrOxjcT6ZhvgvRtd2SYsSFUCtlm0aSXbj8zwZ6Pqk580fw3izSRp636P9F
CLjfMESL3WdYsOT2hFdscP+9JBSPse8zWIHgx+BzmHdgxPa6uQRSlJut6eC7Xz/4
u/JACmZZtJolic34j7o5uAveAFhphe/3yuiukfLUw5H+yU5YTQM0DjpSQ+LRRct6
qbgWQ89wTTUxC4DUUNR1uco4/NjD03ZzrqzIYpcxnSzf9K+npdnZTg42PsAYqbOk
oogFzyOAZgXye0darz+/xGfCV6RbSbfMpkk8EDgoNvHVkoWRpIBXwfQXj7ItSIMr
Rf7lQgAKvvqpkzuvidoCC1/olanl9NU7SNoz1lRTi9e9aZjAHKeMysADLPdLWSBx
vTRN5ycMiZS6z0tCDIknGKq3LzuW/zuypyAG9hJkRWhZ9v2Hot7BgI3L4MsXyEFL
LpeIY3FRpU6wNVKaU3Ne6wYqx8MI4CLnJkwFgkz4JbY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkvGZquTZcQfEU0nJCSM6xhmWfyvkPeOP77UamsepkkvLEQ9K95L+DMHgH6Dn48e
cFzZ9B0wn5pBqMWxpDTvOoforinp38Q8ahyAnc8cxJUFu6MvDQFHl3fk1Ph2u+k5
1I0QDSWfYU93YzJzhiGY8UrQF/Rdzit8fUDpJ8CieLGlxx/LuaFiJ5urB5/LmCu7
4joAHjM7stQd6XJFer7UAwohZO15cC5h71d9JG/etQOG6Qn2XwNiICta8wiyf3lX
UEz0lKxXbZiusyD9FqFt2A/IQ41GwDjyWsEQ1JhnMGA5u4/xz1dUPeR/uJJDFDFS
/cmf+QWddFfGZByIUABbToi61BE/UpQFmV1Hyt8puaVQjk3MHTMRksfxT4V9HwIl
5eFLpISRJSszzbJxmmoRbWMMqVMYYYuAbQGPNKmdJBkKL9yIMxzhUyNw/zH9SQmB
rR6zdLcpIfJjPO65RcnpGN+De3NtvrbV4CjOdr62m3sYoweiMZ4jbaeBTYxozi0S
33c00mPcE6T8hVNSGbqefMFBdk19JzoA0K2dpf11A0MZ4Fihi5F6186dCh2U0Gpx
+caB2cNmwdnw3MFKEh+wkLZFsgzPrpl3iW79FoS062YtbNPPnLuqO0/DxcH4k2x8
6Ub6UORzcbFRN+KDWsz6ZLCTBD2moXQ1ItZpIciXOG91fm6LEf3tI2bhMnumPDZ4
SBdZ7AOBkCeO2IY04zOSo/5hiKc5gNAVLnPSZ3kgFuzM8k/0qOZTzej7XJYoTREL
z5PBA3l+1CBSVGgLR9+jtbsFYealg3vAaEu5kL9ubtzoCVa94I8MDqJbcJV+Gxxu
PgQNeUk69lF9Z9me9hY5eMkdI4+pSkLqfpy3Rnpom8gSlf28+bijQiTyCIAksbOK
V2CZfUeuy6376qNAkP3yEwbfs7lZTUx6TooqczyJI5v/2IE2vRnlFxhFOemBJj3y
IXuZUHzyyo3X8E9vDUUO6LC/oxbmdHGBsuqHuG7Y20QgcBFVB35yaMeKjYOZLc0x
CSe3YwA+Iv6QuNH2qQ1U2EOP8tMxjDN4OY6+4MFY6p50J0LHjsChb+uNWy7YlIxx
mFK05BoD7Z0WtJMSfFjaaceI+Pip3h1W4+wngfmKIOeYOyxThOyznPw9ZJ+mut0e
5BBM5izIQOhkshMGQ7ZdEZfH0lQMAdymQkTSzASDjHC/0eNYvA8CHwQtouhA02DE
vlic4wTxpRR7l1OvUAgOyFH8V0ZTViPLKS5iMTqy1iaEKAMDWjADEBrsIPEXxDB9
A/ytnxFtDn0UxLBqBM7/dIMSPH1Wq42KI7byNhxLAoqRUAunp02TiZAQcQwCSjNa
nk3IN+kP/BupLXx60ucMIzYzEhCN7w3HHg3MD358BXA9U0VI+rE6l4hVGCfcvFrg
5C1dGz6OFcb5k8A2Jr4Apv9BaI2butajO+MHIveXlcIYGCJt1ic3HfBAWDEHWlnx
koiKTexhTBLbc5+4BoFcbUuCDxZEL9H2ma49VbpUVyFjTVakug6F13u5MZrvdSLz
pJF7V1G1c4ouxS/yCMnqy9PGhPtNgWf8eCZEiiEd3ZefsXwIFZ06m+c+r88A0B8d
etEKFhWrg1AwTVuFq6H+5FEzq/tEGMSfoKjsNp4aY/hFvRV/Z6eML2qq7ewfKTmg
JYmqfa5Nv8FhMnaCjIe1/zJwrJ3xYrtr2zJpLmgESRc/RtENj2C6Hjo2Nfo+Ivd+
710TQEm4ho20yyLscDYAY50HefrmmjXF6cLYl/tKDS8qONkyepQpddoz4cVG/84v
Oz08HERz6bvBAbuB8HhxHxVIkQayxqmgpXmZxdKpsCyyv043V0fP9EJQVyC0y3Cw
o4e4LxCdLqZGSPANYFC8G6pAhuvRk8D9Qb3cMoIgcTR4WHcAco4KojKSQXOyG0Ne
v6ElPpp2uyyOXBX8g/qcOj1gengQtnHjhMNObepvz3MaXicxFim6X1Mqnrs91EmA
dpzfAX0zpxf9RA25hYMTqnLYAOKJbLA311vX6j3Zecpql1ycINnXuA0FP2lDYEEH
DDCsrZsGdy8y7iJ4frsts3mtRPRs6dmwx/RhgYN9LsOg8S/7S9gtO8F/Azb65Jl8
`protect END_PROTECTED

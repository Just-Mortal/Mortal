`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBWQ7XwWBl37ozKR+NXmubQDfz85Wh6jblyhmt46ym4+CiR/6usGCAUmZxCzxRNm
qqEPuQrwO8xKgO0eEgzOtdeS+XLCdZ5Yv7da/6g8Gm+aosFj3ukDTO5YS3Wdia3y
ig9RvE2fy9dsqnwYg25P9JRYfhEyqom9XWnuRUCoY1BKnIWpGiiYKBX1KBJEv1Qm
Ml8QTookWqOkZ/1FkT+6/9BXq/nMboM/jUG+b8epriRDkaiLWIc8iHZ4TMbzlEEY
0qAiCV5TUDW1HzI7Omc3ky3F7aozoFuIU+zwDaWKOfcKo7bWy/JwHIrKV0OGefwS
btVIGpNsrAnWNNbM3pQkOUazCv/szYfeBJVR61wzhRO/ti8oBf+nr9KIwi/eN++y
suSEvkl50i8jPQGq1btNlIDxqJSGBLB5ofYhJPsAuiyOYuYdCQ/dGnPxchQFyRmN
YtHYfPrD1ejsdDIEfO8Z9z7AQgeTQtL7cNqxl+VtvTChaeQlHRS4hCgLMeHdYNsd
A1T4ma0z+Mjp3KSlbI6NBFRXpzPJ4LXW5BSk6+yrKYRSAAXt0zg1OH0X9npj9wPS
1S2M+SJAznb6GmC6GbDEjzJUzPU3RQaC5FMvuZtL9c7mLNIO3cDpTKmKcyMX4jXv
+NZbUbEmwW3tSnxYj30Q49+xBnLGtIQ1d+IWzr7lyps58jJtJeFvQtqZOlVmdZrO
yFNJanED5tXNW9CNCnM0YMk0Ma7aLqqQBHgZtcvTGnZQxTrPoR8ZyMb0tkAMRYVM
NukkPsat8MZRfGs6Ml6vQiwekJTygW+aRbzCmxMvzWZmYISNNrPVgaCjXUxhwfgo
kevPZvqac0VBbk0eeOAWqZjHWkZMEitQLIw8ngbVwqWdmOxrcpTITBy0BrOkDcCj
inXbHx7AAvYzhJI7ERrj6U0Snz85DtJ0V1iQAxdARUgJyoGPvdemXL/xjk/WviUe
iGh1TzbII2YKvUPz4P44ppOV71fURnHPGQf5/hyYLGCtIzwAZ5ZCBcG53yK7//uU
vuSQx1XHa1IXfWwzj8r1rvjsrB2bXfhfYFw8ZehVtuM0H5FRpdsy/qLE04h7ftfp
NGHCyhXfmcQVhU8Jn2CgXPYPcU9I0wu3eukywIHeEzBhcVbfHhgMcPeMQ/c1zVAY
R9bNeaBD9qUhYyW0+FtgnyJJoVf/pdWKQ1dVNZIRvVOjQHw4aAWKnPlaTpFcG4WJ
vRLoZTRRVN/ViaQtD4iiTM0P0+paDXdbnOeYqeYCcvsXHueayra0fUyiz0vrFRMa
CzdDMknAkE21O7y2y24I8g==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YMnKSG6w+QvhpqyXJTjknIqRULY5uRBfzVijn5mx5EvF5hiYv6lml6R5016DpkiV
V+IHlo5yqjbbZMCRNFJCYKtX5xt2d+ANCZRYy1ByWe8w++iV8a4rsSS3HDiVWxj3
ZVnVgmxAipH8JLxiIjXuh4PUC7p7kL+jbedtdjMqH7LIygtJVlWktT8DwopQC+ZD
JFvceL1gA+nMSScrvQb+tsmI1L+kRHP19K+U10C/eoRK+0Qw2u0hPURL9FmXgA/s
55+/ZsURKtJER0tm2ZJwzrTMYA5QArn/NZqmPGDrcuYKtjFVf55dpwH054pKBnjL
jcBASm/DaqOjbL6cpWMCMW3o3SZJkBy6dQCaEOfztSfCYc61Mc6U5tAE0Mp1sEgd
z+YmYTokLlP+powOqVU8SCSq/KtCH9J9d0SmvCHz2Fu1Mzx3GPoDlcQYadq6cuQH
z5cOQsHQ5ClcO4naxwYp4J2JXlcyLjzo46vI28BuseoVcKUkWnhehtg5KbKOXval
0nKBD+S9zHbz7owvZXTJtz6RqrSxLB6CMA0v/Yc2SADohBdTQ3roxHGlymZqgDv4
K+dsz9zODoNKjlvOSE9+kTTs3iADq+MuCs6H8GJgNWtRIiBAaaiNn1TkvTPiL01J
1AM4o8DThbCfujSylR8APT9x2bIt+P3+t/b89TniMd7f8JYyQCeHBQ9dgomeg6DF
jX60XEegeMdjwC/HY80UtRYo5kFwq98nLBt3Hpg/n8ob9FRVi4P065MkQam3zhaK
/xOJ/zIi6KcJMupg7ous0LNLBK3XDpjO9rihUkt4QMxIB7YfAiCOcBguVJF4CrNs
t31kTaVxKN67gj1dqhZPajwcKigHxDuuFmb1qBvF8jCL2MN3pRcFQ7nwGkuWCRAD
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4vSJjXHUFVCPNmon9giBxL9ny2i9F+miqeFmAHjkCPZbePMbNMkupR/pZLASk/Yl
6uuPDwuJCpV4nMjSghq08EParzVPKd31V2enxV1I/gnVPJsewQ1W2ZexEy5xCaGL
G9QxNgwAL4l4GGhenKSvH64KJeacsqe9I4+XKGdtjGMHIUcjH50BewH6hTOyO9es
L68RloiDLNLeU4AuJIRHS9tNgt1bK04MjH5OPhpMkSk3J5DN/nwwghh+vJ53LcKc
UcqkcebbyNgTFl1pX9gO31t9NNcLoM4tCA3PZy5p75nQ4Mqqlb05FjaPXdqTOqJk
1e+wqJZRl4wl/99cHq4GPX/xqngluKsSwP5/19lr/tTkaqRA66sR8AllDhnN/gFL
V19UZmKF9MAwU2gdgWzXZVkCVMXZuu5DLJSNhNrARwsMeZvFy1AA8m5dTDOpuBbB
V0KzWyJPZrGkD2pW3UnU0ZH7QEYkVqtXIZ1+NcISYnTJ+mh77gEwWDFqoGacjy7G
rWKsrxYMi4iHwg9N9PK2JyDnCs+TahCJIirsMn9RR5geAnKGtPX7jMOjaDoPK0VL
YaPE0J4h9MR4Se9iD8dGxEZ8uBJ/sSEuv3uK2vXkt30YPlYyeRJZmH16zzFCPwO4
4mOhFUU/L78uWi1k2CBO8h+B6LrFKuoPv5KpXIgWUbEyh9Ao2mjlf4WDVOMgmKRh
/Klj6aXHXgFP5MOzPfrr3fkTRDw3qKyXEHIvOyHqHQm6KybviIq/fHJ5kRm06Mmy
r9WAjsL2GNXAMrnwPzjoyMEjzv+9H5Mkt0mPtQwxQsorOIgFsUfvMXizlwyG2Pfb
v+bcBL5+SLAFakwp4tHH1IhBLWPO0R4k8pHT7FPkOy3ynFCtid6+bbuPK5wD4yih
krJFxIoEvqFfeLGQxytKfakCUQzzFqMa185VyXajE8l7CDn+zYQkj10FB34bwvXe
L78SAtL71j6rhzwexojdkFfu7uX/42th9zVDdATdQVDOC/8VGGF1j/nnJL3EsGua
tLdEflpXDGcuU6q2YvOKyNjAzlKAF4wfHWGnp0wNXLBu4nDHwFSpApq8lfodsSWT
DuZcXvrwLMA45l9ivs4VitpAoGcAkTLQK5bysEYE80YyDeUpbb59VCUH5jyzD4U3
9QVB5fT/Kkkz7n3YvGzsbqA5i3MggCdFUi00GLm/LnOBZXzq0E6Pg6T8rijVejAl
QU5EA7V0Uz9loT/2nlAzwaVuLzadSEg18sLAonBW6CR3pQrCUfW9jOKeC2AqZEyf
RVIJ4Z4MBd6KpEpbfi/hNMvpuyYyID0TtHn3Ar26tEYMgHMfqOUzIjnXkTKTVV6G
e4lQ+l0A6hMwzEaSeavw61xPiblfHkw4wYoWM1QoNi2+tHf3xeT1xn2j7HEslwjH
QnwWvvLWABADUzRT0dGi90bIQ3UKucMSAPMMnB/1L+/wFsfGgx0RLeSwkAugbSzo
LLTRD1wgEOWCN3OEzF2sbVgeRTi3pEGseZlSWnq0oS/uiELCMJ0pVRIDvuS2csZH
8k0OVBNMLYa7hH0XttW4oGF9JgV1+tu87abCgDoy86O6uMXjA2tl6pCVvWwNwF/R
oJaVb9+3b1RyS0LEEbD4Bn3efE8/eXpTBvzLjzuvw/CZGx7wM7sqZ9cOwUqrVgiF
XlK6eAp2/yOlGvFGcYKyWlOKWBwi3FMbqJNkbJMR21IV0Mt/Uqfj9F0rPIIcrBp+
KjkeiVb/wNxMmjLn4uEuXLawg9ocSII3GfwvtMm2qFt0NaUuILcfUAuAWwp3y8A9
pRddQjG4p0/KGqvK/3dC3jbuHVDV53QorvYdy28VW04OS0V07X+0VtatX03h15Sm
u1drrw9nb3Ljqg331P5/7zjYBgwX/sWijKz3BCKygZxIuUVTTJ4y+e8coPBSXEun
aE2lvuQxOWf5ia+oM1aopGK5cUZoter6kIxvJN8d+qIBQEiX0K2Moif8NDAdeYfg
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGxpPYYw5HkKBDI0AegOufm13M8LtDvtoM4cRwqy+mhhPqXQ9XHw0H4PxNSZclI9
1RJ4gConbDF7mK85TCiXL7cQtxHtzGf4mI+LnhRztvzJt7npVAX5UMsTnRq9LrFm
LmC6vFfiosgGtxLC2YZbu+RPK5Hu9KnYmuiIflsJxFivMVTMO7x5xJ10mb7e0m4d
1EetcWoFZos5bjxvYIX/267aZWnQMdpUwWaSV1gb5PnbqGYZufNjZ/ZW5qFNtX7J
t5KMEeCKPIpweXGJGzxvQKAkOK+08qEcZksBZROvaoAXGMv8z6qSakGVziQR0V6V
LXX7r7hmiwxJmHtBVoRk6CRBCWN9kOhZquDxXWpQPM1ZYwfnLQqossW/OriYnMpQ
P+lcrLPPm4YjnNvHsxVQ6/IQW0NstzPvYuZHlvTdDS/hBh5Pb2Sx8OshCfad2JZM
paBEVi4F2jwvSlyIyqEkbGDENgN63rONuyRQQ3VasSAxM0MHXB6d+unensYfpuKn
SYy6YxnQK2qYjaMqNS8D6rdAj8L5Q2Fs0ZsIwLf0FZRuSs6LZiCyj7WWy7CSrcl0
Hr7IxCDF9PKlJhhpd6IaErL13tYBCBZCRiDVwl1wnVOYiSqczkARHe2v9ZdUbyuB
NgoIpubvh+2LWCMoBzQ9pfa2WMnKMgynx87C52yVIjhUcqpOictfT6bda3uoYt4W
0Et6e6UaJj8NylvNSUfTVK1T71kJRS8a+g/KQU+pJFXpKBOK3vkLaKMRDcWi4VZr
9Yq2wzU18X3GPgJEFlI4Uu9NAH+MYzFES6ofGNRT1x1mkMMNpuIQxBMRMqdmRF32
E6tXNqmmkurquACf4CVpJ4aM21oZBztIDoC8fwSYtrbwPjSdFL4toqnSbDaDaJRX
B3ZHt9YI7Y3XCycoUB05DqlhPZvevcN3+9Ofmzox6NXyknsug2I1Lec7UkNEKqd0
iBjzaUDA84ia/QyOrRHaCUyOpaP2eHof8ZhqmLNBmDu2+kxHOzE9cQczch/a21dq
HRikHK+RxuTyN4RS1JuBywL2VOz6O1PlOfbTsmMKbAxFYKu/aK5wqdq0BtOBaCsu
GNC/4tWvhxnNRIai1Iv8UUNP1M80nh99fWewEhHk9zGbjDMND5LzCJAWc7Q5KPp+
hDK0hg8jrmZpjiUtyaWYbjBUy+12YuPUTdUiLQB2601cUMoNmFTuI7YYXUA1GOkN
Yu3Mcey2IKcIeD4M650eDDi5WJjXdZQ9YIdnXCxSmmsa2MUTIM9nFyXRqwKwiV9l
HnP+tnhlyEoJqWLlzypCH1LkT3tO3MvUTDlM1qJSSZQiPxcd35H7iSijb3TthbJM
1jN5U9lvYuL3MGfFvjJVvW7yPClpA/S+5Wpzcy1PAwWreLnRkVqVWLKiID2fCwSE
Bfls4dwUUJpCeMxrPthhnyKwV3g2oxo/v1DrT5M/RgxRzsouZpqM6ya3X50XYVj5
tj6SK9UGqivl4VjC+i2SwKl1dnXnM04dYPwpkv2yUfocyB09YzTkpLF9nAqC2kLP
lUMiJZjUHOo5ixRgsTVCdEcRQYE8SYBd5peqctnAaHgNiTj7iDfS7/hGnOCFQ/et
MqmOkUlLFQ1hiSKOaYhTKCuC5R24sxBScNXD2NDuf3UnnW92xHmWc5YD/LWG9Kw2
Bx1I/Zs9ZdWZ7Uig5EHvM2sPfOEVWmXgitQdkEP36sduOalnAipGi27KObGHeBCe
lCHpGNVLQ4+oDQymCXsUD0IhkF4hG2zJvFy9uqCZBQy4JxxsQ4gj+4Twvl+VjrAB
JlbMOLM+VDWGI9IhHKNlGB06Ob0yGIV2Cjda47bWDXj335J2aajS2PRsacLxmKqe
VwbIfLrbmuK3Ck7Dk1YV3xXkRAbozK1KrisT5/+r7hR/HjGTR9oZ9WDYDfbfyHag
Sh2pYMhhSsiL8acU1oyMDK2i6swTCYK8iLzYh6jiK6Q=
`protect END_PROTECTED

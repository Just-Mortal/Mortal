`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p2YTRRg4KuC+Nxv0IdYlNOFBmchbrqrxqaHmap+TQ1bjEl8DpPUsvoY0+DxpOPxa
PRlluJVPuosLAvLkzCM9GYaFq8FAkKHAC32dsoa6ldGFbQ7F6w4LJPDW+BXipx3d
j/EATeOQ0yAi2ZrYgYMNr5sGg2n8u3fz0t0L8bVyVpNbP8m6xSHH9SA20Xp9v8VV
Bq+/f7aeTHqJhwkucUhQAVExxLQ1Qu6F0Lor7gGQIhNO8VVNbSOPP15/Fg3bHrv2
Ysr6l8QYKTnJTXklk6BdryRICEJwpKqUhQx8LQy6KzNnVGpK86TkRJB//qmQ5ISO
Yoeteq3MO7YDwG0sVud2YXeRC2Ho9aHNwESnFEVRsc5ADPkKm+4qJQr9A3vvX+Pc
k7wgbnTr53O18ylQfozFtFzdS9EJ1vxrDUs+80e900IhD9m1ERP6O2YtY1OzBTzx
Uw6ohO5hPetQtVaawqnZ2Of3pmWAIW3W9o8iblmstkWlVtLXacwgxHbzltskIkhm
PiwwFnhIt6uUEGt0XBcbHjF0eyFFDhbnsIQUj3LvA9Hqin+Kx8gGvGw3Srj9d0pb
YVMXSINn8AJDKnxTHyT/ph/4uVOeDwK68ykhRAni/v6BO1msvyiyPPExqUk/FM+9
0DQsU//sxOt1yStXws7En4X0TbGnvT7mwA5ujXi4+fOE7a4Qid5qkK1umkLPdgGL
+oDz/YHYr/Poxb0vUg7/QXF36U0DBpyzOq/djKgoahdY/NNQvI8K6H0FcDwuqs1X
Echi95OHn2tCeTVQ38at9C0IshgduX2tonl5xxospgx0kud3EwfPDpFC1bfT5ool
gNGJe69BWZS12c3eAhvp2QxW/qjRGNqTwrEXNBGhRjNWONBAn8pkcJgjhCdS9TNR
2ALBlx+5WDDhYep3S4GYRhrSRn93324u6qAzavYr6YzVv5rY5iw3mcWuK9nnsIqx
m9AyJqtuRNfGnY+8GXDWcA1c47d2FM0xmGFW8epYMqdGNNGT54RYI+NPLYZgE/nX
`protect END_PROTECTED

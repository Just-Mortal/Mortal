`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vv3kjGAM65R+rEbK+qb8q7GqFyKBQs9iAsZ/gpNqCKLBZd8XcZA8rvRMU3vr7Oez
kaHvUl+8WYNQfm7l5H1kYu0alRtgsz08DUQMCQ9Ki1bCxKxViydTDbbxUnAOPBWK
7RgT7FbxVf0MqnboLwO11wgkD4cRJZoEGdqLOkbnC96zFhpwbkt7OqWLKvCACp/b
4v7GyrULQ5ZGUVcfJXGrEfks58R0gEOFpDJy3Nv7puWSPwQ9fNHxzfMsJJK/CoG0
1FIktafKbWFmaNjUG5iWHDKUCzCgysuFe6GlGOT0aXnssj28nlaUmGvEuwQvEpvb
05A8vroadGYsid6nZJvkp2PoWdEOGvKWPf6vlO9AER68DaJvPA7eYbzMHJEF1vtU
K/kyJBLIuIRvKb5BxtukYULVgvtCbZX9FV4AB0Z8M2sm9RWbs15SBTRuwnC8M7j9
OGa9jBk92c7PzXtb2guNmX0lC41fEwP5Dm0rq1jJfC1NXoBqYniPwxyU3JIuIyqa
4ZRzF5w9L4LMoFOlH5CTWjQ7G+cbJbFrhCp3SuO24kw0rRtcCiIKXyffe7gkIsz5
D8LxN28HODrvk4wyhw3wvGNAUM55Bauf+8J7RVT2mQo46bF9UKbe71PQWbISEXYs
YHuFSBNzu/61b76guXh283WX+MWxOyz0oIQP8BXl5CXTwEA9XMCGxNf3s6nvLZw3
rfGHXUuUj3ruoqxNw31hNIDENzY6hKyvM4yyU7+U2Z4=
`protect END_PROTECTED

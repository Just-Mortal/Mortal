`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/ImZXrS4niEs8/bYk4hEHlB20BquA5ixMddvXBgaS+jF+vozpxzc+zkOUbUlUPd
RxwBGM79AV4pnZOpI8DE65ZdSUY8SmdVGmWICkr5FS+6zu2S3S42kzoMs7HNMRX2
pYac0UKkvaB1dW4Ddi09JJBjQ16Hcgu7brULXJPV7VduEkzRXKq2bkk/Fpv5Gkyy
Rs5bUnyr196Bfy2vn6SuBfljyRsYmI3q8TFAtqCmNXYWdCPzpPDn4EV2DA4mvl3D
ZE6mspaz3gJgb0Jsx3nSy1IV3QTtv6b9JZYR8wzwawMI2mbSMHLTK1Qozjq/GrtN
ylS7rsiMAvFp0I4q4IdWNVDzuF1NGbJgug32yT0nn60Sw2T8NtT/57IEcpE+dwv7
FeL0osWFRwQ0JBqy+AknyZZvpas86cneKvczuK2ZD8rPoh0VOLE0xV0xh1jpSlDX
cTtrVjg9pvjUdYWFgr69/F5XxJCnBQp3IQgWB5VpD7IGHTD/4nlx2JFErQllVA1b
PWrBz2PK1T6mBCwApV/Uc8kXZ8EOTXmKNKk+FxYJcHlApWqxx6SiaWoCgwyOl4U7
IdAlbVHuonbxlAy9v1QRKht5+wuwbICf/A3Zh/51iAnyk+O7lkLlckYPzGmVRj0x
5GHI0X58bpddhaIeEyDs7Ha6cN8vCXMPEfFTBMQ5pX/ih0FR5J1fvSMqxCV5VuHW
77JHLj7W+VUE2PfC/QHow2tHlbPOpWRYOsK0pPVFWazJHMrGuYFYimu0OZOwYSwu
SS3eScWaNGUFcLsVolRuPgSprF7ai/xjvPvUt2bLFgbkvWunmYyCHpZFUE2o/K0g
kYq/3cDfEol8JnYbPrWdL/JFCMCnQHwIWNZvcSlFCd2nSD/VMZhw8gWHObOmtj6h
UnRzuYFi/n4+QSKMuUnQQlfVWbzfuZ4zhi7qDJ0aoG20vvg2WLwUdoxSQ2ByVbeL
g79GH2xVVf0djMnejFPDyHMk+Psa3tRT0O8FIVMofqqbVrXrdhNEIk7T/Z7lZp9A
QpThPWo+0Iz1Z1L99ngilgoCX0SM01M0dd2cW98r/BPI9rMK3g6aF9IV83HeXBtF
+WQrqg4f1pADnUJu3jimdWwec77p8iO0kyjqKRKVxGFnZ1MXn/pCTVDs57ceD+rH
nIghNlKqO9YtGYm0Lls4f7I0maFL54/PvbGHN484smcrefU3LVsPDph6RGJgIh9u
hJqadvyR5wAQzcaX74/V7CUmae5nCuZEdLSP1+ZLLofG1Mx8YZyx2MW4ZUg5wuzH
XiFN75+QBzwNuXKe7ct7ZtvncxZXjyYo0AEgFit5ddxHxP+So4pZC3yRGo5ZEJYV
BKWS0ElrfiMbgSKcfgl7JRuZhByMLydM4Y3VteGtXSh6dWYIbCuWm8g110oEZiDn
HpIxqhoa5LpkpP8dHbkAMrzwtfRPqAYOJ6zdlvDFhD588eDhAFxWE8/jkIbph00g
6up67CH+fuycTHh32PjyHjEP+vnyNmzkNAT03L2Ej2XusGAU0b1MeYenNun+z9mI
82DyhKKctL4LViT2HLcJXxms1rlnUKQPGgp5BzXTPU/0dGZF7Z0q7ZIgdE/3Sq1p
y/Yp6yKXc/NLkfWpAlf8d7mbr/yXP/eY10NAddhehT7f8RkebwHmpfwyRZen47Rk
J/a9vEqPOw87/0DzqZkGhsHymcIZfvJoyEGPKgqQY5t4edSd4eYv/r4ASBtUt47J
Rb+8vdLWOSG7Y3nYE9uI2svvOlinQMmUqu54QdwAoMEO4iWxbLMsXZo+1ODfJS58
SDeYpIt0QwF43daYsNtDRVe+KuRxi4O0xm5teVL7rNntCT5spvmCHxyHiBEHARAK
SewJqOrK1PUCwWfff3T06CZCuxyxf6gdCaZJbGXVgmp7PAg9LXPQPP5LTg5LPQN9
vcrZo4rJPymnSO7T2v/HY1u1GPQiiUzoFdL/g6S+yRu37Ldgc8eexOXVYr8t5OeM
KpvrmWOOuKn48IPqdMmpp3XCtroCVm1hZpsHgeNLSGPMIS8Ve/EhfZZkZ9pEotrB
Xo77OS5Dxn+0DDAA+S6Oy3RdS21gv9caP4xwdeldHzbHx3B9MHGrcC8fe6WjRfS5
aiGkrqwO4vC4vlMWPz7KGowNZfrMIFlPUvJyr23Zqwttcev8tBdkq/z/Onldx7fa
UdwT2Ip0C/kWmgwWfOQXv8FSMI9YCBJ9pSt3Oej0GCZMoVkUOjYmsZkJcZl0lF6M
lEE1J838Po9EjGXY/3ZKhpt5v5yQ9zKD8gF9j66nRZ4PWS9pacYbZ2Owk/zmtRpV
ON0v9AHRI+kOTV9aVCzVAu6xiM0rv7uw+UojmJ8fsgdPOPzIIPRDczvfOQInpHYO
SMSlDZzQ4QB3OGuju2FyQElioIkL9TtpSGR/+jWlEQ5v69Gn7hQ5zeeWSxGs0BLi
t86Ayn/TExMpeX/RzvuqO5gphbVa5VQt7dcve0/XEJSFLfhum54F2KwS8r0+Y6ry
khO7N2AGZyNvDTcsrd5D/vjpZkYC19FLPwfBARJS9GXxetM/wf4zPBCrwzU6wyXR
csV/jCBLAmORN+kOY+DbaxnpxH0ZyduMI7GO8ws+vtjOC6V9TTzNntBNoH9tt14/
I+wiIavDMLog+i+9PTF7qtYQAeFEl5SfkOta1N694XLfjdXDQF9dq/q76qVduVXq
9hcqMHWO55RNqkg770eWZuSmsg5gNtTe1AEtKtEbtGlCVUv6tAMwsI7+jFrmCz5L
Oy4jCG94IT3jKV/iBstPe07eOlCfyIGyE4W0DYfOooSQeTZdWSKQIucxIRvb8ped
wo/DZ841YjFYjLoUkkTdAVA7+yMgPAa3P2z7I+ZYL0yg0Q1ExhULVVrJwYsYSwZq
Ga+awlNMICI1jFV0HHrgKIXYH1C69FAYGPwBUCYGCk2FZAPDKKzh2m85z4P+zUkr
GkszuWXBzTlm7ex1ZOgIrcHGHNbN5Kne1s4rWo7PHTdbLYQcZkaInZh4dVO0JtNW
EexwwqDKGYM9Mh24AzfW5z6dz9xkqwv7H21hQIa8jAJgoVqDTMuV31D3uL1CjN3V
Zy0hP2sR4UsMF9BVg5Abpq7L8kkzJMkRxRX/sPv9r0ae4eRwPwxmPwYLqubfBIfB
aQ5r7k9nPkEYyrelTkEAx3dqKh6Ev5Qz2Y3F4bRslZiI4HJvEYG0OWw6P2uAzVxb
AQQ9kSpOzjC+6bcrFBYS0xW+bFYIOghGv+iN98MphN9B/wGRULHt7SZYc6oZdWFH
Puy+PHAvVvtQCmxSAbBEAFpbIRyPakhFvS5nmcwh/HnjGi0qgI+PmhqxQnbtayHH
ZqFuEyUOZrbKXOJCICA62Sg5u6GFo0Y3cLbhHBQN+8NAotRWWSPNqsxXOrAFA2+5
keHrLf9JXhXHnpHt4pMIyM514xKXUXa9twscSx4JDHXp79/iw6FWAuROLLmhpMPR
hZjKe69QK/MZItoppSD9E/fIgl3N2Hi7Uej6cCaUELX0Jlf/9evO5sN6NXu/ZUKg
mDqTT+IKGQTdTQP3YViI+Qwl0Xb2WXwDIYZxVpb0OZcTPWW+RixI5G0fDjBugW9r
i560qhtn60OA14ENEFWpMh2oP/nPJqCy3Kd4sTH5Nu3S/yAEc6vyGt7qrUs7TwbS
y3WHWyvBQl0vl7jgj5jkqnTCTwvX9jBz8BTXgcOwxTJtzvdj3IZCc19sahFSkQ9c
yp6t5QnXlfWDUy98xz1TJfIHV00bcC/B7LbAGvzlm5iCY9urjvNZ8awv1EPmGbL7
umdqf4YEWWZWjaJ055h7jFtrowWoDbKHHkDaRjk3iuxVEY9Z+r2XE/EYEzWqJVcU
TdfTqOcAPj1aA4xalbrs/damxC97Zo1c0EZvGYuax7AC+Mczj822FXYFZowy4O/1
DCfN5VZMC5AloXQnRmFjCuYGtPUrFgNCreLFx7gUbW/x21KCpxMJxA4assQWClge
l0VB6HSvgm/bIH0HUdHf9TYAbnRfmlJzfggEkXtypBvVTzYVbPSLXojAvSy6FjVQ
0elS+rNuVJnpUccoyyDEZOUqLzBvj+Ah3BS7tPP4cYulBieR461+AZkkuesChIaM
19myKFE6OpaNyDm557SMjTbW3WfwczPPM8PaAsqyVvecs1XopnPxPx5M//wG6Bkc
IVDbEXZC9tbjpJm1Yc3doPNBrbV496tZB5uWfcfvp5dL1eVpfUXroTCLLcnIVDTY
0vDUWlG1628R1xyFLOH1zZBPftmuFA5tAdakj2DJAIPYBzDHRj5HnqxIq7JAqo+s
NWa1fUOwGtoNiTCx6Pu1L2RZbpzkb6chle9oNYv5fZAyEPMSotifsndkFKoplIO/
v7NvaOovNO0LTDTlljmLX0OUVx5+Qkv/FfX2hgIHOUBhZcJ9gzEqkHrOls85DcRq
rBm1C4d6L5vUb5XEsDedZdKbJXyMjVdJrXJWPHhHzHYruiUppkwKU2yt5CgnbaV0
G4h3bySueJY4BN9Fu9536wiRN7jr3IGem/2YPwZaupH+ld6KKmGK+cppgZCoHbq8
SCWI6cBvtED1OYW1LYQXIGuU162Amt92RB1IO9xszn0Aw509vc91dsnhN87BMZ3h
xAmCz1SXrgbM+CfotzZn4ok/qe/GhHaUW+GSViRoivtzUoHGZ3LJ65l/CNnOUXQ4
XRwvUBQF8R099L2oRkj1EqieEz4dmjn+1BMMjBJjpoOflfY5jKrg3JVjG6q0KWf9
Ye8OP8WG+B2Layk0dJfvp+OhGfM7GrPcUJnFRY1DPqAFz3TCmQvLFmr2HmIvf2CP
qriHWmLAHoQ5JkTKoo8tQWhkrgkOUkxgWbbHqTj3Gr2zaaM191vZMQ2O9tp2ToJx
Momn4n+w/Sj0Rwq+CqJxr5Bz5q90No0EENLbDbrf4F1bpAkY6rKQa22BY7riSwgu
nvRAAVsyLfdEygYyITRfvcDqjJM79zlni9qs5dWJ72Drl/kjZxLgqpCRe8j6TWe0
fAFtk30+LDgQ5pg+EjYKYHwNTobqj5xTFYHBCT814vo3EFV7XOAiZpOVAHJeTwBe
O07GxQkRz0U/lX4TsSj8YNxB58uRVKuXT2GkS0CWWF3EyDzEtZNT3ER/cBApjdpU
6FZoc9x3BXNAwyt0RFFzq+6c+1fJxfKQbyoDJ7JknoLdAd9gPS4TKTXyi6ESb463
QJV4Q6N68pVOv25hLuiVgkrwcdkycC7AHmUs3+N3DSoUQnppHgjYSFyH3W0uE1qa
mcmhAB+5kJbqWDKhzqerscvYdV7iwNxVKl45rzLDs+jC1QcHd3usbpUz9+REGkZX
Hvcb+iddFDbapinNN8iQmwLcxXustMmEdaxM6Wnk1zhum+0Ul6JV3ObXMROdoWcQ
CZUz3w0sB9/zvu5hR0CgSG8/xlheAat1ZlWV0E7I5MW4DUnx131wxviNvVY2fht8
SIdROrhlhSHmdixAN9ymdsIZe8qmu5+/o8dP03AlCaLuiJVPvgkM05vn2yrTCWsY
LSpL+KmHR1TWshTQCZm/xxohKCFO3uJsRYBH6KH3iyEdf9cXu4uuGBU2fPr5KmU1
FGoVFLk8l9URdGpxTSied2HbpZPI1Mji+KV/3TlqzNIjBjgACrsz8IAmuK6S1m0E
msUuClLWkNsadMPmX6RZBky5RztGkNJS1pEXQmSDZfPIzLJLYNcRpcmVtMDLkecf
5Zr3TItrclY0yTn5dzt/o/VSxE4skuNSxig5j9iT/8is09aBWGVDiy7IvNIfD8jh
Fa1vZfdfqBZ/dOsrzUFUVywEiLrNs3I/dpJNSfNJlZcCOrOQpMlNE0w440NMjbMr
LPmb3O/6v4Tdh17/ckSfSC53fa1na+/qHU12gldh03XBKYiPAQnSLSVkCJpNZN4o
f95WeaxkfQYlU+IddTFMQQ/1dv4s+f7Ur5jbui63bYgQEVEIQOhvq74qXk2f2eGH
2UxmFTiHcPDGSWxQRnRvYAsPu/eFT+KKIdkB8Kahmd8JMMbLk5Sn83msYlkdIwem
FGmE548nUoaaB6hef1u849r1Fgowoz16BYgAgKbIBQXWKkCovQSL1HILObVW4GPe
j4jOLM+xdloOb0k+Gw7l+P3AM6b47HG+wXl7EnsDRREEMjPS8kfXJcfi/XL7WqPT
mNkfmvZkuwmNiXPRDl10nZ1hIVF5HmgXAOHFwM+VR91g/tbQFPgMXmT8VK3RmXuz
0JCruS5oina5YRpRZqddoB8VTtlgghBTqjxki4v0u/mkbl6qTY5FmYv7p2bPnOMe
eTfSThh7jWle/Pc7AXBRoj1XBosovMdPHIek1Lf6v6ZjUjS6ivRR9XzHQo/8UB0c
vGsZzOwdW3ox/dsgHObHJHG6c6WYax4QfmefC0C0rULv7K3paJJH88Jzum6nFtQe
PzBGldAuKhvOHasCdpnGl2wAG5FcSYIEP/iKqjkqvmvV/JYCM2br7Om+gjW03+QZ
8AxmOUhGwWswy7x1b5nTYX5P0rtHMqCYfox/zB3ObJC7SQRRGMNnnBGzzT9UCY5I
pTakkanmCS9JTQIN+qi+crpGleroJIstpIkwKg0oCQRVgw39+YMcU4CU3PRPxMDm
jZ0K57IScL+RIFE6DrGwqy+1sgEzS5Bo89VQUuLHEaK48X2GUPoOWf+97rVr+cBg
+zKAQbsNuy62Q7BILOw54jiNqIm95TRo298fEQcKI631UZ2XR8M0+CxVXKagcRI6
i8SApqg/SklharUlFRmrQneQXU7EiutY5J0pmCnS0da73Z+IvHEJ3zyiBBtCuD7I
q0MeTw+dqieOeWEtHnacAM4+8/xNPabhOj4Zv0r9WPEk8piwEt6Uvu4Ub1nFgX1U
xQh6bUDXeQ0ctNPUeCgowccNQN5/x0n2lJZFMsQxXqwPQYdyK6jwRW9eJA+QBwEp
66F47xUIY6ii338gOnOV6zStDszytVbr15pFmXMjyrBG90JESZf1IKNV842vgLys
9D/63iCA+NyoBnieWArLTog1qqvmBswvVM7satoScqmqB5DJ3U8VxVoCrjK4Vu5z
UzddVF1a+T/s3d8cnOsdgDssEkGQHql7X2rR93MEA5p2NgE8Zd3bZKpchuoIhEoc
uJ5qEQek7YpPPgvJp+BusneG80XTzvrTtnFkyGYTYCI3MmFB+DYnhPcQGc7U5u6+
nYnty7RJCRza1vTLpECqJoyPyOPTDT6uLI5s5wR2mLqxF/A01N7BZYQ9QUyL591S
VKWa+Z7OpUsScUwal/By9Q4qAEK/fasa6i6rbX5kVcItaTD7FOWKJiYlDiLeDghK
hCAMHgNf8LNDlD7+vogps9iU+hr+NE6xmPJGfo8r2+9tos6GInAyFiG+igQbqzHb
XBt1pjV53HbOuCepKySf0sxBeCKxuYUkKO5qxy5o99LUEjNuI+sx5Ib/Lf/wYyZP
TqsWVJ9zvnTsuKCS9S2+03oDHIMvU286xLhev12ORHCYAvb6XzqpvihaGuFQPV7p
FYhq21M3XDSQWEulq/c/z1mnEK/x8LkN2eBBUx8pPexqNhbrfMo7Z+q+vnr4d8bC
NeujE0fO0pbja6R2gODBmwIeABkyj84pZX2tvwQXbaLs+KSszX8RIp7eO5psasj/
KMk2vuJeCsTq2I25YCRYHgns+0wZgfpKvxeKIhTjJBADwdA9Ei0WrI7ICkUB9IoX
Z2e1bdq4qW0HhC6VVlvqjXObvOW9BGoSxbznbgOgfeOJt7HETiEh637+Jo1Aq6qA
6GJYY0UsQeiZy8G2276H/KUnsy6JI+r0pgxszdjM5/CW70Ylkzs5nQ7CXebA0Y2k
wXjhe/FMLTmmzq1cUn1eukVFIU3OwrlRiSAAGaL7UxkBaVujoU8gesPvu7hw9dPE
ADLO+kTYrz1fqybvnCGe1z1GGElM3CCKSUudpOItdp0oGODNnjCOhJr4/t8cNWaB
Dpz8PXZHnDa5FGLE2xbppQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6CFHf0Z0QVZOmZJ9d9jI1t8JZySOwEsENjDV4hyg95FY455EW59pCO0SF+P4ydO
vsflrAWsQdI5DXSzjdK7CCeXufDxxjG0g3UTmpF6WTUyOvESjc5ex96Nlxh0ncy8
OeZgmuG/iBcgMJwCh3a4jNEku9+YQ4AvlLjpg3DRk/+L+tAYY8yi6ww34MlFE8Kx
sU/ItdY1JpSdawSYrYY4xHxiWlOnr08kqmlQ/iktdGVX13YpBZ+qo5QoRCc0K7/k
78iX9zEXuiJqoh7RR+4fnqKIr/JSqE+ulBqm+1zIOXW2RhfRydWZMxi+QI4TO9TF
d7X43CkCTz9gLGkMBY48rslueTt9KcF18dYwGAMC0aNKvOVnyGPv2bSMJFyvFX0X
8evSYdHVRjsB6QFwYP9moN2IaGITcfy/BeiIBNfo6u9X/Ho4QWXoQZWiLMENM9ui
4GX0tV7WLe/mGzsoasO4533c3uCp84VhtroIXAcay40=
`protect END_PROTECTED

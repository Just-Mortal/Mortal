`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mc+hDL8alP+/4k74LkfUHpjbFVqv/B0ZaeTgivXknPl4fB74y5Ga2yzEMxa7uSfJ
3goruqigAcbmZZZG+DnyBEjjohjXhx8ZMYNDZ5rUaVL9XD2gEUOfnDHaZJcoolux
8xOAPOOV2fs0OErfMwGCqaye7H1jxv4lsoFTlwF0+c3+3hWknLYLgiwF8VepZCq2
3Gpk6XdHTHvmZEoT/LYOuznxEF2TzzuLEHvPvurbyLFmlFRF3LOVRnrv9r8flDHM
nwCvb8k8Z6PMqJWON10ulBIYXjZT3SCHzT4FTmLM8q1I2zNNdXTYcjBApOSgYM0H
5cxpp4sxnFkV1Y++fPeu2obRmfdXj/xmviun/8gdfx8uhidthOxwVw2lP6/v9nXK
//mA0C75++oWLw1ZETrXQE2aSm1T3F7F2f73RGfEEFA4xH2SxEZfWibNwawZ3y6w
MnJjwDNKneziN1hVwr3fURPQeUhd6wOjx10K0EO8CqOs6gakJrkz8uecH+U63DgL
/NrI1ywryPLLZLKQwPEEaY7MpqKc/xJiQIeR5OkmJb5OCR2xD0dreRrKzP+pa+Xn
dbmR2O3QwkP+3pi0GlmWTsuv5Ld5PJGBOx95ksKvbqpwpNVIWZH2RzBYBc2Ia8yY
gK8M3KRRfT+aRjWXEvoBTQeFEDAcvJFPSNfkr7v8IXpS+dkl6Ro4+NZA592cnjgc
ULsOvEdjHPzm6TaHhif/Tnqh7ORRN4sggI+CgFjALbDmIP6Gi93FsOB17UzNBK8z
2j/+2hnbF2XKu00f9E9I2dn6Qh21L/oPGVTMyAfvS8ycSXXfQlKTg4T8VK9VtUW/
nGsIR2s4bJ3UBCFSGw0FlDkw+dlriJUHFgqHEVgwEX7HlkUDw1pcfgRgWIV6Qhxk
9t6bzDqRb1YwOFQIZvxCyWpd3vfP7txhvhFAZSXiwjH6FYCithe6yZhiKenAHC6g
fSwV14+RrqF4gKVvXsojH+FQCvvjC1W9JICNHAW2XTdUCYEDdVaAbxRzDMxpiGfN
t+5nj73HwZUN9hbK5Ia5acUx0YRp7g4QFIJ9+w/EjraNOSRkwqO/qqi3ZYLToMDb
xM65j6r5Z9c5SmKsvMDS1zu68pj0Qi3n4391fxzmzt064z7SWC5iBojKSB3/z7cO
gJJn/9MAucIuirVWyl4/UGBeraYwEPFQMzfl9KnWIQ0LL+2ISwYKKz0LgwnVpNcg
Fz6Z2OB6gk5avf8mzXbXwrnPGqzRB0iGaGHCiUmFZvC5pXkODWdPz4FoODmtQOeT
eQ5demzDNXHYXJZzg+BoZaHNQSbCVeFhu/NABnCra/5OuQ+0FzNo58CJKmrT81rx
I0GAF+DlvXNocHVYgSKBx+gSNZFiegJSIc2qjNcc0bfaNlUtiUzDIO8kI4vKs+Hf
8r6uFLSvoJAWLN/52wEHXKRtd586niexLA+9zoyMiG8auCSbDiuMDwoQTN5hjToC
swTio5hgZXZwWnPJpASrAug85J/bkJ89Mjbdef7X/kp0BDj10+UUmWxJt3zDRHkt
6OYkfudc1QR9m3fQxNNET2qNCWBb3ZnLltKDhCIuiTiKX+bqps6gYhbd/in2rtb2
wHWGf4+Cz8hOuSa+0HKcWDrO5ziAxZRYutvlwPvhPbb1VoFuBD9mGeAPPGUA33UI
l63skQzVHZ/kHAI75rmCbDDoHCZTvdlaDXXvsrP7NlxR1ho80tOd4F7PN5HIG+Eu
r5GYY3pBY3EIGdxAPrK0oLCOjxNoyTdAU1iFO/Xn5xyLoPxxab3G42aP9rsV1VDZ
6S+0m/au2XdfY6yUBo+ZfaC/mRfE0xhiBA6gEQSH+dLu7KbhpA5+ykT689Cayk+/
+YPchad6WU5pHs1wXXp4MKZTp0GGi0ZWGarKN9jL/a7ELw3AtEL5iteUwDrc5scf
p1bcB3Q9wHBz9YuMFJ5GIPryq/boBqCL1Lp0gRMoWBe/EhYE/AakG6G0gwtsj+KV
hPPbwlQSeqUeSxvPky4HjbSEFE7tk8n3SXN8uKVieCQFJ9JNU1Ge09dCibId7JTZ
+MkkUZuhWpN541Dp5zxkozki1zUNaub/FOqZ88sXFEVDYToWajUcJoam5IxzFeKz
4q54yyqdDP4lv9wqscOZJEGBTSE+H9MilkwfuFddUj6EmaymhgzeBFsHyZPKHlTH
5DEizzfNi3DUAK51ifB27svERAbdmd1EX7Lr1h1QJVMy44Flv30xvRudBCgNUGf5
EQhZx8JfxOyhxZi0GtJCnF0uHGSpgghK2bsyDMbIbibAeW8HZTfieKMbx6gywjZI
ACCTanUNA+in4uMcg6437wm7O73O9TvAnljN5Ab4Ag+8k8pFiutFDV2Gt5WG1Lfs
gYk50Qu+2WZzjUEsyIVim9tA8eQoE4EhsUN0IefpMepWrGKMejpy5uxzjjAWSkCp
42FUEs0AvIU0/sSfAGc4rLJv/3kPrl0KguiBCmAG1xqp6eFQkFWtAWlKKLKuBAIo
9SjLfQjxIQmIYBTqhO86h2GRhO2/W0kSE7IINq158ujJeGouJjMpKWUABagZwtFX
9NAQWtU+EVSrq68fHj0nZQ==
`protect END_PROTECTED

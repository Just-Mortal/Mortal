`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nkkVd9EU5cGKP2eMGqIOD/J9a4SpWql/DgxU3KbWo3AkN+xMsVJuNPAciAbxEWxC
mEd7f//ENB7WsglgSF2SxYvDksbVPJTnpgMMSrG2im9BaWhgA9xLqxLpFIH5JDUN
XuVMgHhSlNE9Rt9/LwEDE82H+xNe8rmzqsR+zQpQ+bxM5BXPEj0VE5wyNehA1mV4
KcLUbJT7+tDvxCFkLityMTjb0xOh6T6WsFkFJUNjPblcwtByMhwhNRzmc57qdnUj
cbvijJP/nfvcLAtzu8m8jgbrm5DMCrFFxBO01sbhzFFyOIa/Nu0RhbDtrgJTaaFQ
pGr2Piik+4+7+AFlH+B27PoS9YEqfZ+ADtTcEy8RvU9W0Bzrv1QCJzeiN5UO3wBH
YnSWQLOLGw8qSHb/jWRGqRRquCmkAZQiHGgGqgHixiwc3eCZd2RpWY+zovXoZ1R4
EovZMRSS6K43iM36iajvfpAuJUi71fyo+r42AMRhym74ut6rLIiQ+lGehtx3rbwU
/f/ds9zjMYXWeRwTRcq2zT9rULolD4CIdf782evB3/6R5t/8AZ4uMJdAaU3CoX0X
5X4gj7hHecOz50PiVGSZqeVst+eWKOTVlW8+dF11S9NSn3Y7rP7zbmeoRv0QyPm9
ga8yBQEfgtn+veGew2njjLpP0y4cqkYtkkRA7gFj6Ig5fpHr3ly5WL5669o6yYvo
vTR3DPASC1z1iYDep9S6NrdwXIrLgoTe0z49g1e8GC8=
`protect END_PROTECTED

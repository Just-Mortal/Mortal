`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvAvbcpT9iPkhCqXIt750x2pAD///LcJyMYfVwUc12ZmPPiiUEFSx7tBNOYsPTIb
okIk30A3H3qbh5t4s/i/88vbwKAAPoSp9mS2dfX7nFCWf4OECTmdVijnsEVNx1+p
vl4lH9yT2wgPwf4BD1J4eBpiQDfacT1oYb9I2S2T1jcLmQHhBDVpocPIaba1nK77
+k3GVp/9C8CZfgdsrSftl1wH5IfeVPUGDpTUKSpT8hvhBAniIKO2IfY/dRAnxrcq
alBwsO183cqjfgBskM20gfS2qJsc3FpQFTma3OTIkTKuscu+0oVIU5+UEiLTmPy9
iM6YMB3/tPMX6PCoQohgmzragq9+OXyL8hqk8K3RNkHUuOWNQZtFJ9gTaFKqsk1L
YTPxup2NpKpKurRMIJ3Gpv3Pz+ih26O4WhL36MDyPAXlnrUs846j256m4co45aQ1
+4Lm0O2dLjwf+k+IPcHvX8GAX3vpTrKZ7qTFBWqnvsqsQOnzI7njhs2B7QcGbd7j
No09InWFqh+Iar99CXTTvVyMlEK6YfPWF/fCuacwFbkGAobOpB2qi2sanpxyERLV
B5/PFqOyNZRNtkbn06xUcHeevy71BoumK/WlVn5TfgMULXxxUZJxD57knxjf02cz
VenYKuRqKABJcyYf88kS79zPQK7/DUq3a886iWc3GRfUYkOA/tEF/t8CjU+bObbu
7q07be86fONDXbLFIkjS6z6r9IimL0TzOzAdzCbhJdUdnPGnHAcWee1ktvm71wvl
V5NuS1Ws+6QIIegAyqnipA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hgc9DCxRYBYYk9DLB0Varx2CFBLI5A8+Mm8EDJggUaRkUBCxl2x1FgLK7/GTTqiD
sJsTZI8ZwyChWVnXvAYivg2jF9rsVh0lIQv1aAj+kdFQ0PwMqFFRPwcLYcVdLEz8
eJrpKrnps2TBl0q7QKGvI1M7n1lxZKv+b3tMTXdPwjdsZyF1mEDibOkQwWLZlFab
5KCcrSEm8CvcQM6DA+JyYQUhd6w5JDV4ipINACgVqXwyDMW3Rwv0QQqXq9lBV4Si
djfqCwwI8TsN5gY8rO1fm14pvsuJ1tCx2Y0k/MfUg9egf1MWYymrrwqB5Juef7E/
RWW6lMH358DDSrAffT6TITAwk7tFvyEaZY821VXVqs6/lfbIDROxDXhNww28+Wef
30DJ5LqlKSXwnzhKIRk1ANfZxZZ+nb7FTGB0jyHzTqGqMXEl8iBolGkV8T7A9jkm
+ZfgtnA3Fg8EHFKo/RAwkyVMNiimyNkM8G+qiTJnIysV+5fmbJMVU/cIDrdsysr1
ipUU8ObwGa17Hdw72MxUN8O2hTf8/jSB6GefSnxtv03B9xTCem1d/M9obyfquJot
WJqw7sRDGxVpqHqjH0Wdm1k0jCNMRYDLEPEJ0QzCuGh0wlCcVE48voY6PF87nVKf
mx2zcy6Y9qkI9+nB4SXB6cLJy+ofzv/hllmrF2SGi7VC46tiEMTEnENrizO88ROW
u/sTOJGwsEUix01XOMnvE/CT6MPrqym8TjY9wkQlCxZUVoURlq+joNd3RNlO02Xh
HgueJ8ldiM0yyw6cBLf061Lfk9zbT6fvo7wHfBQTF5aQBSDBxYaxK1i1WDQN0RGY
S9QtliXCnunYNXDvnQJywAiMlMmHprcWxZ7EhoWHEozrM92Bb2p23MtYezdzqa1i
oZnOBV8KpexPAeWuKj1g8FJTbH+A1BQsjnCkhfDxnuRtbJCzXUYWpsaFIZEMZWdq
NhV3k2NK8gXtN7QrWxPOM5VPW8plXTLFaTwLcorDwvtieM2NruoKJDvb+nQRaHHp
jVZvV2Z47SyvBwTkXpg3GKGr1obmiWoFEH1SY+xEoeL5TRs/pJNGbxqS1Y1EUWJ0
1FaNzF8o8xqgLrtrkVkkprIzQ7GyZVDunUGhWkxHonbDW6bJT6Edi8RFsUGPVZi6
zTxprDisnz8CCcDUMn5clwZgZjstBvPkS4YwItFPPt9yJJk2F+0JXGih8sIGqKQM
xe9+y151jD2TkhmPXquaIPwS8QCBERyB0Vx7GeBNKPTlZ9OkCB6/aCfF36ZKG1xk
ayxxDQ5UtSFEEmhjpnNXfZDxwHmlX74Z5PUmPlmnwrbwULrnFarX/d1xMSYoP/IS
d+Q5cmXQFSZeIMrVZRHcOo/lqqcVct4ib7l4zicIffB5UmY0EKxHva5P0YaTZJGA
NHPBf4sQQQnM679wTlSsDgnPygDU6zLObbjMzdvjoBiIZ75K4cDiDCAZcnNRXqFP
mK2GEbclVXPUPoizOAJ86O+RI/OuW1HCCrENS9e7K4qUpxlXPF3V4+ZlTULvQZZV
vTv9spC5ZzOOqCBp6QJj2I/KX+5JO0fz0uccJ6g2nV+8bq96flWav4flVg0ms7Rl
l1cA6ogCUuvjL+JfrjSH3zoClMSxNX/Hn61/g+py/D7qbPq22DGWpb/xu8nKw02V
3J2PdMEK5B5Ar64mfX+E0c/su8FIgi82lo5eCQRL43f88+WKof4dYD1fVkxhv16c
UmrC2gvicql9cNJyJzO9J037rOE8qdfVvBch21BBK+2m9F8Gz4XJNE+tIqlMdvjF
3zhC+HX+FeXbQEkwteK9tCPCL8nQ5IsBic4HiXwxslCUWhp0N6ptGfGO1fQjTgix
uplX9GAlCs0PEq/sIaNFiR7hyOJ2zfof5GTJsQvnCfpUfz6/gNwhkRqrxERSv5sF
qSGu1cveCYJxICav3wQbO9nSABq0YDXFcvS/hN+wrkq7NT67b+42bn9zRh3EMIb1
9YOoq1OEQzSydO2fnqfJWxm+M/nHzw5xtWvSbSf9T9y46O8nOJnha3LzirDGJxmj
8aMxVYzfB49JpjPnsdbEvHq0UXL8aCfWDZ3TsRcpaWWeoOrifUu05/QUPtigr2wA
r/qtUJflXPnGSynSgsRimodG5Kmq1t2tCZrhUUmb/oqvyLiqMb5sTSnLSXcj8JOS
liK65OTnqHnSSWdZTOFEvi6gosDAAU5gXS6RUeDUkT4akN+7kHW8NDxFD0G4EzzX
hbyrQhnugH1NFyVMcUu+tOZNcowIWJ48oGwinWAg+y5RPnN/gYcdzfT/YPvwX0qN
kS4H5ljhFf9QtOtTU+UzltAkA0suZwH8DlvFMEiTfOqGDy/Dx1kLzk7f0kkk02fL
n9kXrejwSyxOHT1Mto2Ab3o1Fzt76840eB4aGU3QJX8SbHcfegmYtvSitnwpo276
21F5yUx1qHJnXIKMtlVdrpBeLx+QnRZEow4qQ5qCrVNlCl8apsz6Z5qeW1MRzPjk
0rlDwu9o/ZuajWRed4nirnME+jIuo3ObsoXi399ro0ik9v5EbWDP9P4C4u/WnhYV
27XLl/3Cnk3roFow9VxkjQABbj/MGQsX6O1Cr6c7M2yS0Z50JszIACBJXdcsGuVX
pJnJ4QGwfoRGuj2grPzFJECidENbMpxTo1G06SP1wpnim0k0DP9wEu+ww53ZnC15
oF0+5e1uEPWFitz1L5ZRRHiuRKckSF6+pf5HLDTyY552Tfm2VX7ftxl/ROpaoCMX
P63XY0OvI761uX7sG2GGFl0B6+p+XJYnu92KeZJXkwObCdhibfNDspa7DBC60EKX
UkfQCcpc5xTFP1etNUoVUQAlbiEKt+d3XF5rEarPa+cltIUL5rZhBSvNuRhUyeeG
HPEnBjUi3OwMORL/KQtaFqKyIDJQNKyzP4/Oh/vv6w1reVdHeVcCRL3y4OKhnySF
EPWGqtbUrJcB8E0fjUyPXggxxYR0CUUmrhj6f/K69TvOdPBB0yiuJXNZcQlHG0xN
wWR/x7Hnh3rYUDCywZV6WpvmEFwH4nY5vDbmjdCdM80CjFO4kRtpNc0P2wBdyZ7k
hJ9KY0DdEDBe97gdA/vEykfcb/yaf1mQERALJT6/eOIu7LrNpMyEFtcBvWZqBEix
pfKc3meZtErWD1W4C0GxJY+awVmono+0vSMUtSOp1STJCOTlQaidv8CAoWwYoitH
82S2kuJdVNwTqZiDORWUrLKGrMYpA/RO26kTsMZHXbebXAFMAqF9PQEJUw1adn28
NKD62vVkkjbcp3CqG7vGV1keBb6WzG2GRVpigFgDmFmTIb1ShHaEw8mLdXHziSiw
bBU1P5wpRcZtwzB6ABBjwuhnVgEkY6YVH6leT9uJLi0lCMGKLh/9lzwB8QuxbW/D
InKTf7Miey2GfhyCAgdC8yAuC0XOAyleLQnePqZSplxaXeUk4X1qv4z9IfF7zA0t
l7Yg9mSQNab39xn6qXcxE6n9C8C30CBejBPchRYEyeUJFchLIP7mVK7/lrUaxHYd
QiRB+EGdukNPPs81dmqBzfpAnRn2eXv5ZVK/C2TDRnsFHXEvve6YmLKZQfFtU0C5
B0shvM3FKGDajk41HMsKEU4spaJ+tI7QkvpyiFW3caJ4vjl8ZRwAvZkdkGj2YWEy
Ty0cJWMPAyrnz0Xv+trhz+XVfbreaO7xZzQ86H3P5kwu/l8WR1XBkwETxNq8akZd
OWeB4MOXpnzkS8yH7VGbnAXnvEEsmcZlvV+Dmkkt8qwHe1ZZWS5H2KtyUiEIp/r2
ykdKUqCO8m6OUWlaYSzzXdYZgTk6IOaEQh1BbTEWMQRpUIdXTpWFPaYv+Ws01hYz
b/thpe92L9KiwHT+RbZ7Zl5N9zWRrUkAFD8eDY4CpMfm1ipj+1SexUL1fTMz1T7r
FWaJFIH0uGPc8MHfo46qIXoMqvc+x9NCtJqB4yrVyDc5x2+wj5+yy4yZXmxJiEVy
drnZRsH/JWnsWxzNmEcBYuzY4rimnbhEkVaGOlOvI2ne/MQuPtJmDaQm3EXu0Aa9
wPIogU1lD3dTnzzSnAkJvkfECITpn9p3SlRUqXbxw7WP9FtmZXsUWcym88kS67V3
XbwpJECS/mw7LX7uCoeDZ6K4N8yf1j6EcJKrBhlBKiIYEID7AZAdk1tyUuuxMpSE
TLG0/HIy+GtBgYzITE45kmUUJO2yssXnbtE6lIb2TVm7hutwbE/6gDC87PQPLqWE
mBM0dsOxQ7fS9Oabw5oOUyBoZMeXbpyhNo1MqFruYAptiFipMHHfss/he7vUvGNJ
07zcFwI657vcLX/IHfz5+CQXig/RE/xsBvT2cI8tjBz69xBxo+R3UnhYbZs89xOC
1uflzZdgFBTb9NiAMEmkyqG7FHsnFKzCtlnMsZxj4tC8jEHUaPfsLF/cjkzOY0qZ
iWW40QRI5YJyo7u9Xvbyb+6TkL08c0p5TXNGCgKbsl4WiSNjmI/0M84zYyap06Sh
iKwuT1kg3/+BY1VG6JKdmWU+yErLnVcpK6hZEL6XU8iemfdlsgzdCfEtRdHb6+og
pM3Sc7aGlxJ+ldVldtIiqApMSiGgHKJXNSUOZZVSqk1nc48wZL9l5wbOSvz76hf+
0dHM5G1HL0/Aza5wLa4eRUpJFe+miy5OoNxc/72e+DzZFswdOFHvqNi132X1EkHE
u7PiSofy9wQ+0J22JnadNQxvNoXMzx3TBmNYh/+1vCKsJn61+xU6GPyWW6YemEjX
HApxsSUYaso/hUadFzCtplEbYmfMYfZehp9s4fFr+LcVct6A5W9/g1FfoHpykCGf
4EiQF0lTLf95E/kUdHP9UTQ/sMgBuF+v51x0Toq1WcahuLwcUNPQyJUEyGR6MjSC
SemUxs4c2uhSgY8LL8rv8L6eXcKNM3iLTpqQGo7sHoxhqJsNbqoXNZaRjSnkiVwo
XSkY1Quq7iKWAARbXmIwUklGDaRz2IklC/rR8cdXlVuFcbGluZG3Kbdq8cY1leUq
Yz3BUl4O+Py1kHMSTtAH0YmIzDz0AvyLa0CC8cOZbruKye2wrJW9OAoItK+zI7+i
Jrh+7QARRRWDYgLxlqk5JBs4A2aSKvp7HQ8hm0EuGpSXVApjmKwiHYZfbl6aLWYC
ugNddEsCotB7B8MFtFWmy/3j+eG4WAh7Sh6rIKij52bzWggUaq/l7GlG+EILdj8D
OaEkxY5Q33t9l+dsnx2fL0zi8aB1J4uQqJCMlMvt8xAINSxVD6G6QjMUkaiKspkk
LAIFux33gynmgKkHgMSQePfpJcqY0iAeJ2rnReJMJq240hKSurtXx/YbfNnD3Y5b
Djjr3H52XKsr2zf0kvu0+zCnCo1dg7G6a6TIT8jX0y/I+QO0uZujDqFSR3lDjay5
Lrtnfo+6j0EQoPf1bGufpQwysbLOHjS1VivALGBirvSPH31eAdpsXIXuSb3/iUsc
sEwSEt3C6xrOd7B2nPMb91xNhegVZmzBMZ0rSUPhsbZf9CFjX5FpZqxa3+qXcznf
8WSd0+Rz2shvCAx389E+C38s3l0n3aQcXajbvLIzV5fF2w1XPoPJCuL9+1A6A9xN
KF3fu5yXc3bPwEvNaE3CSVfAhjXe17TUrL3p2m77s6v406Qzj4m+rqVEbjVZAnAD
Ez5fYfgFWbA9fcI62WlZqcKJD3q6ki9erL3vQW4EJ2AngkEPEJaCT0POPbGeWL/4
tsj55Kjs4oNUVdKPtK4+ySPTB8L75wLSN24G1qC5Pv7HHcAk2a5QJ5VHSJ6qcbb4
yMkodRXpc0c3a/oTOckcjCzboXzSnrFoL6FWWTdpll6zt30q259qTvXeAEkttLYh
zRuNB1LW4tTp/N/lcdwWWdGkfbpZJAmMYfe2LpRuCs/oQr20kawvFnOr4QLnrv+i
8CtzAAHlfTz191S7JKszlK/M0d2EItSWQkO6aNw6RQkc2FYooAZdEj13CtAF7bzz
FXBAeLONvssf01bN25/FbBpc4YtAxuGwWqDqKo9iGkB9a9YACpty9ykftAv1Pd8z
eeN8nH+GoLvbu5UyrzwNQ9mw2MjliXx71iFxwdT+9V2S2jFb37PUnfIW+MNXIdqx
fytAFCXvDao5K7emsPyX2qhaOJBeWMH41ULhTtdRaL+zSzGEokkN62uZK08i6sWO
n7RnystUt55uiNWPZGW5FWtId0EUibMt65920fmWV4wsr1hg8k0qWTUm58HJPaex
HtP36vzSF1w0Ep5oGB0SU/76WVpYwmGKtywDFDAenXxiLRKEXvPzq2DZVmS9eDGq
8xsT6BRJphSDgqUCNZM4a94Y5RBJgTCNi0Tx/WFvgla/D5VnqkD3fq23c3c8arNo
fzRBOFiaT5+AFlc/M7LE5DQmQxy4dDwfKnTutC1P4lYlxSRyKFslBGhbnLLLash8
yVyb8Ke8KW+gxUQCoRro5WLtP3/UhVnp5iJKNUz0oDtDjF4PdSTg3UbqYMSHQV1c
2Y7ia8/r6Qj/LhY/Y/V4d4lHxVpKAI79p8EC985k96Bu73EE7yrVm5Kezk0Gxh3v
BaJqj57l5UFxhlC9EMqn6/gsXAFGO8nMMT5fwOlzk8zjYblz+GpPlYeoZDDpOyoS
nYTrJWfRX1xi1D1WN16NQJRR0TYnI6mzSjePLSWcimKttjKV8Ig+/O15Ywmmk2B6
tUKFby4Ex3ov3HIXHdWUiMPU2bKusMrd3EYqOhfOUfJJ0TQ7VytrHNyJd0N3m9Pw
4muh2CVUu8pijwqSHLUPObuRjx3KNjx4fxqt7fLZDCryF73AWgG45Y8glT9p0Nxh
6ub9U8lUoftokBwl+k2Oz/LSA/x4Jt/2TX3pgptQKohKs00fTZnAw8wlrjtTPoe8
X0F/GHfoi3agU6+xfU2Mhv6Zzuy7R7WOJ+n1AQePs+oquUvRZ76dkIfpDygSaHUt
mHyZ1LIW4fNJwi2i8BaJiD1ee6iFgt7rjVes5F5oYPoSGh4YH/mRPBcN4oY8nlsQ
pde1QBkoPNdgf2iXcr7XYey9NTJkCtKKF9pveLwjeMqFab/xIJjJrSZea+ymeZwh
fgU+hKF64Tt/u2gr8ijU9hTumfHkCHU6ezuqqtDv0riTO+aYxz5NsqnQ+p6pq8Vf
SHvI/zcz7QMqhqiOKKySFblqfytH2QYRCpe3qTNxTI+R0828E6xZKpixKA3Vqj+q
hmZspyXDhR2hpHFkNtuLagsntDZAcGJc24XU6C38wGj5nMUooHkT0puCcyBdkgXs
XoVFWbl09yAq2sHD5p+0m+H/SKHoPh6e1OFfkS7CkH/PZPH74qjnRitzOxk4AfWr
1Ml/x6OB3a0aVxcLlg6mHHUMhwjYVtg/wZsorPpAShQe0IBmifH1Yw/7iOaop03i
zKeqFdnupwoV53XwpPPB+eelIcNe5xQM1b/0XZrq3XHrm+QMGGrU+L+QJMbd2cNL
4tsVwe0ZANklHjmfPUkNN+4ZJLOelmyFXKwk6k29cUbJtdIs95eQXlQV+ilSX/2F
7zqWR8rc95HYdnScE4sb3EnVynl0fBsdJ8rKi0ZEPHEC5Ixox9LnU0/B9mo6/4vl
6r0cdHI++U4HL7mAQxiNJT33CtRHXL58BnivsNWWPq+JGaC+VcK9zqnOtPObqLl7
DlgftY7ybfxBn7YyI+ee9U+Q1NrE51XtMluCFam6jQhAJeD07KTCfcZEG8L2Q9ka
Lo+lW0/ovhScKv0Sl2uOnnR2U96s/+vRQSKFBysSJPfx4YxdGvBQeZ2PbVqcjCoF
SIjFwH4yUbLgIOIfQMjbbQsy5M6p/3WYHyyMP33DTIdZrME7d9X7ptKUJO1MI6oL
0EumsDgMaWI6P7mzv31B02ddimsgJ7sDtGwWbBPhPKWNJpHuoFbQ3hbcFJY30PDU
f1P9OwkeIp+b8I5gZmD3mj5ylQwWgfbYuEygkkxI0YTJFhJWE6PTgGIkrYzBcgNT
XW7bAbS36eQFA32XwB45uhb4HYqoejBhcPX4GvA0Pd9MQwlv35OYHtSLDJSOSFv/
0aBGSNEbAbIthTA8mHToeqtWiJZMttJ7KPcdDI4u3oBfkcXVPvoKMxvJ7qqy/5ii
INGPvFrnDlRFt7TRBUWJd5KeXCySdFz1cY6ENnfC7XSqmJBK4E7ExsfddIkRRxHO
8loMzHZcaz6EF8OIRmZ4wbFvfJzN55U+DzHgiTePokluFlaRZPoawJOw8HHiyHcE
mtEoXpGWMUdWozNA8LeCJU7umrgnvRwjTsEh5PsaaUnkTnEeeYUp9dUDqDinycxd
LSxodU+5wOEjiHJosCku5WTm/bdLBTBRT4UDnXIniGZH+rdxYxFU1bpYLsBWH7cy
hN1ojVOjWVlWm3pX6+LeEpS78p5pQUXngknI1ZbRYfDodPYru5/rAmW2NMRiLnDA
w5mavIcI6M9VqRkW0xIWy7KcHTVnf/0y0Nn9hQsySdHGauEmLIAjNY2eyjA6iJJa
MiRpGdbFP1AVS4dZJUVOUYEKDvkYn5i+t1u6j/OrYByi87GT/n2P+yDV611oIxf5
URD1uhxZKD3eA5q3x2WbJ7lAmYiWMAD/2/ICvTK+lVe6X8kV7/y3+TQasF8DXSie
muUSv0HtepHvs8stpc021Q==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lREh36EMXVoj5ihlYzvafrPoPIUQ04Uf9zu5NkXzMCDbln6yLp7w+DCSHDavJstI
6/dWhOM6m1lihrMp+dRPTXM3zBOsACqmYRwAIabqbccAU8rvgVXDMcDwW0potRrh
9mX3hwdf0Ti7e43GMuA0zBikQ4rhM/z61toLF1lpBLdD1S8rQDvziBUQ1SOIOvKG
9o7LZWxpJtqgu3CsyMTL/gg9l6kVddj8lcS6jPAS7dVb5qICCuDYoIpZTyq8iXOA
vo+ST55Kjsi5dgt2FV6OBjrHMR71GpoCRcKvAACEzUcW77k2uDpdMElmrf0NmU/0
4j4azcMNmS4XtVnCeEwO0XYbzHCHb7a4bidA7fGjOl3ePAl1bHPdingAwemvJthz
bcSO/AFFyokF3FVk24PrSWAA4Uo9OWU4roAU/NIOANiGtmzTlT3TDT1+7gB/dWB4
+Ygvkcil9WPEzJ70FqUOnRSFJmJi086vB/IFRSBdM78ZRtq7zVk3Sf1+uy8CCAHM
EPRvI9bDFJe2ECFy7yzCUnmE1xVoxv5Q1x30wozUxQvNBno4qpfv6jGAQRvmkdEq
PTMjijFclfoNk+FiCoOeI8Mc/9zH9A9MF3Hqt4prHzWMVlyhPqjsJ0keO5cl6lsK
6NbvIBOToE/Y0Ep8MS9I8FsLvuECXi656niPbs6pU4V8SiN4ITjqIhCK2euEZTYb
RJ/k5HqAsz7GXfcSs79CpBwsZ4Ki3tO05hcYOw4D9rRrq3eYqDgCFRJBBMPzjOkY
KzgihFJzpKuwaMiOC9GiKkP6qN51u5Zl3Qo74pB+o9mYKG6Hu73xRoWmEnouw2M7
nPw8iRuLadXEI3Cbrl3nJWTUadqFY88Qd6il3VSHRgkAq50i0oEtkcVtCLtLz6qA
FQSgZ6HfMQGbz/KC+a1mSoQl1bUG5YiF3xjW9eVLSGNpOXMUu0Ze934yf1G1l2ZL
lvjIS2z2oT3NWoN39s8WWsOoNmCcrRkWAZI+5h8OfiESyCu10LzfWwH7DULfY2f8
7qgXjMh8dzN1NZGYarWjPmX9GT9uAJFGHGFscmVOonkaTPqrNePEwq4CUDesOcld
CPNK1JymAyBsw3GKBLq6j5lfrfXWZeA+IJEBt54CcpzIbeF6DSG2cA/lWBgVFkko
4ltP9FuvAdhA6TZBJI/APOd4syF30K4hXr2f8KLO3h2opNbZ88HdOczBUjKSL2jT
z8I1VMYh1ZdK/hM1Y6hW3mjwPhQktOU4+JXNu590+z2Tq2z3HzPexjEc3kCCWUi+
zhzwADZJLoOvTDnZg2axCBtbpB9kt5VL2+B3qwlBLI7o2SBTmr+AkkuB94wK2S0a
VzRryuxNpCMEBHFaY+2XL1YkjkL/a4WpkZX94NG/m4Q4iH+CwBczwt4TahlwbjDr
Wk0H5/AF4rQrZZwMKkmHWltTbdDoaw61fdFvmKPp5expcdy5Ia1h8vDEetpg7Uyb
v76eod9oDK9fQOeWQq/uZXvEyFbEhT/PFneTJ79QKEyPtzHkSLx+DzTfYYtDBis5
khacXxBuh+LOzyMfeK4K9Qj/zPQJrvFXEUQybc38+NcynVUiY+MYQxA5+jUDoTba
wzwZX5kJ0U/ZQeLJN9CBXJb6ze9mKSdPeGeocBFvlXkIgEaYmasSZ0fozV+WVxmg
My4zGlsoWgZn4MEEBbqt0GrRvlKWKF+rowOHZBp8Znx8lBnt3XVT81TiJoN/q4fx
G+wczg6nnsm7ruwwejM4Q1IzPL+HymvPX/FGblRcf/areTZeK5osuZQfrHoQu5Pd
Jp25sTy33chpciR75CFTaHdv+HRASN5ll6WvtOba5SRtUqNeAkh/21qO7BuRupbr
s5f6tKCmTdCVXC+Hv/Q8sXuaTnjXAKkLX6n+BGWU3kJZmdRmRMj6U/uOQm4O0r2z
ZYdbiul2g215WiL5C3vK0FArFSoM8a6mk5jGnREiXklZoqG+owE1YXstl4zt1bhv
kd/gkS81rDf999u51FKonMVvNGPGuIsPZvMJpiOFLwwOtzx/5VTRe39DMX9+7qlq
Vk4IHAksp1Lh2iPrVKCZpEORY/qNp/uayXZgg5CU9/awrkpU0GZXPd8kgrNRS09v
PTmApvlO7VBWKRpeE36wtfimp601jCl8LkhLLLQjJrwuVH7efITuoPhfhiqIqu03
WH7Fpt0tDk563g7d1P25QtEurRoqTjFEB/i1SWTkM5WZ+FcPpVYxMm3pqpin4uAR
5X9h18rQmME2TiKT3dEw9o8IFHj116dt+10iNSOU/J92BHDuFcNPdCElL4VutqKl
ENWMWsYR42ATdvr/ZmucGMEREooloMYRQ0q4LdJUdapVViJJsbjGV4bvcJIxi4Y1
Fk1daVBdaLNXqSx7tIWCTeylHndwu2O/Mc9onNnZWuh3qtZ4lAPbw8TTCBMUkvBD
VQ8fHV6hU0jwOETOKhbzeBrGbIylMwAg9SFYvhrdIUXkRO/dcB6WN8VM3jMYa+d5
U9cN0o7SZ0tXqDbGSmasPmUfszyJj0gKYsmaxJsge6S7JDYhxY4I9XpgYK9EaNcm
bcAONQOrgABf56sBu+ydzkDqzxgaCyCallE9N5VdMVTKb6q9aaFOOPld3NtupD3l
z+x34uC2/GiL2YC2/pJl7z+0dB3liTVVi9o/rplW4EU6+urczmzCWZnuwO0QrMig
jzGbISI8j3wOoepUnBRoXiaD0FMnqBSPUTY+/0hrRIYy1hJ4nec7flFwUxE4F5eF
1Q2SMvpLCtIrIEmUZG2B4/rC3KjeHETGveULZ/2phdOFDSfFRocs08rFgmpDvxrj
rBBJXTM14uHugOc7j8lKWyI9vhE9GFM8ST69vACk8wq5kEuKDCHCBHcaY+8n1+0D
kwCrJa07hK40QfB/9yWAattrWbPuSHg34eNe6XgxrvDLliMjB7+lvUVkZ3+O7SQZ
a3fWKiINdGmiQRa8VH0QvpVKC43vLr33XAqHond2iHWp45VlGr6498TPHPOaMvud
enRf/Agty0j6L9rHfzhqtsKsf+9NVg00Gcyhw++JF4tq+kBN6xfCC3kFAj2Y0GOM
bNEPfp8hydk7wVWb2hYoI64yB5kWFiLysyIa6i4mJsJARoHaDfEdhRCfI2C7/pj9
VhZl6Z2BOaj+HXDlxMabGv4/CK8p4Mf2sesbWjr/oYf27B3LWZeud6GluvOCw1GO
KB3C0rgOAR0LfZ1Jb8JJmrbIMqdGE0WQ5yVAPwSbGNtI7p89lchwOvug9xyEZebI
LDN+uh+m/z9mFrhjfYsla+k7TlJKsr8r7qfEe3PlQqumvqoGIz6QcVZIhB9TLAVs
FMsm/8VzzIctObjTJYKDGc01fRiQHrb03+mwfo941W02ZRJwWI2I+w69wZ22EbjX
vzo5IlGtrznT0vroCirhVbUsckiQFnzy/+0wDEb+4XkepzIv6vWeEqkKRJz77FY0
+God2cjpdWXF3SIcTqyQ2cYq1yOScNJXClh6pj391b/eAunmqu+Rg5WW1bZPm+CP
rgTOchXa00O9oOLoxoYK5vARa53rKflUPmOh917POiq/Qf/sKWZ9kVvoyVksvX5z
NPc1L9Vw11JpzyEsOowJ7bs1DNotLC2Ro/CB5Lg0NDPvD/AxAqqRJi2c4PxdHdbq
trV2xteNaw5cHNgUQsHD0/GqMBJdqONmiDKZhensk075BhJtqxR44RkbWeqdcP2L
EkdhYG8qvoZIZIMYLUUFeQ7eeh41MU0G+xICG/r6ft+mFPUrHvHFF5vdJSLSv8AI
NQoXIkljtkpRngFHaQGiekNZkYKEGvfE0ntN4RND8oMqu4dOTgyE3Z5B3Fof9SWC
BuSb7xfFyAIkpMKWbw3nb9uGeYyITEtAZz+T158j34cyVuC7SmostKjrzRbv9Hjg
CTla5JDT5sVxcZZb+dZvF02l4OKvHgRPPrXXaQDaxlwrJVdnv+2b3Vfq5wSagdYZ
YAs23YFKPP8DXenJAKqM8DVvaX+4MEL6SVq+LjCzHB7w2IMuLKhSMu+ChT0gxxCm
vi/E2NKqwO9MyV7L8aAcM3bzWOdHvIG3V7y6DQvMXMriNkstdN/qKLWbPf5BCzyG
s9dmE8CwIltqZN7mN6oYje3yKAEB4J0LGFO41Nl0WfBpQICwoGLVvaMh1gE+auBg
WY8G0Wd1aJgNwK7nWZ7rgk+qe/KNGD9bNmVMIfojyFMmh4DO3mHIcG/M4jpJxgGd
tseAs9/Rtd8NNX59UUQ2kn7OX/ydfw409w0dolcFjrM5y2SQQcpLH9a1jOMB6pVL
OxpW/pt7C8DmafJkOshbwydBl7vJypa0wLbcSzxcl1Za9NqoZuAVg9kBpwCkpyzi
vw+qnlgbt0Xcz1JiUUm6MWT6eGsVtjJ4QcnbSO7IyXv8PmIs1j8Hc52Qx4RL9T6T
nrKcoXb5UkTwvauTewz8A8ZeFTwedqJ79v9Du8aU2x2Snyyu+aNoTOBQmjxlVYjM
bEgFe14/e2HJ9gFiu7MBV9kigIBkgsOsnlurmxJdx9v0IC1reBQAJVsKGFQHBbSt
ccKS2VtHpfylqMNwXqdwLS0XBwRQJHUJo+t0Nerwo9EPPZp33OQEbk42XfLXlwox
flkIXLNt+NOa/PgSJ9fSAwmgZEVL5QfY1VdgJlm/Gdgy6FRog3R0n3YDawmPjcla
P3L+N/Xk/dPKIkJRn9loAqiKP86KA/7b28HQWpIqI25//AMEd9rn12slVCFMsXIg
GbwbM/rf3RhUzypMDamDj7OPHY+t5PeAJSdtIFBdONqa8JbyTZ9s+X99KpzsiLjh
mihG9osX3vq9IfpH1F4qHA4YnXuFCR3vc0lMluqPel0uoNrRMpYhN66OT8lvCde3
LSG14KEjnDjvRBxqnmXNCKweU9HXfJK+MN+rvYPf48t/MpN84mQHTSeyYHqu9EnZ
MeiH5CKJJ+rxktKiaH1o7eHKIgfD3YpeY3vbxdWtQshPb5d8dIzLOxy6EfIvFY70
wRM2qrUbKGz2G1QCyOa2bOxaRKYqOIZ65dd6IwA9xbFNfxR0aaRF3/q2rBTu56c4
J/WZ/xFTcbm9yMJd7NRMpt8l6eR179nsuE/Yd9OlyxWW+lLoXkkTn83Uej/YCVMt
+Yl+n3yQejQT8ytHTBpYxLW4S0tJTCDe2pcL3OaYvYHIAXKeTNtsbROakEPf6mzl
BrZaNHLLX4DDjvSmiB7O99m49Era3XngPusYZRPLC6NEUbpoJPSHIwI4myHcKa7i
VsKWsF85fiCWjUsnkJFvUHwyiCFr3CyCMbaqTD4+vGg3GpNnWzHORt1oi78TiFdU
ZCkQ4LAkVvl/UpB2iCq2rBdf8PI4AYJitKYQfJ86bettaeN6LQX/OkN/uevvCAgb
DfUIZL8JOIZGR7FpsfIVkk32CLXa32khGfVjHax8iqL00hxKgWAmxbznR2oOlTny
hFBEHDvROES/8l7uLknURAaFxV7UbkRm5iSrxyxR4ZMrZYhSWLmq1RtkePyWDdQH
cxO+6B4mqPx7EPbMVzGebxjKYEA1IlDLUHk7OHBEYd/XqRrp5O7IB93rOcb9uNTk
KRNMIvwbmAokN85f1HbBYdChcs82q4/f8Iu6TT9JEEmUvxL1OTnCTJcxIv/LRTzy
ULUKCMRKYQBnzMYac5XJLmtrFrSymabPzJnosrR8EGDUFLuPeIpXI7VKdxXpPxS3
+ot5EBrULfJNC2ak3IhSn9dPOi8RGWSuoGhfmICQqEcl8Taqa7lRNcyR6CmxBffo
M7unDOES1HQSvV8K4yXVNiYgPHXmY1YDLZhLfSKm1YzCWx3Ul6MT0hnapJQPEctL
EOOm5OtdTNm5ab+1QNbmJmCv47bgwQugLmA/h4sneytBkkKPGrStt6dX3H0r1Dxg
iB/BUv9goyHhgVN9gZNJ3pPH0Uruqh1/MLc2uGIzeLC3O2vJ+P+CHQVkgIbobmr9
IZtiuZCq7t4ashZD3LJpeiQr/zQd5TozNOqeYUlrKw8lCQLbOf7r3VMGARWNwVrv
xd/bamN3jJfJBRRTL4FJh2T49w4D3qYcENK1P+aF0NG+izXRfNLSF90eqvUK74KV
0ywlC35uvJXEXcFxUucr0O8D5vC9pyyy3/EwR48m2CfArjqmyBQy53I2S+st5KNs
8h3VqmUhjz+jb78v9e+nU1R9Au9jYQrdddVJEXIZ7jJ7vK5CJmmXvE7afqQiiUBV
aoGOViIaIGhTlNHLpWAa6kn8p3WLRlQPEZLaSvoQpRLkYsjSaHsQiNdNGQ1pGv6/
XLUXufSoMh1jKRkwKQUMnBGF+eH7la9Q8Nz7vFuiI8sG76dJ1QB7lBm0VOWnJr+x
d/C3yIjgVjqpi2YniNTabcWG4qd+gnvUQdot1rEr+1VEl3WzytJF7DEXCtRnx+Rx
8eN0HMQCFyq0viKFQZraZbetgtyidQu+B13Kq9tV8Uqo0QX36Et63KIlsnZXnodo
WF3Gm0extl4K429EY6vOxh9L/SNwdciEQBUwkCXkvn/rr4hypvOwe62JMTUNu29O
P+V0ms9NIMgf+S2lm73jycxc+/akL+SNv3j9+NPkB0Iv5RQKDFgeOw8WwcgkKRfK
HK7X8hQL90F77mf896eYRb+iISL3jX9xPbT6y/d365p0SP/NR84gAkgzSI8iSaQV
Mifb7l+2dfwhHBPuSCOJl3ECTimQr70/vm3NNhQRxi0PSQ/6OyMiEsHKIfoha2FZ
vGIuHm6poTF3WRIMX3c8HMBCjqM1QEyYkxl40/EZq6XIHoeZPz0i8blEvnPsGanI
JwZwMiS36oR7WATAZcRzNUM1h/Uqh4ZVWL/HkFkGrCdCiaw+amfwLxVgUQMnU9bS
xNOlbFmi5eN0E9sQLVI+Eqddc+MHCfWbeiACF5EW9iCtwAnjm0u475hw6BTJoqrL
AgYppvQbBHxuZSryk8Gp0jYrgzdTO5yCtdYZFx5ZPoSLjhW9D0zkCJX6BpQf2ZGf
z4TTFCanuVVODsrDkP7EKRuoV+CxjL5AjMCt6NVEScBBELog88g3oPwLucYVD8KZ
ivX11yWrVumIXvQ6UHYDLyUm7ulVrn+pdmkN7U9wywrLLkesGGUFl380n2p8WFO6
oZpu0R7F+oV02PeSH2r3WN0R24Hi/c794DeSta8+WVnDY7ib1JQddAoLTZfHWMND
7b5ValODtIQgO/uR+B13aN2L5GF04tkieR50OEmij/4GfXNUuQwk84upYokvYZdc
hc5weLAdWxlvbKapqDCnKxg7X9x0BBtVqKf8o/ekKX/4KRxSZUZzhn47dzT8ecQQ
WSIvP/WELREioRSP3uXyGbC9hE8YJBUABMh9U+zaWwYLa90iq4EhY82XOTVOxeWP
Y01jofA3rYU5tpO5mY5HYH7ZK0XIWtsPvsvgDGz3hHnWLNxwvphNd+xPvAd9sajs
26gmugIo+W4bH3ZCo9uDDkrvVbj2e4AahPATENWxgwsen/HUnHjdV82v/k4PpxP9
l3XhZyuqhkDhYVtldUHwqhhQhg4hNOD0DR/e3rX4LJNA7vBg9YF4Cria4erCsEAJ
LoUsAWOrr5y3BcbmeAplnjn5h11EYvuN5gm/cXpT2uv/GjI2q1E8PFdcqHoEtLtX
ikYnE9rWGWJE9dthoQDPnAUIajjal7BlSArf/SRcBD4p/ESk9VNtHjZ6MPOovgfC
JygKApiLLeJsQOClFYmaVjUt0RwzkV/ecJWBg2oheS7FVQit/eNgd+9/f3/RIVWH
EtkkT6WbyI7nMZtsRlYBJiP5e5RsbUONn/s1h5Jwf9hYW1zrdwRioKchjH3pRSv6
DUDX84dTqWv/7oF7FkPSIH0p6ta5r82nIP87ZqI3Fz+QgvQzK3EvHK4d72YyCNel
ztYMUAA5nY8Xv1oz6g/1GKNhBHTOBWXjeNvMzzbT3ze1FYFHTSuxddYeO+9fHULE
+JdVTNgQp9Eif5F46g8bMik7/cku95ZDJ2y2+tJh25YkwD8X7vayuAm8Tz2rGkm/
6j7arWBcS0P3TYgenY9+e6vcMWVjJrecvs6NyoS9qOM+qI0bmxO4AavwtZBK4tOs
vq8tL5MChfqljlHcJZrEMY0LnHjcGpRh1HXORCxQDA45p8AkJw4cTqjxJhdWxIgd
`protect END_PROTECTED

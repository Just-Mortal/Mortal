`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pnSJMm8ZZSKlmoKaynaXWfgWrU6SoVw8RVRx3/mJpKVmtek8p9UWsVze+Qz73IOh
9D1hYXwVuC5hELrTVAg4GH07Ewe0hLHiokTAXcvOzKyOR+gRLyLQndCNqyK/0dQw
akKojWhQdlew3b89tSKc6VtdgEnNtMdvahdyVtFkG+BmgRU9gcbbQKb/XqyDA+tk
h/cPh8Cj0mZcfDoJWreHNHgz78w1qEPqSoKmKznW6EiOg6g6b5lzzsy6EYVnTde+
bbs3pxy9bm36o9c5zJpWmjE4QAxp04i+PcfQ/Jaya0MNloj4ESs15lv5mLZka80J
Wm8C8tKJbPIKsanzeIKR+mjWvXhWgT7jCAPlcrwfj7hr9tNwZKMwtgNqzF/imgeM
Ae4vidyv/09K1IhH4Zi1HWY6uFwCqkmY7+2uHyX3vbJJM4qaMrFVbA+bVJ6V9NcR
5qHguIPwALWmL1IhFUpb+rE1TWoFIqEMfWEzvXr10hN2e0a5SWmi/sGhrE/RkLMj
ExAToaMOEAwVG0FN8GLqg8WXxRVP8Q1mQpKJDGMDfgle0kBXGlhkbgoQXwNk9CK/
ZrqXHiWuUY6rT6Dz4HGQbW/C1lk4RnkE5S2qj1OLLQupB/SoQRtwVAOi4FsGcM1G
BOLzH66RLdRhd0eqcE/iDM0nADD2R8TxeN+gMaEurks1Hjg8gmTxI95KGuc7/b2e
kOMdMgKeed6UeG4GS+7XNl7tZ4+YC0Bs/3pj1BrqAWo/XRreVtu1pq9bIoQG3btV
8GYsXT5rz/aAoJQ6nXzWPF6OcTpK0TvVum15/wsARlYQkZ7+jA2Ukrg8DbT2S4gJ
562mySwHVkxvWnQwiKlkUcC0n0Zt9oaYbj/g295xLwdMAwFTilPXPBl/Vmrcs8rJ
49xBmkVddgvX/SyR58DAJmjmwk7Y/K23paI3HAGzsR1Z0Ms1xj1zH1//C9qX7Kv9
ezPylzyf/LDiryAY8T0Z/J4UhVFZCuoXg3SVa7PGBr/o78S7lRDZaRc5WvR5GoeN
A6L+GoE47xhB+HlzSeq4DCe39dS+I3Cfea+pPAAFxbwLgLP0x8kjhUZEWWBjcd79
3Eu0zVAKK/pcd1PaVM52h8OATb+dIjR3HgK4wu1biRcRUuRXaxx5Nl5UvbeBK4ft
QQ/AsXplCncIcFBjChia7YISNx4sL/Gs1yvFz/R2QMiV/tKfyy/RNd99HsY7Z8t+
J3nYVWw/FHjNATCzxhbX6jJUcqM5Tsqd0Te/aVdqto0H1IZK2owbG/FAuTXR+AaF
bLiDwmySTNRZYmMkmp/8Ti/6XmYFWNUzkxoBduFutoXVJLCppFHeXNINUV/w2m5b
i8xRHpmV/SKO61Pix2fYu8f+ktEp1GoxE5jr3L4O72/pJyTNsOOrghI/en8E3bkN
wFIJwJ6hGdwHWvLnHB07ASlTTNaKpDIWCbJTfGS+poqe6TaP65DqWggucLTe2AiY
q9/kpDJu6Z415nbGxFs6fIJJdwzi4dVlba7nAI+AAk9M6EtpxfEKOoBmxFe4CTW4
YCgUdORC8R8j+HcDBnC82hEw1MEF8xliDPvEacKirZGdw8LNhYLJLp73lHCf0AJ5
tRw0jSGWhdBIChI+7QP5NrwpPj3ho8m63JbIpn9kxVQFhYLB8nsrFuEcKFMSYX0B
+7RTMrxEea5BnVKpeiQf+exsp3IRYNSACa5hh5Z60Z5/itEQntqpbUVsWmrxCYuy
k7zglVxs7rtZcEZdfCNcPr/zDK0U54WE0/0/fzVAB/k0iSokFCbankRPU4meRy5K
0LqxcY5MGiAAYgy1HNbm9VUtOFyLAntZ7IWg2r11yXgEHCA0A67Lx1GhObncRMpo
3Z/E9OvpS4kqcYpEgbKnbM/BVPVzlAhpQabw7G/3d/8LKwmizoMZZDhrRWjedtlK
OmL2QKq2C0YkfLqRE/Xng87NjJhgcrPU72XYit7fTRB98Su7zdmh6juoamxgb+q7
idjA5Fi4VQFtSXadgnUtg6PKGEHvU9vqhK0xERS7ODVta3cc6qE9G6A3KARAtFJA
bzHaWPJ3cMu09OL4lq0EvA==
`protect END_PROTECTED

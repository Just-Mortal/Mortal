`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RI2n43ljI3FNnXcdveZG2G7UWbdMwlUoUSBseLV3jCGlwOYMfJGPCCU1DZqn54Tf
hEWnHKnClXoD9JrtTZFMlAMkTt1siEKs8sx449YBlLfbXSGRDK5ppvRnCxRFcut8
it8kQP1qub2W9L+iPqOdGB6z4gC6Kdq19hE9Sn/Sw+vpWMQOoWPeFuMBQoILzYvz
OgERUFWx2MDdaTnwSPzYPQbKCLDeG2PL8tqcBgsdjgFjycUI9iHcPpuJrecJo6iQ
za1Mm2CXqPjOyflUPclUoVh0IypfbkoahHgEIVxv3KkXRgXjgEwgKhrVjAbGCvo2
BYKcZjNo3b2EiJf6Sa5KHCV8+pjDOZrUxdzEr0BY5r3hsBloQfPWqUnxRQ7GNcQ/
KLm3bLoOU8d2CiZLoo7uZ/KLQtZM7gB2ewuaTyFo5r6VFMBEYA85G3yi/Vhm1N5g
/szv9IgDfypw88dFuClR8pR+55vXTNXeA+eyeKMQ3G7jpHAcs0SQ1lGqeN7aGL4x
Wf3XjXKW2LEukf9A8zPZkflVYofN1N4ziNQ4USM3PeK2Pkoev8YlMHElLmed+0O+
Sb07cJsGFN9I2A/bSHQdTZJuuZPPiYq2CvtjXjV2uutJ+/l4A1ECbh6ivdF6vDpT
E2QkfELqa/qmp9ji0yjGV4GGQoL9rHA8gREcbYS5fXGnG8INX16MTzX6bs29OEbr
Frrqw/RMXiRoiZBGRKx19jpm2WYimiL2s92hIgFBQluDxmExpI5mYJ1JOVCrEXEP
v+XLw8RmvlHKxQz0730FuflXWWi8xLT2Wce1fFnOUfB/VGYwDvgufZB4VK74R9Wx
FrKsjIOkCCtixV+JlvWGXpUzvn6TnNiHz+XjI0kMpd1g2D7xCtEWFDwJuf4XHLSD
7pScIZz3tHbyudCex9M1aFbFpK1sEmyqTgisdwsfZ+aLzxXh74e3nq8kmLQEDSlC
`protect END_PROTECTED

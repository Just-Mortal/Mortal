`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z3Q3n+mjydTd8OmAMZ4Gkz6wpqL6Pzv1PDBolnUbi7FpCJcdQabNWIfS2bzucg9e
x2yuFVVp3ldc/q+urrcVO+JdDL7BiPUl5eIJy8qgVMirLooEWvHqaAlSHpyPMXg+
Dmaot1HXFxHp9/74DZL6GdL87vdoTz72EJxO5zDJhZbpLog6ux2l1wTMnyUbAKMk
NAU+Xa/KaCdHnlVDS9p4woJp8MA81K00p420JVtARJekW3zR59KZlR5SXlwqLihq
yShOApmxULQFzpXQlhh1Ou5tLBRnrfH0/ozaSRlLw37ZrAcfkn4OccuszGgcgen+
4dzjH3z2GlzEAPQoUXQwaGeQysOE9VX+Kx4jxRqN6rNG1eUaxMB3GXe9YK6l7gK8
7B7yhoRP1FbBw9SBY1C4+Dnswy0kJcWO7PiWgxTJ4WnlKjvEtr+Q5o2iivWTxLcw
JJLXZ/MqyZBfbY0/SORmRGzzCqdYDn6fSuPZVF0mDhx8ARPSu+AH4+ZVJU5XgvYF
HLHKBnODPX4IGd4Nc/wVSQpfHSbEhpxAq25jupu24hc78jS58KfaZVQaVOcABuzc
dzchCH6EgUHylBfT7SmlJ9/QCBq5O2EJiOLnI1BvuEFCQYoYll8chPIsw6bAoLc7
9gvz9Zk3clbHO6ZLGQ3sz25xnQy/GUrn68ZA1wCQQ1fA2b5+y/jyv9eI2cy615cn
KBVhNc+hu01h+un45nSDFGFX4EEdPFnOXCIowS3iqsnwi6oN7XpJxDgOrTDYPimA
YywoBsDxkdABRpRUao6y61FS9AmYR6Mo+iiVylFeCLFFN0YCFbRelFs86hEZPHwY
Ta1kEmSAgWyW4gRJQhFe98zbmxCZ1lMyTUkqZmei3Rt7j78BUy/jkTtFWhYR/8d6
ZCeQ7E/TAy1VKb2gG8KV3+39YiOmVbx+XQN9dJXkBzRbm4wI10GDbkvJ+BAPnPvC
dQuMnEsC5YBZctfW+MuWDLNefR/z5MTLyzAlUYQQm79vBgTtaYdK1CzLQJZLuuL8
2L9M5NKJTTgxWQ8YPon7uuBVXbgGNFPFQlUbub/YUX0g1WQHCAjhPqF+b485IHP2
Jj8517jgj7wHwLAy9an0HwwU9SSBRFRO+y8ZIMwECck1wIpn1VjHK2jGBUX98uvn
2Ns11D17kc8H4KzTcXWJ99hwKljWY3hBc9XmIu1z2vHBof5ekpyhjrCiA06ApaXe
KjbpewTrQfZsQGE3mA2dJR41DQ2vjzxHemzlYA81Y0JUyW0rFKxXal+FS1s9aNjT
U3QR0et6FVj69yuWrkq5KPoWycwINjOGyinZQKoBMH7mo8uiFY4z6bMA/mWENLI1
HITuNzKboJqOxog0LGwtsdTKlGG/LG/JfQMz0dZ4rEOEHdhe9etp063cxCPrruic
dagC9kaDY9YbGiyofmVTruYTIXnOnY9x/UwusdKh3ty7JM1RcZe+IE27/UVrxJJO
IZpzBTM0mR59Jg4Wj3V6Wy2RQ1kLVYXbWDPC80pbdSpbfnOQR6M/K3OM4o37M2/O
UAugkDhidlGprH8lWQ7Xmw==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4aeGFYnhh8yniW/nV3QdV3AMoLkien/6jiPgVa5CB+KMt59uDa624mtqPKfJ/pOm
mGwl6du4bHx251xhLEbvnesnPtr0PBh4rZF8A79UOyF0P08G2GL8xqvfsfezttCp
SpF4SaHpt0GNkE/yOxt6aT1wxgLQiH0DTEgpC5hIBwzE1kzrGcSc/hp/mLc5YHmi
gjRvuTFQbcbVWay0kw+CD0UodkvWUuj/4ANUL2KvPD3qvwOnzU58kXTzDylqmEjE
34V31fnHU2EiyaoV+ylW/vJkqqzIXW2CS0DUkiUC9r+TE5ZcH7TdkQMLZ3AIvjXD
Grvc2CUBIan1snH4Na5LrLq/H/P2OXYFPE10AqeGIG+1ErV/+4EGtIFTYiXvj1LZ
xl3L4Ef2rhV8DyLGAJ48UVT99ur48Lc3GADW/n55llv0ONYXMzqiOrGdgqrQZ6bd
37OT7MJlX3z+avgHsARBxkXe1nBmQlXaI7BCQ3Te8q4Uj9qrPfMoY+l6fwUBLZIa
0rwX+Lf8KUZSRV0ofUd1DQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLgB1kDYFtn+wtMqB6DQ3QHpfBjNVPuyO/3ukI10avzlpgbe1hFRA9BA2n4Xht24
F5OK1ollh9ULovNZ//fzCoQfcEVyFiQ6F5lKXQFKJmBW/7SWTIdIrSe3EU/fUb9M
PeQnGoAaD7lGHINEpDC3XGRpi2DuXPqKv6jLUEEkyohR6alqdCsScPxCDbLBAoPH
an+jeF09HzZhE2t7qeTlb3J8JtuSRUrYcDJOi/e4pZ24cm3DVrRqZF14NLImYKEp
Vsd/JA1g3yBKIJZx2IW+PuSyAwoK/N2kaFPjcVsRxArQOj8HAw+rJ1GluRIgnckC
T8NAbpgS4plKB0rWVRNs1j5/gs/d8GV37bCy52wpeER6MAuxgN3GxYRfAwvrM3hW
D+U9OZyI961z9kmKfOWZB2OtSEvAvJOhaN0zMykbSfYkX3kCvUrJrK3Ge7zbU5iu
Et5cYarIEx3Qo+YpCNMs7BcJ8a+9P0ZP3ojoTc1r2gSPuhCSrstTjp2HlqFTzCjZ
KA8blYVk5Aq5RgCF3YJSsoa6r6FkcAIG39ImZUdRjhbCjFIzF1EJOzD6hzgJ0JRm
m6ECwzAPWZm69rCvoUT3ZRYiDIOgHryqVROTSFR1vw1zvBWT39Pxqa/CwUuczWgC
zZS3UQgEQqodnMXdcVvSJlE5MqQkptoVQ5TyH8T3fyni4FHKxEP9hIjkf5UipZCH
GO7U6nDUQ+yCYWK9lqYZNYvdhekxNEQ6ycf+ftkk5mGb7DfaEOxJqh0icb6nbsRp
8K/KhrTOvFZZnm2aLfAiV4uuYtCG5dhvFdKFacuOOU91tkaiLN37qa6oxvMuuRPy
0BRAt+yXqpeEIjR2b7bsxc2152Vgp+aF2wOD7CdfqTTgAclJfMOZ0Po+OzcXY+EL
9Au8WJ8biYHpSrb2BK7Uz02P5f6F660L9iYHx2QfYvQ81WR2y01PTdOGsfHFU8wG
AE68Q6vIkOvImShzoGJvCKm+JH6lQKx1d20yVlDNe9nvaDezIJV2PgXqvGGMSHU+
w4kdZdsOhw1q1z5wpzG9+wnseyAQfRS3srBM0R+u/LvAacRxmgcmrVqDaKx+n4uS
`protect END_PROTECTED

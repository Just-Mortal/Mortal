`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CxJmTr7wYrGdqMWg6x2c6wBgMdC048ez6gExtu8Ae3sMXX3lWw2NsPyXu1jwGUer
TUrHedpMnvdCX8l/SYdd75cJ8BphhWcCVCVjUKmCn/62aIOXY31hwad2Mkh96Zxm
5j6OtzVoVfOaQ3aNkCiUiTPT2pJuRDOmyeSFemqRhewY3nNUpDFO33Q++AsYfxA6
+7TeCNIizOcRF5+eoszbvljk25mpiAuxUAJnR9uOUQTI06L4k3fP83lIl0YDzEud
5YMj2rbyY3355GquQ9DGkbZ6cIENdm98NyRCLoXVH4vuy9R8fS6oNuoORjmlpZP9
jrfVUNleMEAt9RaYxeqJg1UIviipEQA8J+mf2dDjRmrZ5pRSM10rJK9FsL3X4gCM
GKK93qrm3A1cJANy6rlDdWwSoycFmSpmRjjRS7Cr0LmfHKAVZ7xD/JsYA3Hu17zH
TuxS8Z7eZAha6LbGYn8qTnrKCG20nK2SCyBehWx6I/ZMWQNtgf8Ci1vLMCeQZVgd
6GTGEJywrStzgkBQI2NPxIP/42ONE6keoqIgSmYD0CK0q17ClpsvGMqt1YYE96Qy
xPwlwB9Y4v0lWE4NLLzyBSjlFu9xe1KkW2Qyhf/qldevBeah2UMwLCy76Bcc44M3
3W2n0hRGsoOWqpSOD6okRfRMgnYQi/ubY+gOVC/uUUOFaHJgZjpv2uP/ZTUXeMFJ
8mKLhdLVWLnpyEmmnInjbbItjuoKYvMLBtMu6AeqS2/zpFm2udpEXrnjlGSshbic
m7IYCGvSw/vfb0xE1lQZ3UleQqsZtxAG69ZUQFGFpCSIL0atLks7dTyGPoFXQ7L9
eacYkAre5XBX5HZv09IYgx6JrNlMfD72p818VjmwpAmolygHmUzC7nAe/iFeFVHm
tENzZZ6pUrJKBfJf+i0x2xKe3cSiytX1Vj+MY2eYd5dTayoShOhp3b05kZLseZDa
VjDpdqpMqTKBN73aPO8S8yiatS1LTapRIuPc4dn9/MtJnsz5WB7LaiawfbMKIb4o
6skNFIHEvNlF0PnvDUc1xE9pBSCgJkw5jjVzE18hpbS0lBd3mPUw0SIbjwUeCnOI
4Kdm+QYoFgYyjNs/e2ZdfceQxnysqe5e9Dl6Bzgf+gZMVhzSRbBpgJNVmOSR5ioa
38Yf5aUs1x8M376otWeoI3wmkFB7SfjLHD31tSUtAMeVThsf3OzbGFuyWFx9rPvI
X0f1UoMMoVcEpJXHEnQtwN4S3zf3+vGRRHPvS1LOcF1bGTMSUc9dpUMTb/7DcP0s
+aQUYrImbr7G1P3YRB4L15nOKsaTJAvMfS5VbrbzLOLI84CN7ScoyZFJfHB1PsY/
VgxugWDjLCmjrj0aabn4Ch+gjnYI8a4e2FRuhlDqxxRLRvZ53V0rqFeDrxUODX8n
TFBFyeMI/vwKu61GVH6wHa3KfJjbiwP6cyYazLSBY9xvt2fkxXJAfAZYqko47mlG
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hhwagf6HjcvqgrVIrbwX4n2VbuezVx4Uy+vqtG5fBs6WJUWtYUn3WL5pM97nl0VC
pUcvPImKiRsnscHWz22YyU2NF995i9qpw6qWB+C4i5EZC13DWHKhxa1jiyl7tr4x
86WxSQLzs6j+11B4pcLK3FlMIrimOl1ExOBszvj05rEl6aX9BCQwsl/tst8Ynnw3
YVq1mPpAnRuNmcseWHx0bTZNiC7LBhyAFdeb/YkVuGPunCt3zcr+Pg8n3DnsrAIL
upnbghHsPWGZdzAdTBRkgsc/lRT1ZCzYl+bKM1csHGiLTfzHSx4wD+vWM3IyKSFo
5yiZUiVe/2XrB9LjKEAqT6zKfx9duw1qr7K4pNeQxJuIznrq5MQmcH2/wSB1mQop
2BJH6b86M8mnXe6sGPLpBMQ1hlYzz117TFSOL8XE00EAFfAVxMMLN/qxiO51APNK
S1BlSW1vDoWrka7dqc4y0y1s1TgRu7kPKq/+1ylgL97VWlJkRrNRrUX0nhQ7iAle
4zkOQ7cYKe5E8eXHDHg/UICrGdI7kEPKkxDdpfuB7FaFFzNkO8uJeD5GwXtQkEho
oklk8AIm6NdZIUubJW57VIC9VkZ21TGvMXx+W5QeYTxVNrE5W416GElfXZYT0of3
O2NfwB+VgnwOZjdJzvsFClDBHZCZI+gcWFf9g3xwmieNrwWNDkhJfnbAK97ciZDx
GpFzsz3D1CP4scOV5bGAmFrQiMPr1GvYpZdo7Sl7b24YQkiecr1bYUSdRuMVK1jY
mT1OfSRDilS0FxTBtKJqrta2uUg4IYR+CFtjSMj3yJXLLsG00STMb0QOU7uP58rR
pkbFoPVCADG+CIPwi/fxMt/PbBFaD1I53XOnd9/dPtX8ySNNcN/eCquPfFFAFmbr
V77Mi/mrZwbLobuhkTjlLHSA7OK+2JT7LX84AS2tYVLE0zb3EJAWSrZYN5XUff1K
IKzjiHshqIzKDqaSjHk87ftdjq+dJKUxZl4sU6jbxRrhY5UN5Nlq4OBM6P4c0lKL
Zf0rs5vsWg9QeqDc5ZEEp+jCZ/BApCj1Rffa3Z3l/6iOsSmaAAH3LtdaxB9rAuHG
bpENdZcHSubIDz6QKiOtD0UA2rgt/XHbcAh9SPXgsdN12qXG7rTJnAgNv+J6MYOQ
Z+jcXYdxNhvylEmCedpf9eknGEl/oznWC0px3CoZuF05qjiUg7/69RzQP17zUS1O
AW8qQBe0xbu8kSbiXpcwRt+7ivpwhf31ZkrtIw24DxFEOBs2tHaBRwJbdl4gx3DX
f4oPpHliuW4Yy7kzoiiNMzdPafxSRP6zInqN8fAH/IMxJWzfzJSLNx8LX5UlxcNz
RuVtxF0c3JlBjFF/zS9PnA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWAmwLyGa+ESmTOGp+/Sl2lhI/eu5L41MDadwEU5aDrCgpki83GLspEeVJ7tdp+G
cMnX23V5KCZA467VE8AFvpm6dNgQRysCP3g5lPSAAUZ1gX4xniC2hD5gYvsVcQOu
Tk/eN7DWR/oTTGnrqzksYWOHuJwrdXXOzO4Lcbkzmn+yV2GRMrrnWfVIz26j/rP7
uLpfSMnnjEJMVRTlKFZuU5YAuZQsbzNwfHAVI+tghOSztydfBUmHmh0s/oBiL+Pg
1CuJF2nljC++3wHeAC/zQ0DLVutm3wp6Cj2M4rDv3baIX0HRiedc/0wgeNOFhf3O
mau/wd/o4V3A+NpSpttjck0VdSAQnMo/fZvGnSTDRl6bP4R0vq//K39YyYsHuJiL
G1UbI1MPMTXuKkBJ07sm5SC9bRycMgNjdHV/rErXc+1O6gqpP/B+BXoyVN1tILPn
w4dYdEI1AV4IvTllHmnxI77EsG5JMgV+NRbKCccrfZIUhdvjE5W9low0Ya198NGS
kOXlWxuqyKTtnL6qFnkWGQY3+9J+f0WXMCGQZjgN6dIzbEdJrp2/oCpTup+q3sxt
9dB8H+qcFB171x2P4wXfgMnb/an/4+dgEhrFfyoJrQj4FHLKRF+qDFkPYUer3q/v
ImISpxOwnMtiTZ/YM8dNrzzt/SaK5V0ffDRucGeHT4m0h7cOPW53tc73Yvb1QfSP
np+fhHSp8mcJP7v9UrO4+rg82OnN3lei6ftXCsDEmQcan11OMYd6tJJ/e4n1cupb
Tgcbtm/EIkRGzk2xyvTThv949RPRPxYDR1/YZlwif9FE4Qn5TAFlO3wME0oFabiC
Gi6jAm3hUgVf3KJ8FIEcoLO1drYF7hci9WWbNC3ZikpFrMNraBnsMjKYiU8pLcsO
T5hOcREhYjMAXh357ZjAoJTtROOL5Qh7RzaMiPAzhKsD4O45N9QeGk/HYj8dM7MK
n/tCo5TMKE0k6KxZlX/MdjOvIbTazdxjTy2lJGdhu95bxX+4D5bqaKlwmXKnuPJI
m9IhFqcUVqTJHPh9cMgLI29+qtH/7rMpi/IQHVMhj5eNgRNsEpRjRi2+LG7x7z1j
2Iz4qhlc+0gJw4MrGNyDZctnGnesA4+2ic1B9HChvapoXF3nf+QMIFJlzuQ4FMbR
r0kwoizX8F0tvRXiEJqnZGTwNNhoM+Q37BD4EpLv/RtNeOM0m4ixZCaq4NKz9oBS
ibUvwdGi3/RxqumEfxIWVM2AGiTR5ZLS2hF16mD6sJB3m+s+lm4yDrmA5cOt8CKU
OHYAypOXbLFBjiCQJq87OfPESVsRxLGksbkiiFwIwMeEVjUSlcXWKEST0s4tS7wY
un4NpSh9nxwdRg4fuBuUuAI9iiZwO93vd45D8E9wJyr7m90H4LVd7GFSfWMJyapx
acGuYu1mv/KaDdgrZuIePzUOdO9Jq9qPGIBQpoz6B4jbIfuaxg1WxRwsO+m2qIv6
16ryHuHCLPMcKxM/NCtzRzw6fo50bhgo8xemUiisng+1MgZSUYNekozRfAw+NPNV
fnx9zK2UooxEfp1ZLeeYeszBMOBTB+FKSuWxD59a8nyYvZ8YyOroKkaXwnw8oZH9
JJSQFynLjn3roxlCmioHROCRVz6eKWGo5yUGDXR3OeYCDsRgRzyW9b407dHckPUz
K1dLsND3TEwZwEY59UOkJ5rm1rnO65mHxZ75UfnE0oQbQhU1aXH7EHoRlvW4CBS/
q3OyjuLl3Xhh01CybwwlEEQw3HWNd5NF9YLAEEeU/c4qQ1lWmBNSEuMxWUrRig01
F6tRx+0jW5ruyG59DgEvEWBuB6gi0eOmtMeP/fz107nP9N40LDuBG3dVwxw1ulVw
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJ72DvTOsJoclReyVRRg8JM+i042VV8l9rHrJJU5qmLQR0e5oWRjssbQ7xYpjXms
ZdTnQFtG04oo+NUuIhwhjPqW8JXeecwmAm514DAFPzwZqiKxISbRrvnCf9t+ds9y
F9ipPjx1ckvGpObtWiVeDvi+69vd2GJqRYaZDMeVuP5CEo4Hzql+FEXNVW/0bBcO
q3aGbiOY0d5cw/UdZ7wSxzt5D8FxXujSvSh3w9Lq2rVsCNACwtrIMxaboWIsi6D5
O3z/6Rbr6RmiDXC/B/p1pCMCAtlMZEsa4F+u92eShrDfvmbLV6p9JK7Tbe3S1eYD
5BUFgUtW9vs01YSPihNbfnk6tBpdnfRYNFsN8nCbR42Z6G5CmOV16HMtZS3RhMHv
Zuye/dUmMmym1ZEa9zycxiQlXpKuN9J6L0oug8u3lnQEkV4M6Ti+Pr0mDOhzJVqx
mfK8O4fTBPyNlPWnBQJx5IR6Iwl43OljAPa7lR8Ch3S2oBUlbARti55Q6C75kVX0
M3yQ5AO6j7/ZjXUlfHJDWOKhVqY8ZBaAwJP3nuRIDJSKaUeXCGLTzJPOd1jhQ7Gl
egECVM9xt/7pm9BBwci+WE3oNESzWoxb/EjW5vlCGmrYZVlmyc2vVezLisg5Xo8E
ELcQaUmSIrExMbRxR3mFJ4cfZY4ztJHfbA6IWl9kY0vDV3y2JNHAKhAWgS/TKVxN
FlkVkXcpUct16liUzG0eL9NHRSjeYyru2KWkIsZe5hHKv8ly9kQ1VPBl/6fPk2QM
O4y5T+s0HUhnbahD7wUuZTLRtfvNjzO68mHyXucdTk6xIs1eGcuHtEZtl+0bpqBk
q2VX+Lljhaj3XvbM4BVAP41eExem2KKE8ywnjX4uFUfUhASy4jydGNJGy2/UyWVm
NR7BX5LjsR1/U0wblyQoQFqtuQLTim2OgrV/OYMJirHHAhp1dD1DEFbYtksdDgWV
uze1Vd7kjHtcAMtKcf6y2JiN/V85cmsElHWZ6Bdqsw6rgBshv5HbdYqe7DBa9nf7
O/fUocv6P+jt/hac9XlmCUMA5KFma4BcTVtGCxO19fL72zyko3efguh+A+u9FATt
zDkiOAc7Xl0NCNY0YivDnvTn/fU8tux5SqGAuci/OPzSGAhrNVjUkXX5nowA6PbK
CqGgJBV+x2+iqUMkKFY80dHIkykytVoHPBI7uABEGpGbnoDCgJuidifxclIA8gdN
+R4BvbvEfgY/7EtwoG7PxCjWWm4kCEPbHAOYXnhZB5jMXqgMHof5nKb8JrDBpOBa
YNWwcqcuiFygWbDEFn2mPxGaB/1lYiZRxHNU7COVgr9nd25JLhsEUI4SXo+gzr/2
RbtBDK5PSVI/2ixv7qnMv7LEbCAgvqGYqebutDxjjLGvptP/ScZWQtC8tcBNZWLW
PBfsw7XRtxg2Vt+Ok5YS8N3pLQcDRbgZP/cppiuggkIv97BwH6nsMd1Vay6VrCEl
vCtnyZuX0RQm/rFCWl9/QHWoC8ENECPRsw2tYMPJ77FnZuR4zUDafIqIhppBRmjI
K56YXBtlJsxgZBiw6J0epAV997jGFH5P9nX/eJ04bVas8qPNdkqm9SSM7kdKS8uk
TNTBiBOX7LrLCEBX8zX3nKhtaD4BTcWdAXi5C6/dsdIm2tWjIlk8eONsXoU7rd07
+g6sddFQczon0eFfVHhAYT4a3zgwfbTfWMtAooNIlI1+u5z0fICEj0xVy9WY87Sp
pn/Kmxq1XRc4bmL2COwksAtDWw/spAM2BuMskmNmaK9hoP/lzNXzpefxbzG2mX52
sAZahvJzNiXoYecViYnrTUWNR1lclzGbAK+/Aj0bHw7/WOSiH5gZQNtcSFom6BNk
LEvgkVb/X+Xm0R4tAIv5B7+Q+00+Aeos3+tX7huorywtXM8lzuH/zSxPPDmnFITY
lgZQzyHqYvbwQBAyEY7xmNSznVjMe+5Q9nqY5NDVoP9Bovc72bM4VwRlfkV+r0YD
+mn4jA0lGUuuJ68hids/ibbqtdW6qdKmLSDLOWOnR0GvgdohAkT6RswyTM7sPb6v
C9b9NOpu8j15n4W8I/6H/ZMD3ePLK52L9/XW2sDRsM78DIy3/baPrJNhjhJRjAEu
zJcJ9FuEFjwug3QI6vGoqBayjgRXR/oglMElV28qiD5rI26vnN0jF9ZRhIsgUHn8
rNY+iVJQL1vWsZ/Oz+/fCf9tNElVDDCsD/A6ovmQeEv5aH/9E4r/ISAAy9nIgHdq
H1pDE++WwnCGKGbD7r9YgR4X2oyuv7BF/yMM7hoYzoBVNip5JA1S1EnSPnnRmHXp
8ES3pYQHlBA7IB058R8WTtLaMJVkD0sPdItlhX5HFkyOCJ1HDe92b89CVVxVnXrT
SpsBQttYqLf5FZ2fKOvdFsa4S4Tpd4JbQjBTZ2/ChGbUIz2nXX23t0XhUps9FK92
MAAAfWmehpewQ2672cVH/qFg4dBmmPDyXprW768XOwbIU56meyiIP7vHE207hTbZ
sSBXrF7jJZ6vWkayr4blv8U+tvHsI709xHx0QAPV+gnhOqZPl1XVu6vaO+9fYDL2
5Vy1cCnnOKJrrgW9kaulI5neCKQg9pzckWgCqBpqtHzwJKEuJZ5wR06mo7RdUgkM
yoOIPXc+Ny74t/9v7hZ/8jBxAUtnoPAKrdBMV6esDkU8EgOXX2UPzfG8O8d6690H
r0vZwghlGRLn8Vcf4PsV8yBHJ4ztkbMaAS+XqXI5altUy4fQagycBio7m2AYcdtG
K40h/JaL8vX04ZhrxCDWNL2XuLZxQkoLCBIWHJsKpnbbrjiqtPRwCII2h6DDdF6M
rdQVKesuZ88FkHFzv3oXJKI1RCmDcQTTUFwld/jpDtPUJwOPldhffyaDavu5CtNk
7233S/f9c4+g74HGMevG7elWIemH6M6OE3gQNL+sZ4vbSGkJsBvyURGdtdaIjcvy
0XIBUxhRbhZqOKJq/t7c93WKXXtth6GsgMtnNyECwIVREBqzXgQSwTwZ2fe9fI0d
FaGQlA+RjjSztVK2JKW6SMUijKTxqR9FZVAFva45rRW2YtyuqNOfWmgc3FtcIc0I
WJX4XVVjl8u90vpRiO9Yp/UgdhnybDeLw1iovAYA5OgkdUdwORULGuHt28Sjo2tt
fZ5LYoYDr0xJ6RcJLzXl9rkzQsv0PJX1mngObX3zw5Hy/RrxVich7P/4+yg+8NeY
48ggNjLUQEVTWzQNsDVpeGrYCaA2PjuKgrVZQOpunP5MMtmLmxjIagEJeTztl3E4
6/kKT2Iq4xYu9i4MX6Ltne4S+lpCqdaDBK1UcpKx08w5OpSIDkQ//D1Phg+xXqxu
gPeme9G1fJa0q1n5fny7PD2Pog/db+/Kn0bL2Z2Nh6CucTmnBZt6GGjcuyYj3rEw
VEicVA8ciDWbKxM5idxmyjudOrZYBnoO5A+gWtPWKrHBOsvH0mygYzr2Uk9ioVz3
miIMmoG3TVeK122zrSTVEsn//yJsUJ5fIUt2+T2srjpgDNoZ4oRL+91P1GmpgjyO
Z5HGR/rSHIMT9SQ4R2WdLUSLcg9myrMtjXZhme3Rd9xJoIWfKMLFmb04rE4Y0RQb
8yoye8QKVqKwo/eHbLe84oWHoS5JsIpXXNEgev5YhQqltNJG+cMsOJpItNRx1UgC
WdAyWuL2o7Yv0Dp4Y9F11So8xk2aviquOJ8K4wq0KRDC9DitqbTClYafK4MYSQsA
A3Yg1UMtjdWvOnHX82vTuXVwhGERwQrT7mlfbaIFavPDq0youpi+NB1EbUOGoznn
0pi7ehCg8t4WV2RYipREuAJG1wB75g1E+D1hLXRwc7eqhdXGc+Wa1gOgHZn1xnAd
9yH/FU8xwiSFQEdjBqU11oXr8ZuuodV3Of3skt+FB1RUZuKVlcJLo5d2MTDADkE2
iA86P7B05NeaKoDjpsd2jcxS5zNfDksjrjsFFVYdwDkDOMVRA+m0CFtl1ObTinlO
KE9dL4HosZgHgIkjNestjFkc9hd3ZfHNnmhdQ13JPV+pHR50NA1AF0gFMJrKiMDU
Mxxrc1ruXiPnYSHLGbGr9722vqWo2112ZOoO9XWzVkOYQ5FsNvJLRpYaKdb1dX7Y
RlzGEaTniG1WPWuQ0i2xLwVu5E63XrDVOXhk98X6avcu4ZZjqUMvzYGJPET3CMmc
4KL9Kt3ZjP8gZTR0OGpkRb1eoj5bo+TAOkroWUY8xMfPXEwgqR6AUYnLdyBuAgLQ
CBoTYO1uBE9wNzGg4/31tQkdmmvK0p8m078z0p+Ip4oDo9TAPBorB1NqgG35idOo
5Ys7uuoO7MK7kABaasRsuqjqsTOFocPR0lL7nq5BsPw9OSikZst3nLNzeRzinwDn
eAfp/aDuAcYK/Sb7qW9hyfeA0if2bjq/+pMtSUoKxmZPRLgz/+pIZiQIpyAlwzMK
KbKJexS2wXLZ2ru74JPWynP3iOwxmX/1reIkVvNkZ4JopszshLUF7/Eun7FKr6Pd
iYDwQk8ax4IxP0w7ON/J8hUdmOVErRFrNUKhne0Es/cMdpVwOCV2W/061SoWOO+L
3TwpwW5IlbsSSWMN0Gauc5vCnvUNq7Tz7JATMnzHMHxJO4LtVFtQfkbQNsP3us/9
8dE0IKvl5FAzQzOSKggc3UQ+jLp2OU2A0e+tlg4gceIQSj7kxRXhEwT980GkQN69
8TgVA+ofuudtxIleK31RajCGfNbADFQml2+5tMlDdIYd14rWz+WBPCGDPtS7dBpA
tEnkhkC1tTDltegje4eRXgkENPYxJ6ZXbw+hcWs34ENLS95jrZiVLVGHXTehG8P2
LkaJQZCkxxYCGLWnCUTxfks51VRWd6HTOh6nfGTKwA9/wZ0WGaMl0DCdo8NDqcMY
JLJVTDhc+sLnv+7u6u3z13RRQu7bKvVGhiE+YHxLlX5SqARqOXZ1E8FO5WerUtHv
hQmNQt2yZQ0f0g1zDfJITfgzh+l2rtnp0h6NAJgWuCgwC0vIzRdtJgvVMQisfjzv
ees4tVxAXmoOQK7xZULkDZcYc7t8lcpw295/53XM7pP/jLyEDdpGHkH2c8jhUS22
LDMKqxW/KhvYBjpa6va/NtGct5kPMS9pS0LE2Janjqlves10lVoc4xfMsw91ZmB1
oskHUKEdTu6q/0dKwRRAVR59iCPEaW2BkpSTW1+kJEVrhBbceOO5OWS70zH679tM
1VAqwSchJXLsSqMtHryMbr7hJu3Gtwta1zuN4E0txPYTbf98wf99tvTBaEeGFpAZ
yEg7Eg9vO4D2bN4pMkZpbyyWiBnSd+2ajgBwnj64wKHCmq4HAKBlcwO8KUgUAC2Z
THAvtEyaAwR1KBwHVXROsOaDRQHQmx/jWW01zakDcvXtmMsjmnJsdyFzsjhuzvpr
zYzpk01E+2MN4S2n0QJLgxDR+tLSh/wxdOltgvDxUT+/Hhy7IyZL0GrpCnDk7puk
crM51Qag4kAnNa2L+tfKyshbmRzruIyY2JtKB/PXW4UtD5/DSaXklKYLikxxac+z
G7Qq6dieXl3KiWkkSW7ar2CHJWUJoKDGELyJOsq5W8BJrp0spj7TrapAHpw84Gjy
v5xsYhsP9zKNSzCDIJpMYmdAb63/fdfmhtfCgk9MCzOsS+wWK3iXRPFnV+apabyJ
rgwdvWqAJkcEvZKF+/xLwQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+J2TD1c8gbnQ41+5NtrBYMsEgiLjNo/9Vncm0L/0jU/qdGxb+7WragWQTM6eW0Zd
W1r+ec8b4zDcLGcFSElW17S5hLLxrbelG/g6x8R+DjF8RAVH0s4rgh/HWOw0VoCT
fs6UABG8fIxLv4ejPbldaiwvlJzWb6MwDNgJkty1oEisCfDzN1j2Gca4B4Rb10Zl
2hVNjj1rSEScJx0fyL2Cs+qPS+6fvKpux5WfwNDaQ9zqsd/EmIvd18FfHSMjZkjR
T6Gh7yuYXaH/Z+I2glhbviCMVx0NvXSoBqOYd2ehgoRQzFUe9yXkLbhI1hO5euFL
imP4e0N/iR+VVb6LR5tFtXPNyzP3UKXhaPEz7VeXhPN3qjhAdZazFeB3S4RsdYxr
4ymAgFfrEL6d3FJWbevDXJC7T37yriTtYbTDjTBLHr+mpZQRc79KBSWtbMh6DD/p
MCwGt+HN0GkrqSC/hlmN8YQ001SiyWfCpH8a+xvYjLhjUKu0xn0hhLGbEsqt0M7H
KSIoCOC9Z5W+8saxrb2bElwtxmE2q/9WpiB1tKwHgPNF6bfKzRrfYwuX4pXN7ktP
22S2vy2fUtVDuZJpan4IV0k/k2Nj9IdNfzFr2iVBjnHZN3QhUAltFNzjGgbdDkTu
hy0pA4628HU1paTuGhI7y9sqqgjJSc6+Y/v1mAO0JWb7S10cp3jMzsbnrRzlfRQZ
SYmW8fZJTMeQKDvZm9ke31kJp7V+RDSuznjFhz3IUvazYUYTDxaz4UjkfBdPTLJz
S5wRtW26EagSaNbe28nztreCotwfetz/cwY7rAYF+J5CQPVFI+uIGElMyhP66l0V
jJ0TAtgGzRhvL57bjQRy46ixJRs5d9RGx23fl7re2n9U/vO8ehopIbdd8EgJoM4/
bSa2Su24PyTxJrZpf7IUnDIY0UXzzcTexWZhIp3KxtCFUq/cxQ2OiJG+/ywd9Wev
04FCHVARYp4gGXqkUbTv8Nh7HD7Kik/cW+UboRiWuRvoeLn6ZCapptjBsr1gqP0w
RLK2T+1RjuQzvkSaY5REZ6HRbqgGn3s4bdpK/flWMReOJj8znIogP7fg1l2FiYWV
4vuKzl5NOz71KWIZC7hR/mSg2UQHkOMvPwcuJYbMIOXtwnNnQOXxAMk2yBTLWMcE
robKRwY4y/VTb8qfYLvFVw==
`protect END_PROTECTED

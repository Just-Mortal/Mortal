`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/88My8MqIVL0MSbHw5gJ3uI5yK+SNR/cPmCtadNGeyM7SMK4jy9zJmwRqubOYfL2
HqIIYmMP5DM7TRk7o8Hcj4Kw/4DB/rOt6srXpRvs+pSvulVSFM5YgPSEv6cY/bEt
e02qslaSYazqoB1DoYwOwQpevTUAGhiRLMJ2htlsO9PhxSt7PukIrI8KXOSjCd7q
YCObw5RZLUjq/UNL7JszLJXDSsZVxDpbjzKSZMclUsYUGXeAaOD+XRJN/LHsXONY
O3V+3htLY6GeIloeyLGNgmYVN4NDGkhE1FS00MG1W565aEfqke0mtFAiGTsv3bIJ
nPX11fS17bDHX45BbTLoEDlHbGKTHJ2sx4TMD9BdFpi9QSZbx64yeTixojZyhSXz
sqNO7RcuwzGgXtvG1TVlNC5L6PrFsiVC9gQPKl0vb9MXcPub+ShAVX0RY3iqig3U
vy6cJXZehIhBgNp9C7EHyxlHnAYihoTO0MwnU1499lfDJvXQ4ySPCwomVjuQIr1w
1AxsWOX+MD3NuxsvQdqm+6eRoG9e6x1IX8kJv2grAQ8o2BXgNw2oHFbt4QMEvrFb
fuYT4cE3enu52dzMZvtrROxFmmthuEwDNORj9bN1yptkA6hKbSt2Q6QjQeiKb7Ha
l06kRY9+e2tczXsYUHzd7R+GGziXghA1Uu5rsNlhM5p/7U7ecYqgh2EDxgWnUmUe
zsfCtFy1KxY2e8CwuYy7jJQnW1gcmBebs8a0f3z5MQF01pJOi1LKRlr4GRhT0Bei
6VZjzPjuviNJ8ItV4vETC8BqtwcSuk6VCjJZa0npcsNrB/f+SGmnHAFtcvOTFHLw
I4ma3xLv5HjzXTrHJEi79S1lus/vNL5m0W1IOlBkspKFCHrJt1zkAOCHLlzN+JNY
F/L1lQi7qcbDIW1/DDj+0QvGC3CwAGR5IQFSxhL8b1MKc4Oil9UdTXqOIeoPoxfJ
mdF8RfVjwZv4Iz3oM0h0ITBOPUw4LWlgsJ1Qs1u0zDcExpUeugyshfLvnNn5OcTZ
J+Chp7xRzouTIlP+oKUBZO5RnWRrnH/8ClLpdhq9iS7pCxjEPhLCJpyqtphmA1Kr
aoDBRrzIb0eqSVQj3UDpVHEmG2WsMmDNXUODm/QT60wqA96E5kW+2te/O0V+dRaX
MjtIWFYUuHHSTJ6/361A7J2VBVCH9UZzUJVAjfD4isDO1Q4srOUxe3RnYacxRluz
D6ZvsOl/oAuEwC24U3STRA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAFT6Wmx1piwvwFex2wilj2JZifWQ0pXmcOzT1TT9TGR1BdE96e/TyELiu28zodJ
2fvdFXVbUyEG0vMq0gEBZU/q0y9gn9DLcmGn9o+uewShhRvb2ru77m0gHlDhSJhc
FIof8D85UnVU3k/B737eKcKr9abdrLHPNKEOEwnbVuoT7o+BgcaAWbmCAQBrwFeq
5CmfjPv9GE7NCnccb+OKNXxsxtO7Ji9DxjJubWXNcjMnYa+MsZQXagHu4ZVImUTw
Wm4fa/atxeBGihF1hGi+1TZJO5ttc2yCmoJFdoJkSI42eKlO+f4XLuXlUT+CX5VX
7qni85zXe5z7eu4dnO+EKNsxRROfYhe27uG0OkGy9KmWFZq9qZRc1hg6a6d5wWA/
WK5im0XZmiHyBUjbGZIxg1s5DC44mHj5OoDnMjovKkn778ObG5Wd6hXC7QyVQoEE
M7ap930pTlz1zMJoW2r2o+E7/FL1NK1AVnZdKAuLzSaI8tBJzwP6kJdBL1Eu7o0N
1qpFbfXwji/Cj3U/atO+UG+56NH2emDX2TqBluEeFiIviwEol9g0kRC5FF4Okp/0
RQ+wcM743cWEZ77pxV51aGJtGalUKYIvF5MySvyAMRbQcRoyElksIgBNo0S8KtNY
XAi8EOlNmOAlU8ZqPpDTW8UQvJwzBmiCiU4Ux+vGIpdDK2YimNzWLpT2NxnHwkgw
7cgzR6C6hQgP3m6XD8jWlIdp14r+UuJx+u1YAZVUV1LKpj+Af8oOFu3n2R9dekAI
h6yHEopLXfxXDPS/74JWKwq94I0T/kgnSHxJZIlzQAbM3XkLQ9on0o1DHKXHGjP+
2DZ8vKVwSbmneFaMWyRmep8BkHZWvNl958LZBmpYeKU1yD3B4tpQBGp/TJdTLXRq
X/3Jp4QjSLmA024oXEjaLEnpMdXHAVZ1uSQoUWtgCJOQQ4IeeNrzmOKjk33T8mYU
efO2yv4SdHVk0ndw/Y5tnSlicJLFSpYriD6mMBfcy0FMX+6SRXiFzcHi0b8M72rg
uGa3cvYdpxf50TTJ65G7dZRWbILWIVA44vFXxplQ1pxRI1QpY9EacBQ63LWnEQhs
ib2+6WKRZixZENKmjdkmtM99ssYohMwwW/H4CNwHxibxVbKgFLI63WKrPRV0ajxX
9ci8v5er4OJbTWJ/qAPydVaoc/mkjG9kn6nMFYd75pMaS1BjeKG0/e8nB1isEMtq
VMAGHTe45CjEl+BKSB95+ChNQVvD3Gb8rw8Fpt8WOxqOq67jYw1fGtACWmyIOeoz
k42jVFZWbuyW17LlRMNZA1qBhlCfJ4Kl8VKbYSDYGTcihah0zIc7bzA8zsFEnX6z
e8/Lv7uqyFBgagd7p1lteEA/mAZQGXQfZ7CYdDwotmXI+lWELJJvbdTMohlHVkXR
KyhBoobbKk4dlPZu1saZtGmWLJE/JKD9IKfCAoAuBdSpACnnxF6ioT3ClIGWvjLg
wwwEaR6bFyrngPYrfJ8iNp554gGb+bThcokbDAxvztHW6v6+jmamU/dAGceBr6fy
OjhXNW5hmYzoKXOh9eJ0uww/jq6QpplmBQlp6zMlpKS3ORoHxZBQkZyzoyGMXJ6g
baYOs/8Z4XpR5VnXNVrha8ZFny5ddVYc0Kw4U/S4DtHuXI6y6pt0l2KT3ClYbHHF
ng0cdrIQSToBuBD6jhBj8uWlkHO0ePo/QJuR66CovNadsSouoIDeaO1SGBJ2nHwf
iyjnJ2ZNcG3zifnOYrhKWmwR82MbZ8XB3N/VgLoCCHRYPxiXn0Jk7LcApOFR9vrz
YIdZsT54R9QBbG4ELUkWPi/Mc0sijjonnjrVPvnNFBfgPIGgLX/LbItE+FHWeRWa
KGfqXtklv6BWebIt7jVqfzL65PY1mxqWdMmEGZSDkHk7mwGr2im1rJ+GVU5PELJ3
VP8fIMuY5lA8HtLBBYJgMDVDp6USgQ9E2goLhKIKp/vgAjhumXc+i4EuUz7UnWE1
ntW2ak8Cizr3KoPiSs7CJXxqzlgjx3CT6Wmd8FoqIu5vaz+hCLpwbxYpeXxIAgnX
Jn+TB8iZMdrJlS1/5/PF9f+e6hUECtRdxOFu18vEZ/W1ZUmDwAj/sepaMrQ6VSh7
YN81gXxNreCkv2cf6y8fTCDD23Vv9K5tmLfZhDYWmPAcO8DAiXADkx7XaLd02vgU
KV4Hbz2vskPapThiHbAwh+28u9QMpxX27IMbYJs8LOh4IaN/HUDL69ozxVqljAjT
xc058IH/m62EdGl5blrKN6KJPgZgtjqkUtNLsP50ok7gYSbJ7INu+c5PZg8ZoDMv
MpiQqTfHSYyU9wQZCsFrNFS0CwZKoT6bdPWrHV5PQywmXiS+ieBe6oUTJo22z4iB
IGVylZBvyD2a5UjcRXIReRXzfxMKwRsVNTkOt9CPw0z2ss2GAgoW1HJVuzAwtJz/
Ul81/IeqXngErPo8KEbK+Q23aaULhRU3HkV0RoVC53jeQD2/MpDO96Ndrpe/oxZi
V/FMjZiiN6eg9R6nxXCjlL4Hgk9nnatZJRzESzVibQK3rtO6x+Q9fccicNbfqI7/
0pw5te7cztCu7+9S8HgallCH9DAFCY/vDYX66qwwNP0bGatyTcBsdkmnRshIPcq2
0UIEQfv3IpB3Pqh9hA111WTfME/Iig+ufBfG2S/QKVI5y6ARgYNSm/al5jrrbnhY
ctmA+Y+a/E+CMjxUC5eW5dv85v5eIh5Tz8Te18C6WIkpCkZsEfjANTQjDH2KBBYM
YJ2rbjnnzQr9Cr4/OLHQ1g==
`protect END_PROTECTED

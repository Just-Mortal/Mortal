`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06RaAL5xA5arLQWG6uADAkkwRYgHqFhudE7KLSQgJSxYSEL6aFxNxDSaQEtJfz2/
H3H9jDSk4+20z+VEKwcHS6n8XBn+1CB4IWyIx3v+xut7o7KUjs5XXf3cmMVhxv9/
xBaY3LDaMMCJbWGKCLUfghFlJCyDumlbtynMkwRa+sLAz5m+N91HDx2Wd8o5UIZo
xEabz/ieMPIU/VKNNtEbiN37h5mDO7HoXwdGu86xuxYpJVrkt/IlRsOdmwld4MSV
/LY0UlNAZMBRkkgci+jRQpI2hf6UVHifUV4+pMUfJt69Oxf0EZYSNTpSD22tkb/U
TR/XRRxZQB3f4R8Y/uZrNsIr3w4bErLQgOd/8m7qCib9AZgM8p1413t9dzXCODoO
GO3C+xIfGHm07xBusAdBVLBm4d8sfF7G6wbLEskjEvgjr0jbqNGxE9btD0HVUL+E
3TAktn/a39YRXsdqTATpK/Ih990zcDjLpHKjI2QmbS8w8shur4v7au5YESOdrxyC
yaK+54Ft01Ivpu5o1p7druEvkq1Zj/uTYiVBxtJc8KUr7+Zbdz0d/Je0YIARI9Sd
Y+f30EO15HSymgTCY3RhXClPRnK3RzhKY1aWfVIue4k=
`protect END_PROTECTED

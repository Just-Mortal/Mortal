`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bJTTr0uXv62B9KxHA4H7UlwHQrzk1yHX+T08Tl9dmSdDpQJoEyd+LWF0gtLPxcpb
fv6w3CHJx8wu4n+8i8N8OQbWXbBw6M9r09LzHATRNaUJSY/VnqN0ls1isqVo5R+h
ETCrX7ztjnpXA/WX5UebQrla4Kl7lKV/o7Y4qFxc/VdCqmO9sisLlzq3TmJfEx8G
qKDargYvBzYMoGKMAStpa9HtKXeXxBkKumpxKCkhaDdjRmgoAkI9D3OPM2aTrHnx
uenaheUT2g+noJRztXZwMaOACJynWDfdWTWaz9ggh4iBqCitE7MoZkca5gXhervo
fGYIimwM81YaQH4FmoZV8eca8p7kWF0/6skRe9xn75lnBtvNmbiQNNmFvCBTjgAz
FbLOzPRUTgVA/QdJ1P46VtCk+qHRYoq4DS2YBCcj1dxoNgNEudzsVkFzNKsz9iY0
o+vtkqA2mu4aKINfN+k5we30aggoJ5cvM3MqFeeD1PrjIwINYJzFbFUJKhP9FGyn
MUaekT4Vlu0+XoG/FzPz5GNcQWzcsx9b7JXECnwLUl7hQ8fxo1hednDUpmNZDQpD
XajEJXkzGAtyrUvZaA63XOq1NQFO/fl0Q5NFMVk4fdBapQxl/rgAq8XFv0QcIqAj
CbWXvWvYx+yXSyR2sVKmyFvLSfxeT7HLPvVpS1Y4Var2W83VB74SF80ghpxkVQxW
`protect END_PROTECTED

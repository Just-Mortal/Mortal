`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A7ios1usdAsDXcCemzXbTv0kX2HcrBv5Qe38+xaQp3DTe4BjkmracXZb0hemEaiQ
1trIILpUt/OftkOgX+WDkwVRqdMZLs+KzHmsQO6BYS+FgyyEpDsbRIjV340kuR4w
Qw8HLEIfVp3qZ/F1A2ZN1R3iwb1Dd/Q2lhpBqOMsx80imrhSVBn5j9mR8GwS6qvR
tWeEFn9jcpQ5pcuOUPYbRy0szmqf7cUZtZBSo3tQWNRJX7/C9gkAB8tdsxIRTZYn
anVps6Vk7fC8IiYfk/9e+kx5Af4uF4/MI3ACwu0rlIEnmDGblYyM+7+B9IXDo+0R
Zw+CYVTdT4Q6T0KD4ATwGvIHIS+1d+MaLD+s862AB9e/YviROfZoKhRoIXXxLz5T
FiVbMaqR49JfATIdt2elAj7TjV35KOQGd61Icqc3iNsyyPYPCcqRMUaWmhnKgGoy
G79rmXXrjYOCkqviRNM/6MFQDSl2rSuCitCyfvLNlmy2kuShDsvM5u0kAkcC68n6
hYgroPOXA8DGcjcFJyZl3LtjzW+be06zEtCt+bSkxofHAd2OHhD1lXuLJlEdFO7v
TItbz9Qj7pC/WL4plUgtnjA7b4DqV0f7RGKWvs9teiJtkLyEE1a2Jm/Srnm9NwDd
l0i2KHbM9AOuew7yLWC4WfWA/6hlDImyXKsXnGrqZsoCmZtzzsbgkgDoWh+Ak/gd
7dgic7pz5r0XQxBfo35FeuBQilRVTd6C1/FogwGMAep/DD5lLQOCNnyt0Z2SbrIn
ufHW4TKA6HcbNLI/Op5SGSWOIRwHZiB0lcpuZlYFSC5WLiE0UjbyKSU/tocxpelN
ijOmT6FOY6wZcpculAPq0EmpH2g+Cs7M/kSLvxhtdsky7wGpi1UIcN1RxUh+1fjO
H3/VJiOLr6heWZvUAB4mF2xfzCdN8rNDTdkr1BcmFSBl5PEL1StefDoENBRT7k58
JvTaqBO6WxFy4rbwNr5muPFLxzQMvZCI+lNOEaL0TdTpeD+ZYdx0DSbbSzM/q06t
3MIf+8fNGRMgiMcNKlJs5Km1EPEUvghyClttswG0I2yRiBjzE4mc3b5KsDtQIEtM
bnrLp8FGnxg7rcY5h4tr13cphZfmBs0nl/Yk2ILwH3vc5QY3bz6VTJa1kk9lr4gB
idhrWQEiHDAatLokx2HH3TwZkell4rXeNg8I15RhgjJbRQVXB3EWHbKUlu+g07iJ
l0uX+RaHZdGbrmjXM2HzkAYU/LGsvASZ7p6kzmo0i+JSl6W7scThlytSSyaXPp6p
KAZIh1yl0pYJSwFaRqx60+OtFNwbp6L0XiOJ4LEVIoVnPdbWASsyz+oKlmSgyGLC
4ggqW+bzHrMCxU4e+y+ip7/GX754s7hGK0S8MuMLGw/V4Ew3bEmrH6rObl065L7+
hVuI2fL4IGx8kPKGJQThb4+8atHFQJs3VGqpEr/S/ovGVKj5ooPaXUrb6PcwE3aW
n/ITpZzNcGdRSXRChgUG/aiRbpfiyO/QHQYXwhjqBfawoS53u/HLysZK7PVk3FEL
ubI+AD6X9Mo2QEBB7c0HyKVZ2zyCJ3YsPImo0oB0963hhL3XlJbi1bvYRVy/C3rH
Nln/aPCdosyjeDLtHSj3E54KS0i28Gqop2mz5Yenae0+L7bVhHHM7g8YLeqNJyw3
YjRN32Q7zLRfpRONxhK4u18L74HRdWqGkTQZq32FEpywDnNi5EsN6Jc1pjHG9ELQ
PqAM4GRw3fSfP3+RiredN+d4kPJYzUez1MKtHbB3Ni19Wju05811ttH/fh90opUc
Bjiz9Ptk3FuX5CBjy9vplYm9QCkITYbEJrlA2/XEBCS884+DPWw847UNoy7B48CP
AiyJtKr5H8soLhbmRgeBTPeDCBx+MEqSNKrIoKfy2/4ge6L90eI8gMG0lynwVKd7
HaFwNPmDTo9J3gWSP52xIZll2kD8smMVSovV6VDgHYx9Mu0AU+Rww0MxyyJkS44J
f/PcRpxJxdhncEKR9WuLAI2xRY0G0mwxgDv/7dH34ISP9EVe+mwzuFhE/h80lwKX
quOTP1WJp79mpImWGfeeTLDv4kLwCEqg4jv1h35refQAHH4rIPoUu2E+1uDhZMXW
r1YrHZXVo4Ox6Q6mQuaKSvtK6JQsKdOStdT9unpkVhfvnNu25N5accAzOwA4l+us
QNSYDfOmbpTE8+N2TiFnoYZi5iAx16/EG7YLn3dBfpYILsF+W6UavdJofWQU1u2L
ZT13KlHIwe4UKSAZjtBVpPn9GYKkDf0NIxi64VDwjKjo8YXeVE+TItU+GDGG5r/A
LwGTYUdbjadROy09m5XieVgfEIeuvyBntVFpAtbz4IdigJUCrbgzZ/iIYpKvTy/N
Nn/M/aJUkGHAyITLIanG8EDKoAPpXeHWTaM1/Z/Wppaj2L0mW3OHCSIVapi54W96
41oXkjVyYs/VkY6CZo39IDZk1L1yFSZWP+zv/povmXeY5piBqB9yvSXl2HGrbrjA
73KR6OU+UAaP6xwL8j1gDfHyzoQlvghJyCXzMy1EwdPEAdG9U4nJzho8Gq84wUmp
8XUv78mtuYJLQzSx4hdwJmIlsVQ6vS7IBoq7RnvbzF/uYW1/OmKICBIZJ2clAiqW
hixzdHY2/9yjIQDRjxeWdI2diyT/70PQJ03OeSACE2gVzr9GEM1Miwr75xXBy0Xh
bSSnM46AE9Y/NEV/NLO+cxcVkRQg9p0XaW660w+oxdgnQaGsx7XOSjOjU2hzVP5m
ztSJhrdaPMGGReyflCmEFHgRSmennANHMdwHrq5+ZOj1vkau64n6uHvzGyY30W3s
bSl3CAfhv0SZvMBAayFzVjFvzHHzuINepX64zDHEexyKKIjqxjcfztz6Pm0XAWIK
gCL1qiu/C4sl23Anju72b/vvizG+rYJa/8rt/PiLXZN08vv+i3+rK6ow21AjahQy
fMyGcDc99ORigeSqREPpDT0PDP8B4TjEf+h45uRxpkCLHxyX16LKpLukZ6Pn2aVr
M3TM0gaQDbmJj5NJzz11eA1zCXadTqD7mwwEmev3asvLV6TYfQk+H3My89glOKd/
s4pAmME5f4O+4w9JVyAsqnBKGXtnqlXlN/emH9NtWcgFKjuJs+bhnrq3biDBmqgO
9AEVbXa8cSEuPRDRmd9s0DKhi4P1PqPnCwV52k8hJRex5vGjibmNiIVRrTxcZwiX
pYZrwvIV0Qo45gUMRawAzLVYM/7EswfGyzj4FGo1zZMalWfZnuQnqvjMQVL7s7g9
CAJkW4LCsYFeDTFUaCnjxeHDxh161PpAdq+pM/vYdZAFQZiyQjJaI3IKRBzTVAbE
ZC72Jg6MzBG8DjBlqcKhiPVlJKErNoH7K0pRoRQsel4qaxJRpiZBRm+ZqSb84exn
XKCYZvHfeASD7XzHu/v1eCxxpEfFkJuxAjnAr7ZBRG/Gp+WJ92CAAK5uQfqHun3A
scZf3/z1sh6WPBKUiXt3ikgQvFtzitL9WVGrvN6c0laI7cride6nu21vYxSK78gZ
+JTh9bnP1iuGGZY1rtlGUegz6vhMWvXQrHqvu5hhDL/EqBWkgAcC/QouKNw5C6d4
U+PtoEyF22ur1vNVMS8yjulJBbnfEWEx/cBc4Ho7xkLKVBpyL3hHgx8Kr24yPe0i
jqwQqpHAwxezOQtRTxeCEOZoYB+nuHkbyUW0k81aDSLiZY1fjdOds1a6D1v6Iq1y
oybrSfaYRnbckjxAn6YdlkTiKCiOoczQMqQXGvP2qtCUkXXc68sfu9tevPKAWnjg
labelRfgsKqOFv/YzkH+/b/HhuS7OHlLaSOpUAaEvfrK34feym1CuHXxfHiK7lI8
uTIzpWeNnstIdWzSWrdILu/hMH8ubiPcoBOCFteL/wZQ1wzEp1co2MDVXB6SoXTX
AEVQILh1BA0KzdmXupiuokTfR3flR1/wvzOyqZ5rGpQNcRuEkfeF/PUL+qglfMim
irpqhXIzG1CZVNJOQsGScfTAXYyV1y4dawQjc/uA6akVFBCUOuqthgRSgyJviClU
uvEpZgDBBs9ABRUOemiZ1J+HSsxiMj3TSBvecDPzvpuxhGYPuDzmh4Cl9U5Li+Lh
VKyWAJ8enGeN5IlDpI6ITSPKPBb0YT7hx8OBOYo4uZLZOqc0Gp51qPgfl+X5pZqT
7hzUIv08lJGvmtMiXmIpNDjSdV/xU+fu0UrkrEfWGPgaoWNSmNn9/t7h5OZKS7A0
IsiSIkK9Ep3BNWeeXOBzx0v3PTMVRvDenHCDB+KBIEwUKnAzxkB5EPYxPE9CBajC
+7MDrMbP7g+Exg6H1+117KU1wKvtGEhbsafmXsf2niJOjHdNHQVUycK7wfdJtMF8
hFUouJ/W6E83RWg8KMQKD847APkHY1hIhwWbf744f6jYTVuZ65BTUup/Ltc6uQMD
r+jTL+p8tI20zAEPO+ex/J+StxQAEp9BZ26qfSN4utdyT/z7AJK9L5aJTh/9WgzQ
XEi4F5mAVKnzJem0QfrtorYVP45Y58io989hsfONYWIWeVARQ97089+dKo7w8JFA
99fNOlJ9ioUktdrr8xVyQBfRXvOi3FuC99A4q5wDQKt2exV14XBBjpJSQ2etRYo6
BCoZ0sOQ7k+QquVucOW7ArG2/VhVLisZf7SsMvC4ID78GdU45wNj8LPRJpS2iCsO
oWEy8hB2fAbP1xevIRresH+XWU5hNoTp63Eg8fiWcx3nMpoX1L2B24MS4/H7HM5U
bbfDFTnuwxeUWKcFaG01ToD51htbJlWH8kFn15CncBxBW5nkFK+I+pltAaZlujhe
BmTMjUuk5iKqf/e9F1MNuuO/fyxXgm9CquV16vE62Xt5qF9HXMEioHKJopnstI/L
tR3lJPJ5qnzDpn8RR21cal3cjR4j2aWePqDRSHO3LE+GqYKT8KVa+QHp08vjZRqQ
i4XZsBdXppn8+67NrLO9f4vIT9bCIwPiPUvTlE/YrFW0qk4fn68dQwUphr8qt5tp
bOz8V8oRjwDE3DFmAivIlfFlWycocR8EhcRSGIKbfu9hsxh7Lrjcp+t7NYwx9Ihm
mqv7MLMtlOX/W+MZbs8NaDRyG/SwfMsjy8FvEW0bbOTCEW50rds0tfgTN51kKoIH
W0D6LHLRk++4hfRUBF2cspOfAQw+8oARdWlmvzceq1ujYz3V1PzxYsg9QYC/UgnA
Y5Kxgx42nyaSWvQNAyTypzrranG7Rgk8P6a5pnRrgdTUuBN8ujzKgpnbX3kez8S1
FnCLTsC9H8GVK7J/uU4USD2D5qqnFa0oiGRZ7oFzEUE805a+X0kU3fMBZov+24gx
PUT2+4ZAq+rT8gYdFFk72CcQMliuXD7WTPcf4iolZxvaXnRcc5jOX8DlbMc5z90s
Qy3kj+bpkPxJxUvl6RyPaX9gO0wxYwddVMqsu2yq1W+1pFtKV0nRAyUOiqE7KCk/
/k8pTO5NmrF7y+pKdSDGL/9m/asuvB6vCBDJLf2zm3B3886lvvbm3V2dFde+YN82
5kPrKUwaF28yoGPpMVluY31dMeZSrHwK7NJ2wOR1X+rUlezUVN8Pz6vPBI+LMBzs
aiyecA2CuvU9Y0K8oO1GoMnQ65hyS3Qt2Cl5fNlqB1aMOWNLAJ7Xi3vWwxSLSPWr
u7cfF+yKERLlM2F2h30t6oKP1lv8a4Ds5ebKeACmHCuUxN5UOJIfbzJ93ctzktUA
YV9nXMi+lYmb4HpJrU/wOEcw0gkhZTixDytoLvrQPpjhFbDhYQOi+NdGj9ml0Nli
fLDoMYEnBuoYBsEKrEbtDXcb2wF6cYHHwLsU3WXh3xPrWXmzRbqxl6dFN5KH122l
dqZHdpvcIvTFj0b9nNVTifJYx6x3CEzABgWYTU/ZAy8NMTUq32mxNjs+H2ysJrku
ltqhaAmp7GvWnqG/VYzWlCP2udEOO4wupXHeeate5nO5k0H8CwkTV3gFksQ7bDBR
uRgq+9K7zYThbuqzzPOKk99Zg4alY9kN8eKaTqJPfx/S0AB7uR2DJnjem/KjmV3x
AnKHLLJ27XuoqU2YC3l3aQOVC5+4rG8izTyqNe5ocdQMoIMWvLEA1bd4VKUJu/L1
jlM698GEoV8uJHOS5DSiBl5rOgPunGtMhZJWnHTpryfMherQlJDY3vaXBnLqKg8S
ZrB9rlY7eX61Z9opKpHiYEftQ/aHp+aswHAEX/DCDGp5hQmBn1bUlcOCWUJdMT0d
gt6sK4u8a+0WERN0cYp7Qof1z+DdLkPPXktc56VjQdAdpEZE4VpxCR5IQzRXzGDo
aQPXLPgebD2D2wYU76nGLfFE2E1rfAz/qzCOQu6kr6ZEiiWAMDJVT+XiK7KEL0Iy
mEtg2cGPfSpf6uhalCWnzHuePLH8lK8P4q7Zc8ZQezD5UEg+n8m0kUeS3nCsY8PG
EMZK7Tolh9ckIeCA5OcmCIoQI5g3+c6X9dX5pQv/I0PlKe/rUNb2DIAxIDEXmTzd
KToFeMb+wfEgS9jH0bzpoBOISif9mdq6e1pbJ7oK15Gx6fPiZCd4rcC0aOHr4QfN
/I9PfnQ0qxOX6C3hl+lUqClvp6awjXpJO3duPuZ0mqHx2Dz2VLO+bkqurT/C7V23
IyxqYyohDWtqa/e+l3GMKS0uNcyTF7R2cEQPQae4spRH2tfqCHwG2AeNTLU6hAQP
MKcB8AVx9gMH/P/p/2VpsPO2ciffzW2FCb88wj8zONr1ZCr4Ou39C2Dn77jGXrfJ
1ANywz1WCctq98J8Q7eI2+517RZfYvq+PYXiHV2n88cCYb6hWHKZ3OLAHJ/LyGGF
U2HwyqqI/DXlDAlRlqC93X1P7XTOnCDpL9RolCxFBX5ToHU1drwQJShJ3W/AZcKa
b8FGLF1M0f06r2diLVY5byMkLxsknd9/WxXZBJSOS7HvU8bfKieKciVzv7FLamw2
TdFhbZYgpqZH0GyNiJr7wy6aG7Dng/RHYZZGCPRvomr2A2+zqz3uiBHfxNvFMlsb
avBy69skV63K/yocnCrAOr2k5LU++HhAAZmLJc6SYkGU0vqEIIqi43rkcrUGQoLt
QQNZ2bzfV/+BTnlEBBABG4vRQnfg9bSvUAYpZuju83vn20kTXpuMRqjWVuO0Ru+R
KXfvliZO3AwPImZP12fWyTZEJoHHWe0r4/LxOUBzPV9EbTyOtF9UgBTgwQ16zQcZ
G9I15zQnTFHJb+6rR0L5t2dlXsxnWE7fQ+RwddN+qVFR4UANNpieszV6H/+J+La3
OWjOgXz/v7ynzx0LJm2GEh7UmfOA2ZJcwkVA/mUNBUbtJNt+odBaP//7nHKZCVFK
y2fqlPuEYR5H8D8xhnGxetwnPvGe7PgvdGrKcswCedGDGNELeWWPrLsIe7E5zT5p
Z+PlCqn0Y8l2jwmCtK7zQd0BtMfwogW7PAkV/hzuOSDYKJ6vg8tl3lu6mnZSafcx
Iat9Exm9lesH+xrj2j1WTXYlciGO5tjTGn2rNhOZ5HuJQs1egec01yuaG5MSiYvC
nQ3EyOqaAF8zEeDsD9rCKmjPfuzwQ/GEZ3eRhYGuUgHxbc5KTT9EckF296WWJufn
hOliiXuOV1wZQXhpZNryoojb+jMS4MotraNjNOb0S4ebGo+rMi4ID1TNocrj9LHp
UfNRAeNsP8LvChoFR2spT/X1wbBT32GxBCUG4AOSwITQ3INugn2lpehLFiC8K8Bi
uSZW8CdHPSjAbLVgOtvkQKlD9Q83172JP3mwu85mr/m1PU4F9Qp5HZNldjvkgaAS
LRXakYRs2NZZWEwZPkQtni0biNrTOLY/lzKwvYVWd5o0PQECQ+VBAczhvgJASC5w
KUpYD/yloGn27fzqtItzXKfbXrJMWoD3bImUciO+NfHr0XG0F7zI2VSiQi4HkL5i
F4bUKqi3t63r0l1v9Yufacxh4G2KjJ92aUY7D5mr12FkQcFz6ROkMND8bbJiX0Cv
fID9KNdWOlkYfkDDz/3WGJ0BS7crzZQjTWFGrjWO79WYHjjf/jlGDsIlPE6+2ESk
XlntPiG3AfstQiRkdmA7PxakAnY8HjVbtDod3MOP1S+JHkd5uPCLwXaZfeKgFWcO
wu3wnLfFmOkWtLG6k1mZe/w6i3UP3YRMtOkMCn9jQHFtxedGICsleVKqKqdAEsUg
hKlPlyUH56XYPOXWg20DXJl6gJSE7/BNdAU31BgcC19PK1Whsv0RB/ywqpKQazka
nC/DjjHwOiEUdugRAXBAwQRbZxtB3Jv8c/2R+7IGa2vvRPmDKPn+TAncjfFqgl1n
zngfxHn89La/D8KX9IzNhWoM6jgg9uLHkeERNXTf3cCLPHCnfpazvuHfL7tZiwAN
wHm99F4tqefuPkczobBGuj0cYNm/QFbQX5Xg6/obOmPJhwyk27nBHbBFiBuoahk9
8p1gAHfD71Bv0ExqKiX53o6JhLnF0XZcCUq+IJsVAjpSnmxhZZdhbNHMLFrOaygz
xfAu2R8lnEz/9my4n1NudM0KdANucyWy78dqvQG1hUcfXJefVVDNofmrg++eUpgn
2/TGvosq3jbAJGR5K96jwB4pEy2tVW8yt9Bk4aXhRK0WTqygCp9RisQG1pzX8CO0
YyZADEbQFuu1iXv2Ef5SQl1AUUAjqfOssupi9qlnOE60QHub+rqCKJxNTb0uKyUQ
8PLhD4xp/eGBOQ/mi1GMZ3P7SKaj7PcaAziqcbSPH7DHRZ/iiw/HXA+CBlXHmA6v
9fwNYLelzgGTcWYIEcKeC2n8wTdqpWMP0ngXZLXUiV6fjJZFjHqS1UnHHu1tp5+X
dNoc4xBBUMwUxVdjZrOmolTbwQpW/4D9XKmWztEqMfzpHkrkfnBWfLcnKKKm/MiA
2dJP4VU1NN5zm+f6TBdg9DC9NZSIxE3lL/fqdqzX4ApMX3NYcsFkGfGrhHQy3dhu
Ij+DA9tSX9P5X1H8VUJFNyBygAhxfdzYOB1aUG2tofFj626avwHvJmuCbTrVb/X9
wnvl9J6PjiCQXKLuCxAxmy/L9fxmJ12YlB/Ra56A5Q9jtpJqutt2MSqVJigEsdZ+
HmuAy8Agc4tocT5ZjS6u4iDtAzG57Rh7Gj3+gOKQQmdnVQvRNxLKDrbrEqSOCgsZ
bDGza9qWtQXSysb4zC4cP11eBVXgIuvKouCsFmyG5agcmPEBD48CAgUAjZdRKOPF
v7HYOnS6nuWAQmt6M06evdK4qD3341wv8bgy82xp47CPpWch7kfe5TD3cchvqib1
N+EzV+74NUxzP9TghQCrHFomM5A77D3enKN2tSGTZVWU6PCu+aCgQ7hxwjG0gRRk
elUeiDrgBjh+BIndYpXZL0wOpfyKK4WBD3nOko/r42gsCvwN/ea/nVqDcf1t0EkH
f7zpdtkfPDtZIRgFBRvYj0JoW/p6o9o7YXk6cwJ3f9HeWr6D8y6B2BBFNWYCpL2X
8N12vAzZ0vEYY7dc2E5sC5ESAwIWGGxxNZy1Q+ywVuS3fY+KdhpeNhuG0veImvJO
kBgBUL7edCXUJZ8DtPD6LPb5v+W9YyhrB29XMkGpLc/u25mL8+RMYQicYug+zGdb
c3BLe8nrVNzwCbeZbEqRFJcfp2oMf6AcCprHwaIDtbPb1cDIk9BDBDiZDEsSYJzA
nHrPEK1Wf0+xPp/Dz+R/a3hwEcyp+wTMto4kOSiHf7YbJ8EvGVe446SWQj2SB2Q2
lyUe4ikmtJlSegcN2tdK+j97ZY/Bugcl+7JaYSj64mG9DbBDHPUJfPKdhwh/rpIo
V8dYLnM3kDoNtXhIkrhwc9Z7g7yFl6fOnZt5Ahi6+E4WPjtKTUwu0MMRdfrKV3DU
VnPEFOuOGnD64/fdV6CmgLOuaTju12HxlzQ+4ZwltZCCofa5DPadLbC0ZcD1PAVX
pQQ5nZetHBeBP8xFGyjPN8+SpCTlkARB8dwWRF8RtnE2oh+NR7aXSdL/+6oX9iTC
K4fNQQYHxovWjVtbwQTthAEm93Qy8Nka8HuJ67YFzs2cKytpYj7ifJ+isgkBEL1v
a7Jikb5k7aa7jQhFA5fhWGkJANU4fM6jyzpoiw/lzi+e6RnGHX46IGqXalPErYbw
4dRCWaEfhbc86WkpENTpdCDWRDQy9zP1IumoRA17sfuV2NOx9BoT4y5OIJA1TVjX
pQsKKhGp5aGCCkfuNM/vV7n7A3pkKGQaipPD0dN8Ycs2BVsztBUdBYv9ZX4GT0Uw
/HJZr3cpKZIyvCjrj6iCKgr0FlGxl5D4vIoVirjifdTpVovSIy/S4lrIhOljr5zx
/Bih3KZ9ivcRZc0182xYlmPcJOcaVu/9oXZf4FQRicf6XidDAWZacwDtTS9K5XcO
bqyyu7LramEbScO9ID6VQ+laZdl4R43RibA1vOePyp84hMplzaxAAsdQRQyqHr8C
pR0qlfbCQ/9Cc9hGwbFpmzOMzEswVX5/aa9HRXdECb/nwBOznRMjAQwUSvTsUG+d
7UwsmEa8WHfSToZ0bQrac14y2LnzJrHlBBq8ys1VREOVu4y7xPn92q3kjMF9fYp5
vqwzHNJvxBAvXZHZ0F91Y5D4Q31x6mQnIqfqB5tkqOfhpHdIHQzOJ22wdtTGoLrM
t54NqwoagS/LbIXySq8AYO4Nws/pXL+5bgI+jB8O51UaBcRsHVzvvH7h23CCb5+O
aTq7MM387WW6QvEVeyFb0A9+X9CrOnKj/OIKrQWYwDdUwTCFMnfQ7ACAlLjAHxjv
qYFmCT60wHDUC8xt0k/pBPHuwec+vrXmACSlox0wJFZ0t8ysLLckdlmXMZGBC7gE
ABZaZkFYyT7RA5KPlUqIo/IAjEjXULh4f7cThWGvIh4zqxrU5ExjMDUNbTZsKy6v
4uMlIvQipeqZ+bO5azIAgxZd/TEMD6Dl19k5CQp1+ioe+A2LTYDFyx7UuS2vg5nb
6qx/CTM7P8DKnc+xIQtU/A2WKwzhl0ef4hPtVfey7PLQ0L6BsjrGDeF1pH4nUDTS
LZSG8KAJzkmBvmopM7RHwFGxVBV68nUvecow6vcMCqKrbRTj1ETcKcuhJzN0S0xH
MZxIH4l/UuGruBIfR0Gq1zZq5JpknO89KIEf9XWc2Tw8iPcDDkiWlgiI3mtMJRMH
u8nCD2m9ieNG1z/tjiqEQvzDi79hIbBS1x5DR0QSytmOpJ9FnAqnB22v49M9ZFZH
8k+SDZ+Bc7Ch54ZtCIglv6I8SKIvgy3f1UwS4yJqent1oNWLt1avTkGcSX5gJdH2
HaCuJzpeNCs2TNeaKsHaekOrzWrm7zHoLUXlLtHR+ZNzjlFTD75x8Ybsl21QcelG
6v36yE3VruB5VQjTv78JfY1kERZgpShOEvzkjGdmb9i8MaAhljC63ezRTAp1/Wy6
5YxKaExCni17H949tNIqYSQMb/W359aHFsVjgGkDAEMojiNLsOwpqcQLyoGoaGRx
GtuaJ5mUpFZg1Z+Oa0vWWbVFUHew5HGjrKzV2hKC2rkYHNKJsgc3iAueQ0U7Jqdz
VLta01PATzplGc70ew3OSX3vUHut7edDgClfuzGVAfZw+/SIpZxrFhtBo1Ts+v7y
LwwGOsvWfBTA24sx2rCzlR2cBLui/c6wWZQbK0brXzSl1kqvhqQjRYgJ09nT22wL
9Xk5BaoVLe/+FqYA6ZjFGbSB/SJ+yjouMagj2Y+umd9g70Oj07MvsPDdskrqwrvH
ky3ndfuglfuX/+GXA0XHD8mxFAHA5mS46FsE95EOGVLQyofwWblr0l9LdNQAeMxt
iJX0QXNtkqj+7s3phBN0phlgRIr2ZgpHUI3nnWPSLDvkIdyQ0Fo++mQJo4DstdIq
YLeqED3Wl8AbgTRaSWHpeAoqxDXmvs+clLq5SU2Xgy8U/WgG+DSG48fBvgY/Amhz
udFneCc/BrGxN1eh6YE4XqI+Ij3TLMwSi5JmX/utsOq4UW5W5WQ6Z4O2hwoXpJ5b
9HNkqxyC5x/dpfUL36Mr+6TWRyoAypMw1fA1A9i1kwE8/gjwAlQb+jkf0ILki74Y
Bdntindfdj0hAAc8uuwj26/oagCwtivnWDsw7BdnbNR0DGFOjNV1CNfhQ+dtbESj
RFnhxJzluRiT2Ricbdhh63uiscPEy8Zn0tWKb5yvhdJA8DJHB5lhuKKmXQ3Wbxq9
bqEWfB9fnFc3FRWEj7Gy4BdNJmzZWoPKrK07D+qAAv7aAFqS/OYnfYyqGwmZWy7a
vONkrnxjpXrkJMfluI6EGe7GEBAMmyXyHR4p1mgtOpRpip1GKZ+/ahnz6EeDe4/l
6hedR4cN3qQBxyEd5MFLM38DzzcuBbdUcHhUZ/uqShr2/20xY7+XhhsQqLlkV7VY
CRW6ZhR0i8mlfu5ZmUCtRTLhVVC/uo+ImX3426h2VD+AFAqJEVUAIQh2RIoYc1Aq
3803IziLxMgBW0kiKH6aqdcishdI9d8kP5ub+ftNW4Zk0vo3dnmd8ak1SpEC1l4U
PWG6DfkUkbGsP06+aOlMN13Jo5ls8dpmZ6acBusPLbJ27h6GpcWGnldN1EoI1Qpo
Sj3U5TdHbP4tX4C3zSgmvr/XO0nQ7kMC+ZbRPo+fQrAW6oT5x1LHx9sIGtbeztN3
awXRkII1q4svso3sGQ0bKzqmPc1Cz754rQP1GbVkOdybWeJW/2aiTxolzJZok6ew
zcOoiJSZcxVZSjZQ8tU6wTRqRhZiUKlsu1VnF2GgAyZiYOSJ3FmtJNx+1J+K+YSG
Rnl1Xy6eMntbnwvsl323HPh57arZAeY2AC84UjcWYizi2ONLstdt0/dxYke6iZgs
YA8BYVQGG6j07NhNNa0H/scmLGqo8SzA2EtUAWNGKJeTPku/hPLqUJDFkantUBrI
JxTeDBE/jhJT6mjOc/lJ6ofLZ1OM5qpJ2lZyYGvQ0yYfIX66/kO76ZG2AveljAFZ
bI0YcFb1XsOfj1+0a+Fd5mUMxm1aygxQpJX7pu6DGvE/KTj7xDi+34WmNBQ8NK9l
dKF55FZCAdKwSBDs4ADRlvmkEpgMiORAxIfId7CH7WNeMnfNeprUH8P4XPB3kLe9
JixNru0yksXvWIgNf+qoP2B1AT8cAmL/WxhCUAMPtZBlth6w0/Ls3Z8S2ZTEndvP
5OzJDa3i25pOFTohssxeFu7JAQs+VY3sMZHrl4bSVD5ahftru20N/Ornlh9Ewgcf
QVIAf8p+2S3AODyqiixfRgtRzoxMuGwS8J7/gAk7IMju5Y6krOjZaufr85WvrKCL
M0vDkTefbVRGPwxYP2Wki+CgCkE1w3jWXBLRiZFtE7y19HdIj6lfhsrWtYD/GI0n
qris2hpwEFFiJhrbrWJ6iMITjaZDaw+LzS+zTLrze1+/8e0uhaSH5nReJsjZFwCb
uqgI1dyo9os9Q7rDGdc3oAEATyIMuBNH4uDZZr4KrvZytVhbJiHmd95p+zLIo2oy
XnPDPnJkCrmG6qYfBImAZaLQi+NjkoKWiaJ9MzHSpMRdQWmtNz/IinBrLGoNw5Ur
7CE8K9F7QFREk5ltLLwE7V/8UA1Kn/9oXvGFDNXUPyVZwrnB1rDEnZtVHN+n6zQC
A/q7zT85xn5wxBGo3Ht0khgp8XwHG7CX4i7exeFRREQg82/dj3LtuPeoqpibWGdq
RT0IUi06Y9GNArbBZ3aLBGkTDuWTtzSE/26qAnd48U5hy0bIZ4bcY6dphMbFYtok
DOA/dM+NQs+tdOkJSmbYFBSqy5457pBB7ws/BTBg7xHoZFWeD12WNecNhaRsu8Vc
sycdSbOG//thBwcsD4ikfzzW4utGvKRlafrZyE6W9SBUHuvT8F+9P0YsVq+o/LNC
Oob2X2PpZl+sLKjuZF0cOUTisxK1KzL/7zoaqLpshr404uAV2fMPUuKXcBVe5n2Z
gTH5bvchynyE6J7z0IJHc7vgjzr/g80jUUsJIooAFw3HxfjOrO7W3rsdOOaCPpZ9
obPA7A2q0s9y+BU0ErWtXqA+BpixI0R2hevxQX3dy6fIko5lPCN33xiIzFqvmTrE
n6XgTy4gL3L8zuVGLk1+sjEC6ddPqxOymi9fGsuSk75kXJePGHLBZSM95kuPZ2Um
PRxhqIVmuxpY+KXE0N39k82/LDlZ1YFqYaTEbrArFjRHtcerlf4ZxMljwp8Ro0tR
+Cmf9R9snFLPtvOVF9NbcMbmxTEk3E+6T7erRyqGrajGl+duvlCi28Zb7H8lwQNS
5C9Fam0MUCYZ+0Gzs8Dzxxxh5ElcM6if1VgFJ0gWJEitI7SdaLopMVtciK0TVCKP
B24PDM895Lqw0ca/K6Ybv6zQd9ij9KWIpMQYdpafGhsO5H///1JJCA2/caIqBs03
3pJkvOZj6aXFMCpbI4aYEQMbqAxAe4zhSnU2sRgKfCZIKW9gmwW/qLA0yM3GQ0Gd
n+hsQtGlaP4wbOvJDtoWUybTQYFWE+F3Ui2Yy2BOu0j20ABzO5Ri137E0l8C/UXp
iMHG+zDS934b7+zRR1sYCSc3D+UKBXUJHp01jnjFSrNzj65vs/i/9AIVCWTklR0l
T/685v+p+yvn3Zul8l4Gmsg5V1wq/o/KmY/5lUewjFsS6eGchf4Ypa7HuNmWb/KN
AALwNKdj2PK3TvaCpzVcpi4besKXkUIYtxtZ+f2zkeofQGyumsQz8BaX305XfBNU
EDDdaiLTFuxoOdRKtVkm3hnekdZASrRrAAk8HMi7c3FXHX4iTcAli/i5dExR7ZtJ
Q6yjpvkXO681BDd+kvoEJBpANHRPjEPIXKn5PEny79jhoQL/n70NZ+01K47Y0zft
LBUO3cy9HL29hkoR+DSiP5k6Uo/u3E82vlV4b14BH1ksRdk6hVW0R1hugOw0+8iQ
JjQtP6rAKcSsiwLJk6h3IBo1mgFm3ma40IvOE9/dCk/vC8dwuLkQtsSaUVHHyXFM
TccsgVSPqk/41VWw2EXEoFaNwFSQ0C4Yd6BCRzmh1YUSrEzTRqaOEaHD5FaOEElr
IUCxd18FBS08O+swQWvo4aqYFaIpI2hhilpcDhNyM8MhTaCOAn50oQYYKpQ2cjLA
IgFwCUqvJtPhIHTK1Ne/qbDnNHSVJHcjUUBrErwm4WKOjooB9knBOAsz4gM2tPRn
ODEFf8NXIxOSSSV21dm0udqr9q86yjJFo2aCTDG5hxuXQadwyJnaWU+GCFluR9Ux
h55NnZ1IB+aJ6Qk5QYZcErAo6pRE4DXcRo2icS7jlz3CDcC3drhzTwUeuFt3cxOT
9Oyyodq1TooiPlGzx9p+0YvmFgPxffUScl2b6H77Xmo6iJqkZDL9scSHwKap1BA5
Iv6pHJbs8r7GG6P9p2m9jDhglg81PTviTcGgqKDNV8s6O39Fr3+/a4l6nwV+Jdfq
MG0ZhPBku2SdpLd4mi9uz4qioqOwaUQx41G6XfGwtXWLB3ucYAZxf0DxpHxmbrJs
7W5mIPyBo/hX6Nf4lnyg3QfnqSHU/byQ3bGboGt4T7qmUv3q6UuMceEHwCJAPDCq
qDgfim+ULk/51DscxtKFqx8FJGbT5FNmC1cZXauy7hVFtdHYWv1Ae1A+i+7vCfkX
W0WcQJw8TDAr4Q6uuUUtLf8nqiSFJlPIH2lJrr8cERDEj3rHxOTfM3BNU0+jZfrv
F/995wgX4PjLDwcFScGjOLbAiFYjDG/sJtKBFOTKPJpsnNoA+3frTVqHZ3OzjXKb
Gn6RuNDRJavIG7vhH/pekuTyX+agzGzkn9LOv1qtJTR6Z2AkRi9mgD147/Z5eEcW
stG9HLSPsFl5zwrVQKBWyao3fxWOdZYwHqfrtB4jenyAt+FebeCL+ESIQ/4hLb8F
Kb5GFRZLc+tuNaL7VmWxu2pAUwHo5YLLRM6T//zbrLe+YSAGrbLudZqams1R63cx
AMuJyhYm8mQm8zKoQIlry2lQLln6JS0IPJwKsZfK1PnLFcTybdV+8rmoZWifhz6Z
qKPDITBgZ1Dbhz2/XPZs7BaaI9EsbceVrq9IH/ufPe+GfZrPRlFJsU0XwmNv6Kzb
PxbpmkvRx7uPYwbO2xb9aCoNkoz39sZpgHeTbJOd8yjLFMpzLtJiCXQQNSPlKF8a
Wh+MQJkmw/ckxBFaEoB8qzCVoI1bJQRG9YibcquKveBLSJdjbVjiWuZ2/UXPtUF8
ypI5tUrZuK9++fb9aCd1Xj9jalHmxU+IQhGVMh6tcc1Slgx8uEU7BhQWumPvZVss
PmH0aUXZiJO8jlJXgci3uWSDE6/WvnXV+iqsK6Wkqz6arMj+bQhlOE7WfM01zors
hTZG/XXooqfHL8lgyhWN9psW1tu7xB452Zac0B7Mm4YD6RjhwRBnOLEjhoQlEF+e
PyFTfQnCkjb/BXnDOk9G4omIfuw33NxUdqf05yBgvsVguLWR5SS8SB9X+1TcX+Ut
YCBlnlciDqRfPbWCY7WQy12rs8npoNmfVqLDDysBqWtox/M7CNQR9Qm3dqmhsXZV
S3EM7uy6muhg4HnLwYN2UUctu3195eagzUN3Wm6cNVusY+pXJTLMBLuJnU9Khn2u
kuOp1sHjVypWVi2cXItgzasR9yvQGFrbkt6vwcgvlN5NRdmfeRF/6K8+crAyDS6b
2NWqoj2TJtRmfCjsI5hEfaEBjzpezn2R3iOs8IxmtZJ93wCoPXPUiiHGlSF4hsIY
OneoGlwpqp55D7l+tEo/RsoEiTdsrZRETEt1JNXwX+AthYFVOa4FXFdVeSINnIVH
eyW3hTHg0+iOSWDXk41EMIlcnyn0vy57SncjBXopHwZOKKY0Gutc80zN6imy7/Do
+15DcQ1f3wK68B6iwgEmeVQbtYWfUyopFB27L1GFfORu4fKT+4y4LRGBOjeuq5bU
N9zmmUh0LXQ8ksdZQYipYTMzNK/Sv3HYmnBEkRRmFHYU9CubdGNjQCU+gQ2F6swf
fMvuw2UgsHN2ht4XKN4sLcgWAFeALR9lne9aA4Kapp++HflVpyWcmY0HO2W5SJBW
DVUkuZiSEqDUimka5H/1naNm/mL13/vU5FGU62OYMKQdvHmICmc+JcS/hLGM+X2h
S0Ofe7AvYcD7hwDQlJA9bhJihO+aWyqD13U8W+IzdU+Eg6BmJ7g0D2u/aWb7lCbc
w5QJOj9QoKNzCJPpOjVP+5sQGFnmIL7I0oibHNQ4iLu9EpmL3zf4bnlzJYqNsRTD
ij9YxZb+7tbqmDH+6Q5R/x5i1uGzwYycv660h9ei/o12t5fyV5KOPK2XptLuxWtB
3G1FewUktgbg6f7d7zGeccoe2AM4vy38NX6mTQKcZA5hR0/vH/Ia0sUd133Tl5vo
iB5klkLVWFzn7AzBlafc+o9sbiStJpBsb+yDRATab5gvgGRJtAANSgiQSk9Wsq/a
6glvfbIqWdYpY85Ndtk6YlZ52EdGwPJXt4qsWamaSNwszxKSUEMj+oUT5c+ojYBz
tyTo5deSrBHP/AgiZrWwJP7Y3UdInhCF3ycmw6FZ9tLb/THbyEu5vndXs3n+Tjyf
oAeLQIU4mpxVxAsYazkK0FOI7kqAGYrPKAAWr15P+B2jWubXrqQqhfWtinX7gg42
RnKRCs9TJpCWiuS+JABeHa6HeuRTwnI0FkC5JWNYpgf5+V5JKywg660P1wZ1xEp6
fyE07GVCgrtHIxGEGdt4FPxX9ENI7RCfrKDbXYnqCIQH1iUYhldm0ZhpWtmiyaDJ
xxvqh6xTjKORLKbfuECwPZ3uohc0tfxt2gWxmfcqB0DGAW0U27s1wuGneHeqYQRr
0NOsPWUd40vleIQbNQKFPFBJDTEFeBbxxYleBxgryJcelCPtW1qFnC+6GOQc7r/W
ZP5XITrdx2rUMEKUq4FKyiRDFXJ96v0GZtPN/zrlivLaNXJ2tKWo2lS/OwrhyMQ9
oDmtf+ItVPrODhVbXMSBF1YmG/IRLLm2RzM8ycdO5H09cWqAUVqnF8WLZDZRtlLO
0ukwNoHTxEgs3CbQi+rJDaBieX5iyC+20jxkCz7BFKEKL1S5iqs+h8ESHF35QFeM
chNeBeDJD3X798XZU3fV4qyW8rjxxFBKlMj21VbtpWpDVYIoqqs3ZZWs4DE+uKOm
qgun4p16w0LiMiqwJhH8D2l/XFdD1lRJZoSpKWRx0NVIVFpqwNDphoxrg+TLR98l
irUpoDRECWqdNbVNiys7uejEOHcREFsDWrT7Ap+jzyKEuGMD38iYDEhrPY+4LNvT
CiKX7lrdPkbx8umuIuP3CHke4+KE0Tbsr3I6+Oc9Ts6clSKEkdtpN6Fhy2nnLnCV
ihDykQtHW4/3pvWy955xdpyUHgqx6Ch4j2jknyAfFhzFuWm72Q3yXWmqD003ajQb
nHI+6dM+nXheVNwwkBcW45JnZ76yEz4NkvDDQL/LCghRp6nH+GBIWPEkkjau9Xaz
oQB4Wm6fwemakkFnhZWSgvkSLH0axTadEYLZTpLy42fxQ7ZMGCrkqtq91mhq41Yp
w6MLgRPQQreaD+Klhx+pfpQIlvk5NeXPoNouuyuhvOY7kCMMJLtYGIRhZX5tW9Qh
2QFGaL0RfLZ2AVA6qGa4enAxoYHl6XH7zn1tSDRv1bsmouTM5CXNAyo/k+90cSVb
DniO/hf8rmvc0cNI3KEdmSQeZ+JrqIMCzVjJW34B+qkDd89P0umBambEAfIMNaU+
MmK5QpfEAx8kb7VXVFYOZXN5TgdDHcFeA3B0+bCBOpmUMuzXDZ7rphs/19OKbzOh
VfCOi2K2S67WpyNvI1VLJO4PcIBywnO7eJxtmRvxuyyhvn/a23Otppji8uIOCr2e
gNGvzG/O2om+0uN1TvjE4wWXLtHVj/KR0ayRPmyrreyXT4JECD5DldWC0fS8IvYX
GWqCXFwFrKSNEZUO3hYYWgb9XBCJjN8LJeFNh1/Vg+f9GAZOr6hWG8k62GBylPaV
6ivkmPa0hs02NGs/kuaj4Z4cAi2ml53EmLTukTMgA2oN/fkAgw9i2ZE3sUcOLeyD
3Z3HUD/OC4gfNrYNk/ng0ExO5VMwFm6m0BeugfbpuoQniC5/PmZTV1fCT/PfCsaY
2QSSNXK28P4p5RNhAtvvzGL7fQSdQLNKLkt7dGqJGLUDJPo534tHOcGDoQi5eVGr
cE0b1H6VjL4Idq2Z8ZrDEoblMpXHzwOsIxUUJHhGmv42rfA+w8D+mRbOLWK3Mr0Y
Uf3URyKF1DGijNFy8Wcet6aUDjyu3H6yzEaDTTxJp68sufreuesG00+lWdUHEdF2
o7PPjGzjN4QREI0DFKaRN/sLPcSA/iECnbo0C8hTsl8wlsV/UQLrs+35gEmqX5aY
lxRDltpHqgthbInnmt2fyo/T4XiXGNaGMjb/Qowv3xJr/Fl1GBOMq5vW9otEX23l
Ta2O+9K7ljFYnC1DYZjRnx5U0vzrQd9rP5kQZw6ivd6ZofMI5SoqCwHENezIikje
/mvZaSc2p9Hrl7cSwCGkHh+gy764jUTp5zj4/AHSPUbt/4+HkWytE1KFWo988DkF
26mo1nuaiSxF3nEVEqSYZHVvtd5CKml9KW9CiwNzuWO3ufQLEZQBnsNCaJ6ARsZT
tt9thJaJWZyXUx3FP/tjpPO92uMK+Nh2thVzYN0uQYbv0STEH406j1a+SB1DqyR9
2sHUaHFjXNVO3w/BUV4olehFJ3MOxG0MPeUiEZ5jK+T6n7InjSuFUV3l/uvIwx69
LP6xttP6+uCIouoxbMcGzKQPXH7QC/ooBbjgN2fDWVWf9da9oDG6tzhqlXcrGDvh
p4y7dp3QjVSPeHf6zmv82h5tJk29orkr69Jq1ZyueJb/EUESHDmOQzVZqPZTRHr/
T6BvAUmLC0hYZspkknZ1lkU9Ps42aETCeb8YFJE8yrGLPQKDXMtqAvlc0VGAGODb
P1lKqAUWpLVrWuQhFcCZvgWkH3oVbGscCdiYPtdXWbN0OzRepFxV1buisRYRq9OW
+SSPHSkAdhFNlgpyJbmCoRKEC5c/sAolxakILu9dVE4n/JR4az8k4T59bAlG9gKD
89ieqXNkHVyGpr8hz+ULGvDVBd4UZ1LnodCCxsJp7uBL5hHK+rUeeXHOs5khvWaQ
Bv7RhFFcvtnTiTsUKiQ1hBPXsnwMwXt1AsBjtAdJbZ0rD3S7nCrSBflSxyA1w+kg
Ryd7yTSW6kke+N2upzt9NegtYOQWKOUOZgZqn1EoHYYuY0KlgMQ4iIP9DG6l3ryM
ThEZ1qZWtY/U8V5OkWVmUTV34Rg9s8VIes4u6htct0JTsJn4zWkED282xrRkUk2q
hnobelIdObYSMdreckpRD2TpYm/92BhMCuFDjOAmezUZEigKBPt+YnF0MTjR6JMr
j/C4ABKrgAWfwwytuCr1CQ9U7tlw/JImRC4En2aZeH4t3FaY/UZBXDZH2oCD7r2N
GPNmOVzxLFsrOg9eg+Zw4q36WA39Hg/lc+KIeHDuCDVS9Xg8SC28056xMZVJg9GB
gJs1UZVYgvrh8T3SyND9ATQHL3Fd56/bKASke7OQcmGBiukYnaKTsQqgp9aiZnsV
TLSIKdCSa1UbPCvq1CDrmaM8xUV+LZciabrf6h9oZTgRItQnNRg72HPL3zrCkbxd
slZFCjDHAB2L79RBZn77ITUWsxhh3VHnK8uX2E9ugS60emdL9fFItsehmZwPPoeV
FZqFUZzbaFyHqWjMdYIcQud9QO3b4CY4A2wXJqU18OkMkLWq8WqyBh56OD9TQR1G
tiBvp/xEsjPQxFl5QzhQke1uc59dfbfza0dZQCXFP247S94ivkF1PaG+jb1XJVJG
xee17eDsIXGdEbBjEoDWts5PEH7DK+wY1kSwBGGXtLjiBAvTlzxGOqCm+moVF9ZI
w5jDHvnkjtCiYvZyUBGb8K/IcTHailLI+7owZggTo4rCFEKQziaH8ymGy+Py9Rtv
taDYFMtoUS+kc4PmXYfjoyQlZr5hSwRKFZlTUle0CFC1Wgtr2tttel2RoUxwk75b
43QMv1xx8j/392JsAZLoEZp+rxHr9MfeZXHT/KziSG91/zSKCYReNxEzJdl7EqIY
nWfE3PiEgbTQrtyh1higs8GIDXpsa6aKNxtOQED7uIUmTs5no0Mnjw54janIi+o4
cjkYVloRTLyczFtvUKTCdP/KMRKs/vY2V/V8uQZSpsxsewWKB/xaAqNDZqHWQ/NM
xXUtBDPGbbjWMpQeqnokWT2c9VAovY/tUjiZAbUfVQzlfUeS/a1FiKloMHuLFuk9
bBMFMaYMo10HXQ29o5YMVorw/OL0MDr/iskeZ0zIUuuR81l6QOHIW3xOUHNoZvOb
OVJrHZ1aepwUVz0g5WqChlX/nfO91taMbrGKf0kLmBrcZuGavdgk/qej57gc7B2G
mehuApPvddJv/Nu8a/K0IHc5YpcROmCFRGX5r2Aejgrjwls5EvYKEL84xjihXvXp
ka0+bdLcBSLLpLKE4W/Jb9fZp6cTBL1KpHZZDxKJSQschQyrWpU7YFbzzxOorK1j
AWG4rgRrczLpeKfcpvaQlHyN0F56inpeVRdmApmpXX+jPhzWRDjO21ogYVPouN/K
/Rp6rHgrnaQ2d14Gq/LUsG6wRff/em9jaRox//QpIeLFx/rM1QGY5Boi1oZZ3HJf
8UmybQZfn8nc0dX9uDN0v6C9y4kjaaPsykaV5WGqPbB4d3vTwuYj10qnYgkXEkIs
mDGvBVLzaqWOO7ZWKhf5Ajqod46wRYVUaRUzYPvNC/yLoXtBb5tGl/y0hdCXp8DJ
zc+NAs6VwnPJySBf2ldzlYPdTgeaLPXc3hUrAa8ilJvpXh2s2wN4B0fJjHdclN+s
YEdzifCn/vDiNuz/vtLOcw4Tyy+SNuZ0kGrO0+TCIqSTHMsTDWrFEM7udiYOtreV
o8ECDtMdqz+q0lDJ+TlEAGTCfaMaWx9/ypzf2isET7sSoCnjCJVoQv/pEPRxxBOs
qntNjnZlz+TCEZjJFQSbpHKHP0mBhkeOKjYup1e+z8HBjHRKr8I72yhq7ipbBhNj
JCahJHcvFqvEyKI3ov75G55fHIthC7KdnogzYThZoQ/HEyTugaNCJ1a1atnEsC43
84IA+w2gCvPRk95AfjtazVdD8Y65a0lQoLydGZKCWp/qtR4BFyOZ9UCawcKsPxsh
x0PwRn8ZvzEFwoYlzpdMaTTU3E2+oV2nSsadA1hXt+KIzqmq2ybUYeHJEBYr31ZF
0e53uR3KgqrxJa6mw8k7bbW7GUPvsMQtYs/y3w2QEiXvvVox3RDjegwpwCqAKu+w
/Io80wFf8DxhoceqzMiBt4Nptkcbg74y5crHnHoWETYHFzJcmwM2Y1r0/Vx+zMt7
svbgoqZl9zyh4qsxMZW7ZFI+I29D0f+dQ2AF8qGaXBO16Uxkj5SXrxlo7SEEuybi
BKaWEC9AMZ7f65eJdQ4DI8xVG3RSoQmATiEWyZVP6WyzydI3xRPe/eaDXDYdRHka
kWEuSMmbeenk7O+inPhK2oTMFpgSgaWjWUfmhP5w7y50EgU+9E89KXEWQ27KcahN
bjfiFkifLa+Pgqf9BcBCaPaaRdpOrz0PghTJwU536ygt1lb16HeKOeuSBdUUbTla
Mh9Or5OED5HCwrfXbpFX+Jko/idFh4wkithCjOp4qNYVkl7EyP3n3djhZp7ItyEJ
xh1cAaeJXvQzL/+BTGFnUdnw2Gk+LHi9MTs12+P5xQbcMW36/lXaj6OwoEvsKJLt
aN9DTLLgkbbXFXv9lVYiNmOC0m+7UTKAmdQUgjl43n+tfsC6AWmqMIQHkrE0MkiT
ktmpnRO0Z21YFVDyLOuj+jC+QfPFyYXvERxjIbIfHekDdKw/82CCCWi1Ta0TkZ48
TmOgw2sZoAy+HjlOuYg7nV5y8VVHKya1g8I4I9GSB93BtrVqLl/E/i/+/qnTwZ95
hP3kvnqWhiZpym5loQNHuAxLfFjx6rFWUEWrmZKZbvKtjWuvzjFiCK50wx/upNKC
+8L2wDZa4TMQ9aFzkuryeowvPZpMI7amXuoXjVi51cTtSyEflfMsxZuIMTgyiexw
ZVID2VxU6Jdg/amVPcjR+A9t5WPbKkKH9BF1LUwUVQDyVzcMp7ptBsXFYo6+k1g5
ZrhY+npJl/FnpEA/D4jM7R5wKRD6KW2XKhFs0iUrhkFvhBZeBZUMHzyrKB9RN4md
yXU4ro0jEOhybq3FGQnGEmSqtdTaHUZO8Pi3azU0n6kchUmuDj+UsAubjKZBJCvR
CPL4KIxJMbp9F+k+Y/YfUayCcm/y9V8PZk/YNodl9pVQj/IM1URwkOVbAtefRxje
e75hQZhm1B1D2WAYCcvcHKAeQh4JzRgkCdrNflZTRHC+viwVIledh68Y8Kd22XD8
fdmMAbUKWEkx8KUknSHS0UgbiBuis4tc+zTmCMC1F+NnNdx5WZkUs+MSXKj5+Cu8
5sPp3fgGTQ1LJX7VjEH2aAdwlWx/00NivTVeyb8iG4Z1B04mL0GDZaoEfIjaUhqR
uIIh3sMaZUuk86EOL0WMq39Jxm2uek7EF+5nhMG/0iZ+28+/Nhx6nEXIMCI6gIZJ
VvP6CjohxKVVcuqijyrKMkcvDfcsISZ08dC1RTbffCmnYf7OWo6DwLfS6//glEe+
z1jL4MPFjsDXbILOMKMYAxQRXDW7wFptD+MdS4rZysHD4YFzHZBCrcB+2bL6x3aU
tMvjPVxOhUyCr+QKa0IBQm+OouEb9jw3fduQAPFVmXmaLo1muk8Wh2iRMFjbjijH
BTkNFKoT3JF5g9qb/6vCG4SyWv6BtllkujulKGrJ4H+XIK/CikWkjItyeY+mxbwg
m0hqdOavth410+ZOcBiOMT4nU9CcYB4Nnm0fGvr3fHMAmqLzOdoCTLxvzlQg8Rvj
RRHZjGhLBsuv5Bd2Y9zJ1gAIawS57Wr0RvalYJNoFrSS8JbP++27ByaaWxCrjvYT
9JG7hWcWjqNMC656eShTNMf2c2xtmCorgqDzI4ef0gYe6jNhHy0w00pgUDMgyPfm
N9zJEXyG7LeugK21lISbVD/g4A8HHJhEcx0QX2kpRK4ugAdVESET1qymlhL8Qf+Q
VyJE0BxKw2ncjuE7nhWXpP7SxqeRcZL/DJJnnFJh48tcdjHJL5k7jEpQDK0IKaOe
eqik6vsII6mnP0phMN4lY1LIy3L1yJ9tJ1AAhIQ+ZhvCMv9YJDc7EAsQaFDYEzCV
UOdwpI8aB/gjg0Uhwyhg77hw6BW+C38VJAH5H68YtdvnP3hPQuhcZnyF/Zzy7Ald
db8XPAgDGaTNedvIqGUpk0wt8aqtj+U1VZwos0fG4k1DbUuXpfT7B80F+0X9uvFW
MfyVrjjhmZYDecLb1LZUB6VGZXzqmX9uWvicrpsukEwSWzmj0Oxaxh8XkJb2Q1w5
N+w43bOgT9IHK6nW8EAbjkvmlrE1Zd+i/gJpIFQRMCSSdpyfF8S3GGcgcRIeujce
VAD8n2IEbBkdYKatz7D+EwwpwcwG2J4ZurkBtr89nkaR7r6lbRw3Io51D3aHxKyH
Bri75fooJrjw/YJTFdERmNbIs68/OcyFxmz4ibzqLbwKwihEWP+wpZce6plSD8BF
ZtI0OlYeGluLX+Jog1qhb2sqDmGvLI+G1/MCOeK/JmaxMVhBwiivS3FOsvjoNY+B
Q0xp6Y1UyTi4Po9l3I8qGr8RBOFz8o1pwTlooiadj/Macc1IQ1kgHcDJ/I604Xtl
OaIkwA3hNnALLI02Ir2/7G4c/DnZo8JNSmIRrdZ6aOQZ9f5CXpEoGp8Mn779R8Dt
wXihI60+NhE6y7+aoKdnlW0Pn79Bj+4NbbrfT1ufg5To28OT1xI6N6wQHH30zB53
y9O4kuTWkJnQ5631qVeJ3fotUKAPDSq+Erti6xtTLR6G37iXmZKQn4lQjcLIdFHn
PLTRQYHStf1OQws7mLZYbaJPTVaPIR7OlXanXbTq+fYX61mln9IR0X+oP1dztSGY
2FTrgAp6i7wq/IDMe2TiicqlRyPr4bFSd5H7yCLFU/cdnbTfuqrpaQWgiyoyJpan
BmcLE+VziGBZlmZtiN0Rl3jOh9ZFTKYvfKktULnzY5/clnBm8GccsRjpGgWTHNdk
u1ZXmQMP54cQ8XlWpG9rDtHeSm8GqrtpKYN8PvhsDlMicsfaVV7BkKh9mf6m/W4E
DNkl5hQOXUt196fwSaPK1Gw6zkz9OGGvXag602bP32ZtLmwrjzAWa4GyzB3cqFvO
NZ92Gc3DgPVwgtKHZaydmdWyE/JICPUzl+lYDBuwt5F97M6MqmzzL7FPr8nSDvso
G0Hg44OtchlhivjVqHRPwg70EedOx/k6TahlJakPjjP/JxnLvPkhU/s5lhnwpdfC
m+d+rJJ5Oj8KopMVZ5Z62pnUV2QDRm02dIpJG9ZzqaHedBamxApJIj+UbsSG6pZ4
QL5WAdBOaSv7Y60vtjkfJXDHGjiffWOh/t4T/sEn5cGhE+Tl6yM13Pe8GXZoXQd7
FdshYBAKjXv6IYlvWZMEePPMgOR16cIZYyNLraRRxe3osZmvuf2j3jvdbjI55/sO
cuFdWPeztmmlrYd0ewU72UYytl6IMxBujWjHqGdvu6plELxKY0Bx4KAhSUoLLI/N
fwSiN2WGlf0PbEDsuGgmDXyTv+D0QY84+4KElRnfOA0M3XpudH6DbignZ8OYFVK2
owjq5YJZdFnJokHsFP6WVJjrp38F4mM8e7bhYwKey6/zJl7wFPS6hLDufNf7Seb2
epJeygaDj6Ad7s9KzeJ2nFOgxFV2OK2ooIEnHRBlcGXuMLJ0cfvTywPxNVPpkgqe
coV+KClknwEXIi92Hp3zNOMDwkZwf76QCjrC2Os4Tw9txoSHpZRg7n9D/1AZ9LCO
C4AUOutQlzBd6Pf7IrOUiPW6M1a+lHAQwNdyls/wxG7TTemRJ1kdYhhMyrB9jqv7
xMM2lGGE9hPttFGDQJIIOJtTZKDWRdAr1CtjnILw+zZt8UV7TSVe3jvoEqZgFPzr
R27tmtD8OIqMZ6r+iZBLWDFWDHDnkkgK3hJ4rFyuLMPSJbWk5VHNURwu7femD0xC
e8cCWTAaCzJT8badYDqxUAGhWTG1RG0caAaogIlw+Mk2DNo43WgkFkvsPdDsrYrQ
ymGqsuFSoEFkBD6Fp1jNVGl+x1kwlP35q8dGzI2iILF4cDRIiNP08izyLvpGRfxd
QYgW0SVdu9WBA3pU0dqmXMDMu2vlxAEtUbMcjzkOSqCu4A40GQjUs8saiTgAVD3/
EpRJOgQYf1SUUP2K+d31e8B6J1Xgaca0GpXdD5XSxzyUkjUJP8auu1supITIn+ak
4oTVrrtH++jzJn60DTtuk5o9fIQu2ZeUAYOW2yKEdt45TDxj7wiwjX8dk96ial+s
+O3C02wlJ5sf7IPJi5PaDK2iNhd8HfD0E9auclZES/PHzTMMi2ZO56HA/xzEptVM
YVVoUrZXACbLbnv50kPHOezd+LinmUH5WqwgNUPc2b/mvhzTDKknE0oxUugQrnoB
mGwnJzDaa9SH4SRmbdw3hnsanCUU8Qlf0wjwgtOG3sBx4orq4k8ws19Yq8jtiDd9
i5sXPiEIEpsLurGDY6YcvcifaSBQCmvbv4EqefkJofhQpv/T2DqfhzeEW/83j1HF
nfNy8XUnQXxSSmDt1fs0jmf69huTDABsXpQSVR1i852U5XW4X08X5f7cukhAr+1U
B8wOd8nR3hZL1KeIWtuRI8MqZJiHQuWKxMK5qVvXG4yZ/Xm/PAb0MbemCeOdkyM9
4pfRuSYDaM2TM1iJ4aOd5QoHnKGfx++UkKEBKCpe5mFFeY4pD327O8Cc0vOM7LOP
ewIq9QBLthSqinm4AlUShhw1Cbj5ytTn4KM0Ouh/KZ8/Uzi6f4zxhPatbCEKzdu1
APAq88oJPVdB1AzRkV7/Mhva/IvK6gcu8WnTbj+nVpAhF2zHW9+UALrdCSoLW+9C
Jh9wprKmjGLo4DYXaBy/5ky5x+pRiopdwzwCKELIWZXCHu0Dmsx9inpJdHqKLW0m
7l9iWT0ZuuuEVowTFxdScRNTejQWlvA303llfZMQ7qJrZ9UAW+JDO95tKgOfiE6O
aS98S579rne+1pLQBrzcbJYRCUz2CCvl8LrzfuNC1gPkapz+1YXdFu6erMArn859
Qh5+TzAW8aNFoz7fbXDpNHjwMIWAi4wb1PvV2Bi8/Q23FrVM2xyZrCAX8V8gAJHE
mhFdGXHGNVCxvcT/PJV4O/BJmmlq5ZX1vQCVB2nuUHpQ3mH8/83gjqfdKINUiZ3B
lI7YaJKjS7T8T9HyJ7386DYwAysa8Joq1mWNFepk3PZa7uRDEdC22A4sLCXu69FV
TbewPjuco3cT7uzWc7cHCbcQLF4sfJk/fOxPR0sPEwCfPHdP23ezH3wjSGYjn2+J
clLgmsWw1lPFNBH56jPWcIkO55nWXN0LlzQKtjP5315NMp7ajE/ukqlGHi0FtxkN
B31IPZ/zjWCQAzCz+vk5ryidLmz1JnVV716tFivp98e66r5s4ynUyJqfo7clLJ6i
oH9L7mFpyhJGe3fwthFqJ1aoJiyUNvwQBcG33UFJFC98aMJ/kr6F5EOyDurXZlQn
o96Muh3H47E+7jg0Lmguh3D2pGs4F3fJjVIDgl50WiCm1LWp1zCs5H5+0hC3GXzl
RIV68N5ZpUNF3hfSfjWyv+tympXPIn89YUEG9qxw5waowuG5DTm1cmrdZm9+ZQgI
jthg4OP9IqLPHi9CP7zDnUsnMLr+6yvcbbtem55OiJ37c/OElK45LYCZb1/e8FiC
aQblaWQDQKVpRPVdbP+qYhA3yq4wpWWDNn18BKyixG30eicrG0ksmEFvuCViFccU
cyQV9WCxvdtVqASkTX7zoMqw18QuCH485oTLAsEx/SokVriPL46F/U+UAHPwta/X
38r23n+j65YYxIycuNHdKFE+C6iwWGDM/KZ5e5t7J4k6J6UTMDYiWXihWWVSkSaa
WAOP4PZ1eaAH+oI8dxDCFQONNrAYPt9yGT9HOtb7LWLKYCVxzXICOtUwkGL7A+DZ
3feR3gNJhe87v1V3XQNxrGofnL0Lin7F82Ee3DS2oPk+WlXNPyHFMW2UyqjiiBHC
wazhDD4aIx0VlFx9gvPdpb5xCYS2ACRDAehWEceyLqcqnF2aXDw6FPSszS+D6S6Z
vEFOCYrvyIhQ1JY7hhKXXTMJFoLDHRwiLlAvnLCgN+6QH+6JV4/wNf/thCAvsPLk
KB6itu9EqPS/RWOmQKwZkBA2jWlVQYcmPUYdWa/AoM1sLz8xhxzijnGzN/Vv2UqJ
ov//JFL0J1HnkMTSjXRx1w+dtxu+NX8THpoRvngOdL7586lTfYNGW5v3oZ7VzgYD
sQwNpdgAetisDwR1WaSeWpYzcwDvuogKTFBCEMBSLD7mg2shf55HMAhzKerlFszM
KkwcREn7POHAr88Hz+r1buzz/8AMsqXE+CQ6NtfqTBGdbQi/TcO84C1T4TexULhf
+JmgMZnJktUmknHDHFOLCcy31rShuqYpKahcGuSdNkCCXO/aEAtXHMWuw6EmZcKC
FLdGXH25KeGCXjNiqicnpeoKsjbDLrTRkoOtRdKce6xqFEkr0jm8hs0fUZrPNyFy
O2BrvN6+rd9bg5U61Sf6tWKmD7qvo9c82B+0MXvji9bQAhqgPddQo4RaIVvyllHu
lVGhlmCgouNvplwHDXBhsKpPPoufEfu1J3BgnJHmifq4gwCzaGMgOESNJt+RfuU+
mF1ToZy+MxaXsXkErg1Dfc3qdxRR/CD/OUJI1cZgr3qUqrNeTj23CzEcfVXNyE/Y
MKMpYONWMgQWOCsqfiKC5CP1v1/yrp5rpOISK1V6vEH/OyH55xJpU9zTuS829Ka2
3Sidrj2rrc9Isu6IYBvbCRpIG1KUlj/xWgHfVrKHjJNLXj9vOkpS4f04jqzohZuh
d7oaDxEoZlo4cArsgjOh0n8zsryPk89vVcqECY1f+5/aZLc5m6gBn4Sog1KXagRA
YPKpwAEWQ2cqIp442U9bjtq84YlOsmfB3WRHTzrkaG4uO4/RYdI39OF1ljMoUi4P
1Tk0jQc0CHTbxfcyEHca28bZ5LDi46pUH01QpAvsySymGeDHGWNo9lcTNJefdvST
32+5t/o8xnvLo3KKsPHc6Dl+R+8KjCEkrHuEYL0ZFQpWhTlnO06XDUX9oonNvW2O
cAn7eItKp+73lo4PloNizZf3NdzriHEORhjHaMqCfF1/epT8aSSHn70BFW4b2NhH
hEbsfobsukdeMEM6p0upGDXq8YcfR92vxy79CVPSfHzFsWmKktpmFldjG/sCpAUQ
Pk+lhGxs6HbSqEsj2HyIRVNA/Dk1TM7ydq0LCdjsgvrtNUktuHT3LoVZb9qDn7Q0
BzpABgjQ2/+pbd/upVMqWAum0+HHSe9hozkPmKI5S6IdwlYhZgZW10cVRvVibdYA
N1Z8ZdVZ1a9l7js7ujvewHPJFdy6C+mdPI/dEihreFM7XwsK2KYTSvRNfL3mfc63
/AuWJgqTCMJ0nyI3eTS1PEesK3upLUTFI/vkrxUGQmw2JjFIrF+ue24roebYw90a
LIhEDCHUI7gHCJaFQ4lBUqA3D295U0OvurvtsywbIR2VIQ4MRwvNuuba67+WfvE2
KF/a3qibvlMQGMyyomaxShOy2UxJrqN/dxhagL8BkyqLev17PQM6fUL4cmBIzEdS
K6pGP1hwLWgJHwDRK+6UzKyNO0RyDlppf4vdqPRWgNXoi0guFlCJ7VuThHSWVBYR
nU2CH6WLX/TTBYpedV7A+3GsR63nDgwYGSyHtyY+scjejJJsd80sj4CJJqdIxVvb
zmGQ8lAVsuF+pblqWhj4jOzL9UR1CTBxx/u2wHBn+bXWv3cLkOOe/umb+/7fNane
ykK94qkQjuU7mdw02lZiebLlOi18GQOqaK+1AloaduEXOMpgz7To+jss2HVOgLQ5
RyTa9XxteYELWQiqhjgXYgWnN3G+l0EKFrIv4v1TmPVWsRCuBZg5v1CcGR7pGiKI
n1yAV23jeY8cPraDWUPO5OjQLjiqBKZQxr3WfR+XFCiXRqlJfxIIKbU0w/ci/cZc
vKvGxPIcXzZx9NTgv+aIIVjC5mBDa35ylR29L0ih3zqvq+1EH80JV714MtM0jD8g
OyEY2FW2gooktopdD1aWNJprQHCPqj83XFWfpQmT9kYVO4Zrgn1IoqOTOuV1tvC0
Fic1GZoh77AR1i7PZ5wV9pG8qsKyfde9YSt/V+WZ4Z6ZO/2Wi7W4kOBEkfT2RVz9
VcAD5katCuKlFsAOyQFEvLsWszFVpsqSw9Zmb0wHpR7DRCzQAlFtAAg3qnVla2ai
AO4dSW2tXkimvHS1fydeKnOH6jUASgC4CqUkY0V+bJ2zder1c3l26Phi1NCkIxYE
xEzwF00cO6kF4sneY2RPA0DSXHYzkMRDomV0fL+YxsekySHFpHUs0IO56zQzjTtZ
BAQxLDUm6PRSCS/PRryf9KEw6/F7l58ooAWjxwQcfL1hgvqI4lMw4HwZEMH68X8a
n+MvX8Gf/nCifpciViC7sYwg0fsv8v2EGm1ghFVo9K4RUe+xgNGiVQy6ojfXBBCS
ytoMeRm/KPK/tz5tMPwIh21ICKa6fjE5E2HNMkyEosOsh1Co8KIfn8tI6kquL6Va
h0WvoxICLPZEzzSgiRcDYS4cQjhS0LxYY0rRI/SFDQPdzTOwcnzdfp6VCAVOGJzA
EOlGtoc62w69jo5GV2Cuhf+hwwFu7vjNst5fLVz7VKIALN3weULD6shYFSnDLKw5
5M0lpdNUhsrluQOMPF1nQ7JDI42RMhdFkCSqbL2pLIPgWgUfmL140cvUgY9OZZnV
tx2VlkENSAc83tAo2sptUSv2weQw7RJR8xYdSZUtjIhtXFyD7OYxh2ApTT+Dgw71
J82uns4gohZCJxP0V90gB4/jdSyNB85o3X4bNNC7PpR/FvNEciZLhsmkc/YnOfnR
zP2cn3ZLlZvBtpFJ8djw1F929cAkuY2PoKoxqoIHQVwjr6zfn+KGLB+q5gNU4L1r
uWH3WnKByxGxS0cj0DP81+Ofg8flGHuMiv2U6HsIysD3WdSq5Nh7fxPFQdB4CJvn
nHL+Ji0ydgT2hvJZBLCI1cvqy/mbzB3ScxysGtLVbWk5tSvaOzPEYJDFIxi3UGTa
dG6tTzdIgdJWQm5BCmw7ELxc3h9TAza4GdCqZmGU+3xQvacayi21UPYazZHtCEkq
5EHHPsrWnFSFGbMngZtdHTQzgXIMgi85GFzVkEjprgX9PkM4kakweU2vRxmz4lhx
NkFTnL6Kv9WgaaC3Vm01gcsklEVuEONi2jIvTGnj2zF3avDfwnvgkKKF5MDnUT3N
ytZARiWlQ42sFxMi2ZKuw7h819NrIfjrUs1BrE4AB2vUc7RY2w7YcCnClxKRjKL+
jT0ICGA93wJfG7/TXr3BVviGSeLxLJo8PZh/nd0ZH4GxyOOV5Qp+5gEsvlOCWAqh
bOIrsHvJBWzghLS+1/F8A1EDufXekDUDx7rQ9GBhE5HFgr9rw8uvo0I3/1RP6TwS
Zv8naW8vZRF7t10IBMGzsLGGZj2Sx+r9fDIosFV5999HOLmwCx68FPEs3mafH0Ks
IMlnRux0fmjrt4sg6s17yqmeLze4vluFkKvUfjDL9kyONWb006VETt9cxcm9x3lp
FaHNKvUfqiE2ZIk99CAc0drKAe6dY8La2Qm2Sub8zw/VLkV/QanVsRceo7V/kxTR
nzVo85RS2iG/IRcePBvYE7SdvrXkfrllxXA34JjCpLo+EFburn29i23Aspjar4MW
0sUbEOVRM9UB3CQRiN4gtJ2sBRHX0EePI4efEBRfgsOhcQiIp+RcyxC3duEpEQf9
fK/aEs6GfxUus6QHHiTlzCWIFK6sxa+DnFPB+GUaeq9+VUnYgY1KxGXcwalXy6kE
F6y7blVkT+zEuhR55g6nGlKs9yrX+TRIyN3uhzx0Q/xdHNoGHh/DbRdvetDM6cvz
UF7SJTkJNwLmjskgVmR/nI9uE7jaGW5hxpE0hKXBU+QeNKNfl4IGc0zHXikgvotk
ANVeoxiIHt0wnzSTa5EM30HZawtrVNFjVdzMdKknpCTBkhdF5Rex8qRfWloAZfkW
6H/1ON40ty7AvBEiBxkhxipp35Fr4RJFrgzHZVa8nHqB5/UH20aMG9CpodvdSf84
XIh713fxv/zU4j6c4TOrkmysHhYjDHPAx52gw9G30DE775mlDkRL5VWAUERQQngK
d/WYRTaVEbsHChuEuiJZNviKX/N825dDCMZ/kYjE7fl5H7eZNQ6jj5vbyswteU61
Xm2St5r30iPMBiMXXovECYy0pslBUu01niAwp/EM/bkiluItuCFA3vymIWBBqmU8
hokMGotFXcMPnWayZMiOWZ3AFCiwrngeqe7LM4qj23J3+Cl/VACPeIVVpay52ux7
5aUxtIRaE3rGiy9uwPL9JP3kG84N7K1sD4VGj9uHzUh2zq6E9oTkvnwB2d2fsThJ
P7X/VZIL34eyQyA2h93r9Ry6Je28eZjscQsxhyCDadl2o3Uuxd08lFQKgbWoaw8F
gdACzaq4oUfVzvLG+pap0F6rHpi/3kZBHp8eP55EAD/Lm8xWjR2jpQ0A8oXQ/z8H
1GQCTPsL0o6UOnoZ5is1VpThuOil6J9WgwVxizctnATK9o+lmNViJS2LoRiZ4bYB
7ZMn43G/Zv3hIlODFv88ZJ2xo1GVXdHuBLKBeaqWIRPLNZf82wiQgrTHkNucI1HP
YYFY3T9We4hO1/XfudjByz/J4GxARHbOl5gz4dTLM/1gkOkEHfGogXZc0TGLETQv
Wja9MTib98OAuzniHkPMfGFA9mfH+l2yVgdCijSnMbkOwxx1SKqIcpKC+QcgAMiU
zL4R7WhUyBK9sVD35Cuous8VunQKpC33txZu1lffstejkcRtvQAVLhsA2ZIO7GL9
Ciowp+MZ6ZoUqHgimMOxuBx62+fIVAkWB3Xe32FpfSB+AVHSRswF3OroBYodah62
SNpXpjZ3v6I3hPaPYO905iOKHQ8gLDqiX6kyh9n8OHouAzzqpejdk2d3cSOf3ju4
KmkjL0Z6kwPs7D3h0PK9Dq1rdN7oT5Cuh4jOWfiidaFBhsZvFT45EnSRzOiP29ms
XiW5+xsV0r2gxfDIMzL3Zl69DIhIKnMsRP0/moAp+94Bm2Xb0gBx8pURf2ev9l1D
XfPiZchOtDmOwjaYqCYgEYBrBysJ8wXBtoXEitRXOWCIXlVoUB35jVifnBGBAn0V
Y9wETrokZprkyyb0/Zyc3C1NzkLl5tFO3P0EFnlUWv0Pasqgts7w+Gl04h7+tPWU
/9updS7xbYMD1Q6chtw/OetW36j1aUvbpM947hXlKaqkff2GMRXLtAqpS3xYjt6i
oCAmmejmd+bVCoHoHOpv6pOeSEJXsImXSFio7NPZ7oa9NdzxMSdVH9qFjQO94FWk
1b3TL+80McGPaqFnridQtovUSkyQdk8xTp2DvfR3eoYaKVnBgck/WIl/4ZJ9xgiA
k9LqVv5gByQ2rBN5VwsLdUA4CS5sZmBt5UN96Woqjz+26LCnQhtlWBaiPp4XpP5U
8gLP2fnjj294dSJaHeIktn2nmAYOzOonmj/+ezQkakLBzmQyFO5PxcBBFZ0+iDNt
KLlQ9sIwG77ECOvUF8RgyaY/WFmrSJQfnGbGH/FIr3SJnr8CSTyn9zi2N8/OD/xk
KUdV2y8ichWEqZ9AYeLTK6ulARLdqlQ+R9lwuZHNXL8UXMEmM1gWjIndbepHFF5i
Tf+3HaZog12x4SJvNgo1ssdWfYC+Cdhgs8m1d2cjfc8lCJ+8FfTRXYNGg0zVVxay
T+dl9gvmdej+AhijZ2v1zyBAw4Qc6ta5abq+4KGIImDW5ysTw8TJWdITv8hh31Lm
Gz3S0PbPmQLEvgRN1XNzW0u2ifiCrsdD0bL17hyGMJsRsstyp/Rl5WnsnktnwUki
qy4uDFVORVszsT2o9PegtFb3G+2BgiCO3B6hmESSQ+u1GjNw0jxkaHnddFY1S5Jk
PToRxheLUHY65b4mNqaJL4zblojstqcgcEttqPUw98eDp4bzTIqBj1wiGKmV9HLo
POshSBiZexBMnsCINX4FZvLRuRrKJyoW3gLw1D0SqD4hN7moVQU+/pzt/6XE8o8t
A0Y1wtBfgrkbi4MgnTVJxiVjkqIhOR3NVCFmYfZoijOGTpEi7OVBxPl0lOfnBDjA
DCwmBivckFh7nxRSCFcBuTs0J8NxU1Y0/xmvXgn4B/eFAcdNXN+UGEerTmD9V4Gu
NERGrWKqsXAaGNZDhq0hIwjhuy61oziNfC2K6QknCIjUomQz6MYt/goWGukCg2O0
y59c4Q5t5mi/vV8Zpb27tN43CHWOlmtLMRNDe3AP8CUtfcsD041vJY0AiFyvDW1G
+qJlfoGzIy7EKb6KT7hgCNrn4C4eu4AR+VlVrSKH7M9rEn7PUqMjrwt7RYhPyI1O
5+8sumKEBhAqjLTwVocGKMc/rVSjusYU7dlFvGDvKU7ZN/+6XqYbXtxDr8aUmlee
dDCxKW7pRuMUYzpeZ7KjN0SfUHqd+Izmw9F/+NakuPv/6cRpewB43YLpml6HwZIX
ROkOZfBHbyD2ZvRkqxIM/8pugoL5K9cbBiQN9O/5MEQ/x3irRnRDFCbQR3OCZnC8
u4pM25PsryrMXVbwevec61vyol+SJ3PvAuElTXkVOBJp32JuGLlqBxKFBe9oKzEa
d0SVAKwfTczKVdgpagxiS+PPrzSSQipZMbYHltxn2H+WZsoQsvjOL/gIifh0vgyI
7l6TK8LAQ10CuUJ9A7UGhamJwofyXyaDMnNMK6OrfmOJq4pKf+Ouop13hh25wgE8
15XepN1GqOPP/O0lgjBjrUHxyXeUlhi/zDUySjcIhiOoshgspVFhiEUERFpfUkT5
yI6/2trMSJ31g/LFhEIUgX0flUJhekGpXEMJ5aL8yYGllArXgkwipBq6O5npXW1Z
G8pqI6LF75TTwcWUHN6E1JCHiyM7k+YgBNfcVNa/J5PqL1CsmFlmsoCopJszC8qd
sTjH+QEMDmPOqDJdGKuUviElxuH+/zYDeVBy1BMjl+g5g9YrJgcO+nq84qfSsSK3
ftweQjyAlvENpcZ5LfexMqL1WjBaWLEW4k+ORpJFQQ9QIQ1rFNo6ODhvEXS2En5v
8tBEDo2xJTRvvOnG4llv2/Ocx7gc+pHJlW0+DIFnJAlD54lMddLUAjN0TIPYcuYY
ouNjFl5jdLqhvFKno5+FbHFJt4Acu3Okp+RE+XREkmKVhMozVSVEGW5NKw2G0Zsl
EOhu4LS4SnOI8kQMz7vPbh9g2NDS/h5RTCxQ2WHwuQrbICG7/CxPTig8SHR7O2i2
8nKDQ8yMWDNSrzRF8vLVkZu7cGs2l854BVz8ErA/mSY/hThLzuHEyoEQtLowuA0R
m8qkmpD9m3Sqtm+C+/Yh3Umt0MXrLPguSaRueCjStwNZXvWxcYzdjlDkx5Hv4mFR
ZX9CYNp/sADD8JkRfjRlvgaEynejSPWQWSAKst0qZcYmbfUlTOWRKkEuEVMSQsJL
d7p61PKlXh+lPTuBF/ClDuQ/JgVLpieFiDi69LZ9xy3a++16Ms60pVXcrsLmOmhi
uKPFo0+Y6RkKfIqAXMZygBy9glyBTeo6PPxOpTmu8YqftPIIE10GjDnkeDmVVEkF
ln7dYxHxQcKG5YPyQ7GjBAP/C+lfRxpUPwAFAbefaAj3yDWUKNA+HACd+6MZLfCL
YI036nvex6QXga/cvprzvodGJ0/iCDzHldkeZMCazJSFrH9AF5ML52f0Uabu7Y5U
bVbWYEQmAA27+ul+Sli3I88FjFlvgSh7YLqae9skGUWnjTxqvpOPH7f2oPUtw9fn
Fgm/xc69PmMC6sSWY+TuZwcSeOBu/83SKmozM5MpiNmuKE6aU3APl90XXOSqC6mf
94iqLEDP3Z4P4j6ueu5rZy5JrawappQQxgXCD1lkXZibv7BJ3aOzjsdEMqObVvHe
7ab1tYoEWTYEnisqyhGLd3TwXhrotlGhjkfwwEhAHu6nkZjsrsDifDXOeOdJfAZz
1VOidMPYye/s1iWHYwizySXNRjP/oNYaiYvD6AwDR4Bnaa4lr7LfpxT6td2HWssI
jJrv7GwBDVotc4qu6D8+GXQmYPkPpoUTUvzxtdreAJdZwX4ATS88Ic2uqM+pfVlJ
OhUJYBJMstNDtiXBVqqbFOaBRuDgsgyOfnzd2xFH5EYoIHTbwxDo9QMeJXm8lyB7
u4CZEB1wNUOfloE/d96wZmmxXwizo6tm7xXpZ3k3LbICkefyjI4BZSLPKvfxOtdv
2JZWr+MakQjIOpL+2sZqUg71uMi3EeZd14yCmcNalYRSjD/uvcgDY+Otr6AQffms
0GOVcYakJ7YmgWneH3Ed2vRyui1IDSSIslbjlHof5hJr1y22d4rlg6czuMqOX81t
yFEQQSEAkiPgnuC9ro0DUQCSBBGzsbp8HxK9riw20cfSYqUYjRF+H7mwOrNB0DkP
E1M0jDExxEbS6SKtZj36JOvLxh0B3yG6hyeDp8CsZxY9TFvqKK5/Pq+C3MhNfLnH
xrjMTnRLOUjbt9sFHksI2xIuooCR3v9hMllBEB2ZoGsM+/qD4tDs4SMXMCke/eX7
NopeFWzGqEz9f2PB0Qq4m22n86aKAeL998V2qRR50KmmaiCtqZqfHGXL6tHkTqjO
ozLYJ/d7sWB2Vij9l8BMm23U3tGwpIlZTscZbemFQ8pVQi35tAMBLRHCfgR8RtQ0
fCPi9h0vGDK5U3j1Nhk8nMb1eF/4zpr7aybyc/+xYkZqqkM327jjKKCHQ1QEofDP
5V2LF4TvZXOb6MImcnVfleHOGfOTkxxlIci0ZkPM6hJc1YOU3W3TJzL2FXk3mExZ
aBR7W7AhY7tWtYVqZwUrOBVt8NQ+QyJFI82BKrr7G3Yhbae/zR0CYAiPVKEkmC+l
CF38DpJWcsHghsDzUwqXckx0QCQ2TJxlNHr5wjolvzKMQv6q1y6xVtPqmV2Dis5V
WmirZizkL45vemdE5wOmEghT3CJjHAsoqb3GxJ1cAS0xOTmPVpjGk5mnkXMKbFb5
8Ox9LQctXaG0jMOmiuZGHAYvV06hmejpn0D9FbfNK6fnvKm/YmGdusmRi7FjghUr
Y48WpUL7J3LfrmW+qi+ejMr0OaDwiOZkGbvsNMjBhWBwm4mSQli2lFFKVy4ATIFP
cLDr6MTlKnH3CScIk3hagdPl7nnSEgUTcVu2YMXf7jeAw2+JDzhQVcA6dgg97KTO
pkda+UcWY0oe3wvXT7OASJoRXsEKSj5ZbI6eD/CAsz03ou4JaChrWfH0ns6iWRad
CuM6EZAl2Hmj6GmcCCKKG4dlqyqsKKIO7CmiY8ugVpLOAB8hLsZaPI8TauvxG9a8
pbd1HiBnf1XUv5q1Yq4BE/FShB2Vuy0Xf+2/nnmWcd0UWqMMsd/BOmY7bz6R2+RP
Ws+dVyM/FDiuA5jKJfnZ/agi6y5g3rca3/wScJF4gsAjav5rZS+2UNmtGRUZ+LWG
5VOtdWwAQYlxGLJa5zpVTY7TYPdJ6yQMVFTmeHXANQHiePPErqs4naXqUempCZ9r
YahMxlznwDMa/U1e8oEtRN1Aj4WAGyfl6BFXGzf4aahcFIEuWrQAkyOcWhPW73i9
FZmupUGXYxFGNgHrstV7tdu97NTE4KRPZU2D61lgExM3Hb6aAxFI3pWc5119Zh6R
G4++gYM0PwwONDSDlKNSjW6yXHRZGD/SBXyqhasIPCXnjIX09vWTilFp8KP0OWYr
nJfx9fal7ozI6wnwiQP8XpfpWfR0wl6EgUGi/tWzkU1zdf078hGs64VD3vmD8/Pn
vaKi7y021JXFdhoFsvCSwb78PC3r2pjYp2riAXgUxSVR69RrckoW2akf0F3fCimn
OVVzKHv9vfiHMGe/asr9FIUEUOSG5hYZdbKEIZdwhn1r0TeBu0dTXzDtC3VoM8bz
v9yiq/9+khleA3s6RZoCAyV2hMINvnbXLwtDK2HVT95oSeVCv/s/wE1YGEQzGisg
FczxW3E+VA+Z7l9sbpsqETiogYWXJ6i8UewR0KSRQZwEtHtshXAuAY1Zju2qdNsR
vIA+85NEIyBwEX4Z7Lp7qHvBHc9aaWn9r840RrdHDe+wBdOJZyl2/K9+TkLHPJPQ
fAcCuexWNhwNMOhTbCNYfSoIyXm7l3DIEaDtymYRX3qfk2ItWQrmkTrwIrQI5Xmz
XqwTrBQ3NE+Z1jjdpyfQyR01SQ6JWhzmmYxwweXum/Av5jLnN44u8C1ecFjWNO2+
987ogD56hU2LN3jOeGWWwispg7ngcDnfSWvtQOUmlXsjsrViuy41rRT4oIy5UX+T
UietTkrbsViaiDEO5lWTnwMZOY93bsW1+yc1sfkr4ULzWHHzU3UAgl4EsS/976vy
wB8uQzFx8PhSiB+d1Oq5ilAYOOvvGRTkyQCTMChL2a7v3/RGfMOqjjqllw2iLOJG
UzYQVZlwLrZTUTipc2kB0h3i2+s5zyyoK1aBK1q6K6GALWeuN73FNSRksHyj/PGR
zy3v/Pmx/eFGQSLRhFMBKxGpsOxbvztN+GWQg2TjmibqZDcVvdtJqZ+cHjG4c3ZW
6bJK5LcEBTFqJYOZhwLzfZZHWuYoqtN1Sn8etFDhdW25I+QY8HcXSjszS0gutzei
ZRYDqm6YvH01U6/kk8jBvWxwt/zhyLillHwcOK2Ul9sUkLEtHKKGDAekGQfhbEZJ
etBInqjTE9SKBn4NzP0kRxHsivHHY2hW3INYME9DiDqPEXiogZIMDcU4l/4791Qy
jUuIMfK9Pr5gMmE8Z8kpD0XkriLab6WbBIex8mxLLRqfYwcESnKFg4GR+ZyMnuax
LjFa9Wi+2MTf6bcCQvpvxtiT0H555HQ1CWkyiuqoMEzGmNqSrdRN8vpCKSv5Q5bB
r5a5F7qGHDg+0pvzX8imMrs5A5sClUUqAsyM8qrwSBnru01Qslk9qGV+qzQjFnz9
NBCT553c2enEeuotGS4Bfl0BB8CLh7LzSS1B4WIMgXHITlEoAcpd2vfxIUHAh38A
asoWT8STUeNh+OoWIGQcUGMyUS+NxINhHCV/Xw3vZ5cLD4Aus3Cxj9tiCBSZ89UY
nhPAaGjMial3n4kgaIz/z2C0Q+Z94HKy3sBQ/bE5prOtdwbiEjFsbXzT1bOCGL9+
VA0upQ0e/aqe1BSWAijvLY1bE3UZXqhEv4s+NOrWR1G92Tqzn7fhJhDHbG3+0gFI
57GiKc/wLzn3/D98qllPlomEQQE6wRXVT1jPzfR7RTURuEhikKOwgFNSg+JR4w0e
/eG60JlJTse6S6uWZSrfAcPibp0rLuMK+lgc/fgcdKz/NpQmpPYkkKZWi9dFoTxd
LuAp4MiqK/SazpgsKNfFWXpWAJ03j/MQ6u+nYsg8nZPc3nB2kXPWme0mC86xSx9y
1PiXMB9GXl2qAzmTtL/tOwhLPkf6CxoDZXaPozYwMbGkTb84qiyLsifDAfNDmV1k
dRgaXlbfhOJjIcciyYu/wYmuXvE8UOrlGHdeP0BAG2Jsfx4XghDXeTg9brj1hK42
rWTJBTQERxBo8bXtm/bCMXWytUZs8Y9trWtNofsKp4nuFMo6C3ECrs3anNjnqLei
00URKgyBUaSMQhRVzU19xwLevC2fljjnd5IV+DtkO7B15RSt3ZY/n6sa3fg/ULeJ
eH4DIoAgylDSG2mQS7KmH0mn12TIJieSJw+FItkpRy/befCsXff7RWUI/TJpu9yG
3aD076jV2LCvyeku1zWWRoAnXLbI3PhIpVc092RXJOf9RGdSvUOgMP9V5rjyV56F
8ObEyr6dhEHesihMjS6ngwdoJ/0gNddEiK9qTpGogI3VCkuQ3YSwZt+uZIsbwwEr
6Pz++dKjdjrkI5tlvbHqT4T2tmuXnDWT2KbWw2EIjudbMVGbK0j/qQUk3Kqcp7pg
slIQBK75FoMNC9vIaYQ2yY1hJpUlqj0PLRVw7zFtypepYW2I6O+SuMk+97FQzUAK
2QoEs9Z9P6QYso3NNUCLXQwuIodmmD5dUyTql6/5x3KKQsIf94UsS6AfkrCNHBTT
x2F77agANVcjY9ChHTCgruOcZgrMfu7CsRtd/VOMzfZMSBlYnQGjTqFTItMQB6tQ
qm1ugW6sfXQsWGqM200cZw1ZglpTp0lCjNVL73myDj1Aw0tNgNjF/FCr71ELtg9j
U5kcHTBbFmrylrD8TX3B27G81iB6Za7C37TBZnUWuX3eFeLYKH+ZztTI6iqEppEm
RWlmVBAjmuVgFXncSy3cl+df18jYNDPMZKV20IFJYk8K8OMyx/zdNdfzpWLACve9
1JcwvTQn6X3oabZDDoA93ZlDOHCZYDxgggF7OBEEQmsvRPtA1LYUWlxNolb4pWrD
qVE5Qt1y2eaUKIw4mxAGFsn+LOZ+DLRfCO9feiuRC3UpuhWtfSQrZJ8dTi+63ihc
JrbcyuyWd0ysUXvQeUh0Ovm/VRs0CqaoRoF4SXF8HwtRTJHU8FJeJWLbJMpcpUTV
QMOXabSMKgzYAQRDiht48/rLse5/mDcQ5RhMKHyXetWdnyKqy0T5hmaq4RjVkGE7
a9mTrdMoEm9pORy9X7VaFS/RBdhm1+0ihie4H6O64tJfEO+p8OKhabdlkrf0Nvva
l8NosCUBzEIV8a10ctqbJP8snicxvb7O/mdOp9JG+wSN/DM7u7I2y/sB/3K5dpQn
mE1kHRRNQqF25RhbZ3A0hgOe6bhc9eKVRT+I74/ZdQ2Zr56MCro0qppxy9BA1N3j
a/vWQXeZ0w2gP5X0mWc019XvIztpgMOT1JkUwaBpOWeQPnLH6MrKyx3b9CALCkNt
Q5tswFtd5TelyWjk8B/8s49F9i/V+3OYHuIEGgPPkinkKpzE2eSWhVfMIYYWr/3p
JOzxcanldlYcErASFfcKi5rlG2ZPxzDhW2nrdYB8z/ZSFIOLCaeiTvWUsLHxWk5D
UOJq5jqcUP6O4xApGv15UwUGQmhza9leCpg0uhOq7+vZS0W0bMMzBUIu2dK+37vg
575spcATWJTX27cx5HMZNLaqjj5uo+EZKGQMP8E1h4e0ZAclJsNs2DFWJ1pLscf0
KjgEnob0mbkQ3Q+5fbxQd6h3tjPi8/Hlvjfkq2qxX3yOToCw7GXjvrkAHfHpeyr2
wkHKcshMygpngdNWFKssGpbdDj44phyNrrpmTP78z5FcBetBQ5LbrBEYzfW/geOE
tCoQ+LLHHBxlsyMdeLVzFQKfrldsWt2jZ0r037gCtup4lxLVLhmMe2dAXQAKm3u4
y3UnfVSHkGB8myAPdCwu/tutF1a+QAhPmirqS/+ligeFPdFjaZ13kCjBrvP8WtVb
PIBCv18jqpc6hABijZLegFvNUxgN/UPec+uwwogxkFLpV0emjprAkml4TDbcMuHG
SPrT14tQ/u12TGBSbD2OdgIVnPay6kpi1tl1W9MscZhGJcodWVArq5j08UgbkrOz
e/E/yrIailE6Fzc6bl3q2niEZOCt1Ls3p4f8i4xD9E0XOm5jaiuqIbOZub/05Ycv
0L/YSIR4Y+BCxi0pu8ijoceonBTj6CcbkBZP5LVyLxa/2SUMZLHgnAuJZDjeZxCm
R3s3sS2acJj+NnGBgPf9iwAH9SrwIFDNFRfD+YErV2V+1SPrLrXWtN2FD4GW0ef8
OjUAi0JVyPDH0VLjk7dU9Ju5dQajYeq8K3MxdonU1kIHXaxgCny2XTZMUkEt6NeG
Na09b/b5tuGibbenIDg77m+cTd5tpvwak7VIkJUdCt5Z9fyPzEvH5TEDsaf3yHOY
y9ytUFXdTW6iyR8zQlAicGkFC9Hj/lZajtxWz0CjAl9zpG9qNMOelFx+AYyPFq4D
bXq8JruuDMFpCFjmU9Q4lg9ob7w5t1blQPaPMx7TORuEO8kEywVdg0kAUd3l0Iva
OEsZhjiJswWTrg5rwoBixAxYbgvyiKKF+FEcA+gogWO4zBiLJVBF1XVQAsn0vBxT
6PEJJEJvHOZb3XZsABvqBq5NePOVXo8dh/Q716ts/quUUs3cyQjgzTzst62vmD28
wjk3LHXZDJg5kC3dGnS7BsnU3M4Uw/dKxopWDw4FmopiYywfvGLzn5/uiZQxG0G3
u92ODikZRr2LHlvzR1sfFmR4dXdjfuOlP2ZZikATZ0ZT2FjZeNj639IaayvRnrkq
vVoIP8DCkIxn3rwyxXqW82FAgNLbw57T9OrhCoXhOR56Z435r8PotXzwnzN9xFhX
f8aD2l8Fs9YJbeY7b34vNi34f1I4RcvnVEKNX3MG2NaDxATgUs+XQpgn4utrhUde
5R8OJ9c0GOzZA/Ol//plTQ98Y+N7++8fUWPdn7uHWo0ndiv7J6w2bMbHGQUfhEhL
t5swYAx6G/ISGSB4A8KF2vQtT3/iHbYTw1oJgNsBdvtA2EoaDMsikclUPXzxPcq7
PZ6a/0n/d1Oqm2xnP2ZZa/m8FHldnDkXnhjZ5iymEBKU7rE2GVP+AUP06oj28bDP
wGDTEBTeoz8fQ6u4ifO8xGJh4yXo6cD50UZ2E5cGRufr651Vfr5H47r5euKF7k1n
oQDmZA6JV3IvgUrUevy/2G24pL0DX6gAxjTgT6vN8sfS4TE7ueYPc22RXXPftyyt
iqlz8fQJp34fIJL8pjFz8fVKQcSvb5W7ghzo0OYUSUH6izOP9bk+UkKQrHiz8NjR
ked4Y6vZoT0AtKLBkE/pfH8wmpt8BgIO7uLyx6H4o5lbrC8nqdxq/vhf2xeyd764
aATncetv03VQ6TQZt74klON5O9gbgK+31jkpAoINnP6nLrjU0SanJ8dw2DBdy8aN
ymGEPQtDxjR6rVaKe6tV4nJa8GwPhDaJFomqDKWoaJa0+nweffwgCKtQ9t9lgaJI
VxF564JK17cdRSCPbfjC3qsH8Gts+vRJsIxogKy5Di6+LQ5+ja98drpHdtTLflm8
8beKqSZlfgr/m4tFf+nvqEFnKFVbiZ5foLncFGLOHaGSqbMy1l7dKE8nbKlt8hgC
eww0ebGqBLCi0Qr18tyeHSltHCjdq2hh7AAwv09NvOOC0Te2TXb8R5TQP1gtkizL
SjTKO/Q5yzRr/chwdOIvgaXDbNjylzDC+p7YFTgClHXq4ftAxV0x3CLitD70sx7b
ItvYUFIuTtotDklizZF1kw6ZcPOIP68OS1tJALefvqogZI+lsLf/Ixxg+DV6DHc1
04rsNLsI6VwfIic048aDltCotthlCet6Fg4NsN8v0ocRJp0GfcYabBtHlJflyNrf
DQ3lfLf8G7t1k8BuY+okgORCaFW/maVyXXFB+LbgttYwDgDxj9duNWk7Xp09R/wy
3iEuW/0kJu9bxD6/wTm6H9dM6AEZD0iWplu4vzc7pYN2DgHbcjQ8085VbBUfpvIC
pPZkgfJsKwFEfqlby+ySHVUGP2wD8OUHg1VwINbd5HFa+pgXjUXsK/uVHQMpjKXG
wQxI93U/tcY+AS23RqJGjdvKOxw/ay98EcjM/r2GTFJYx24QJj0isYIqZU3XclVU
e5/xPTF/mIpAy7nhzzPL+6/BKEeua1yGJ6XEPCImFsspmQ4ycx5sUzc9OvuqPhUh
qvIu2IaXW40x9OKrOUMPKpcRT1xG6V5jlzUJ8W5idcpib5JZNlwOigOgx2pvC+45
8wAnmcNLa3Kc3C783VytyLZemKNL2SpPjHvuU3nbiAs+W11V30Fu+qLPP9CXMyc6
P9aj/HVdQzm5ACoTZCiGMVBkUKszMth3I/EuZXCaYNVT0BuhE3yo2+EpS7/WAmIf
1BHV+3Xyt0nMWbsO1JY5obX24xcKhskWMLUAwVAWj8WU46jeQxpSlcVlMzeIBdKH
QrnJWo+NIvrhXLqGuszdv626WdlJde5Ya8eOnn/Om++vY+zmad0aAZegr2wLd0oP
0ocZCMkXIrkOiJtxYGrB00C1cZo/VS9U0Fa6i8sky8s9sNYoT5f8AgEdA4EWWCku
03xL9hIC1wrUreZlpGSZXbSXwfTvGpV1OIAhHXWl702DnVti4td6PBhB/4kwLwFC
XwVe1kDd5jD7iAc+qlVZ2mjRsrg4nf7vioaBEqvwoGAqx9q0IJQve4XqZZf9GE40
u1qXxQCNmfXC53EprPTqvuIZy2HE1eq1UhlZk4PFtMCpiOrVaVCVaCUPppTzySo5
4+azhDTsVvGA/wMImXi/68jCscLpIVLwpJUWFE+lOTczh5wT2tdrfveWkrMrLb/N
FwgBanejVf1PMO0fMzeR5h5uRs9psmW8rpi0W3iwpXFvzRL/zPrSyVp43ZxLIy2f
gndfyXd4nPAWzEJQObcYsUqfGNwBOCkOmhvhKABjrRuiSUqJ9huqej17jPhlL/PR
TfT288HgPQg8X3unA/wPzt9oBO1cGmT+X7qyeCqFvQdszTT7rd7+OfoEY+FF6qXl
2K8izmNjR1YE+vt24do+wvFAp4VAsxk2ncRzvQWjFM7wha2oyx7V4y9HDkIwtHQ3
+1YfZbRgEGYhhkN+bCp+Gqetv/+ZacuD+lyzLunadR033X6KuyEiB7Vgpt2AzCSJ
EWKdcL3aNUBbPz3zp2GT+aAgL7RlUFpDEb374Sal8SDshlrEoStFELaA6hlUgiMK
8838F4CD/y8Etqcpc3RuTC1PZQxx3azsOIubwhCu+4K5NIc18uMkMpHvcXDZjQih
clcfd5PNtFwBehL7ccgvetjWzySa5nve10r6kC7qdU5gUwQysnY84LM52cuylSKx
rajsFeQc+oIjFYqScHoMyA9lJUh/YgXiphAIjW95OTtTGMCgO4ORH5okzjuutOZv
OL5Uhk+AVhkmPD58cvRAN2RDiqBEpYtC+JMuohlf8VO0EsPALZN5wuuQHewxddhf
1mPo73L0dSv+67zYWv26+K714/DpHifyk6QaoifksOWRqd1Pj7hUITv0DQfkCWh4
2CME2P8Qml349q01HnjVS25uh3ncVBlsfZBHJgw3i/Uzh4fmAMzHBeOvOKvvv7+h
2Yn1dXUCKRaZyVvHPHmz9wseCEPW3nX4/pyrfabFgE5nr2DYDkIL42DqJ/l5CJD7
ehyynj1lIrs5YOcK8FCuIZMNeWjfrTlyhxixrgiKAjrwbwmhQU+W8xA6ZcYMZbhl
LyQY/aumB21WWFfVmBD7bikXN/VmhfLBdYKyuq3Rsl6AHURxq+/IBrkhF4cdQENd
iYm9V94isL7Zpu6moNjvW4OoWQ0MPFwEUiteRZQeiX+oJ/U2PrWtpCr8ToAx4odA
E3MS1ifOyeoSuctzJusEnxw3JlEuBFK84fPI9TzjU2f2rGnA6Mk1ACo825fVQzgc
IIlB900IQrHvrGh+Krxu48EPYdDhnmZajDtpJmPQK0glBzx8/DqDsnu27tqYlW5S
S36VLfzCHeyn3eoY2rWedGTJMsN0fBM30oy1Q/J4ezHweG6CdLXMx1/7SCbWmlhr
9CMm4Giy1FJ9KRdCBqljS3eOa4hfCo2Zjl/AgeGD/YQYE+HcdfZpHCw76qTBiIz+
9IGm7Ao2ZtYqqWl8VAvk2F9I8xbUDmfTBoTsrPvXSSznm6c1CtohC/btvcrxrD1A
QCWiWQaHGXR9T3cNnuCFqOu13tQttltuBUH3cPntzVUMZF0gAIlahjhKv1jjDsyh
Xk0Tfn0Y3zPU69Kgk/pVrqyOVAjADl5nvTHksplBruzUS1YaEVpnOB+j5/riXt8O
Dcah3ZC3UhcubD+nkeRBY9TEE6pCuRUT44yM/btQOkM9S6kSUqfTlKImdzXmuwWx
LeF2wA6aJ5JdQHcK8POjq8C4EzY6NQTyW2OEyqbrxRyxRzxsVGQYQBR6MVSqgjeH
foZvTdaIcML/RcnYxXWjiKaLOszr4HzTblKXJOLavSzz1U2VGxWGkrlIGbe3FUMI
ltnE4pEIzaG2fCmiGqffux6uEGjD4T1zpjC9Cf1AYP3N6QwEjyM5Ju//VPgeJU3S
Hk7GTZGsfn0wT0uq6zB4lyXi6Nrlw3wDPDhANICcELtE0wpkD2wBTYVTmD9HWBWY
lH9NgDL+tUxc8W/bm2YA0JaKvpbYXg8fIYGLSVq0Z++EKblaaR/KfG65IsGahA5C
XVHxf2f5MrRC0Nz6kHyRDBx4vV1AehXlmpCvoMyD3vPCjW2l0sW1G/L4gAmjSlnO
DjU6gfKFo3qCVUpvH/nEwA16cewyDmbV0trr/+fTFpEfOfji99T9KspIcLltP+c7
UbDt4ieSSW6JpZnmR1gLsHxXSyVqHdPnR92aiv/L3gjQ8uXjPSjC2jV2WktogGVN
PQSqFxAqEKmMSfmEgPP7PTHkNDauMd61v/rgQoh37w3BjHEA/MAiWq3JmKLKcURH
C5V/6+z9W8fne3hJIKPT87kkeTlnBaTitF0PlmRAjqqZDRilspLNgnU06yrDdbWG
1P9kLiQxg+ZyLvB9+ZPlVHHphT+tYeDXBJxz5jJrTtMRWUL55q25TGGz1KT9tSt7
WmCoZZZX/Ka2UESH4JODipAiH6GXTpRACEDPtgw1JWj4RQUYKk3txoFUDOhuxA7C
XS8dBwxacct2mHgzj73r/UnjEoTqw38ip/j81TGv1eRqNhAk3hwbMnrV8Nj1kg0F
afs1yGQHe4Mlfvat2+TDHE78bX5ZOINolbHsyKOmGHGqtHhJsDPZnuWqK3hKslgZ
3kGpxkwk9nfoCH8U7PCZdmbuQambLQkc9uBA29kSFnZro/4hODHzuZ4frmNSIjWp
4cpV77SQFdAe8fzssWXZI6PJDJRdF/bp51dmwgN41U6br/XBspWSmIg30VdDBp4u
JyoQeH5jJCO1BLbXR8tr69e0jiV0BzGFso2Sr/EbripT6r6ALsW8ECtLyxRYpjzh
XIIhAhuKh+Ba4jaeDlKPhMOG1FMLkgZKcx7y7QIMUA0q2AVlRK1hdKNU8jEtI4yt
9Aa0/rM9BpdtdmfM44LRch+nIeT6gX7IYGqKVUOLzacYHzqe59H/1rn+azGkF5JK
e0a2m6FRH3hGs4XQ38Qvjonk3HDDsglHxAQH0dybo/4tozEsvEoAYHR8Natqfx7i
+xMmtiPi1xI39qZ23I4c/itXrJI8ZtktVnQEHWdj3XlqQ57NQASs3N8SeBjRw1FT
8o2HVXM4ckCqnh0zr99syUaDzTz9z+pyW2YkzFOrxPVKzz/zSXbswZ04IWGnWrjX
M6gdRfkqgUjJkATDWpCf07ctImMHS+Jy3+RkQS3l6inXm+rDzt8XuT20anRaYT5i
XD9co4GOtlcTLsoObkIhwD/xvUkPBi2jEErSyT3+Gk3ajJ1qMTKdjpYhNK6nPWb2
eIOoCkM0EVxpLL7Wpu18o4FIWNDGzhcIIVjtaz5BIAyl6rs4n9f7L20nph3ds4hT
IRd1AshhQ8AAkjoVQH4Do2852WVIQ3Pw7zr/uXuy3+HTivCZQn8t+KLlftKvH0k5
u2qFq+6P+jhCgP69OGwBj+9SwyyG1qCZ1JTqDyMAuJUntm+mq7aGp1i37QbTMBnn
d4cevJmLbcWUEssFZCUL0FzAUIGR0gjDpoeHxSsdJm9rWC59BYfWveT306izC7OW
M2bVlTGzY+FMRuoI5R5F9SJ2e9hWu/gPoIiwNHYjcP/LFWBJAgr/Ysjk+YtGBxwm
mpTCLrTrApSaSGCnWsjkqFv7eu5miyorBSn+LSBrzHfRL6TlpC7N73aBLLYkcNCn
rpq/8RbSaVTGEQLAfcocwNUt5xtX1fTYOUre6gGcRg78wDQEikJDh2SmicOqkU9j
7VrUU9PtoBiTItg8ClF6Zsjkk6qHjydrhK01pzNPUxh15IxI5C8YWRdS+SQR+cxm
SylxZuxcuTGqaG8s3Hy3NsBoyLtAO0wDEIgHgy/FAIfrF6QO7AEuHer/ZU3ZW4hL
5EYj47UCPDjxHt/QuiypcuX6DOWb2kDx4YCwjsNMzrBD8IznZbU2REyK56aWyRPA
ano9lGr5QitN+9SbinkwEICEntgI4XrlNfREYanPNUG/znYO9qD4dm4tB5Q7gvHD
eacmPA06ImFAFhfhJQAG4r+zKqunVJOxBBQvWCxInrbpnxRdJQ7WePP7QkEYAp0k
UfwGZrFz1s6p0Z/m4r+z5746dY63+yuxGJWQfsQyVorvO/JJpbQQQNOGBJluYOxU
Pu2eZecc6M+xjjPy694ja0y305LOUZ2cm+Fyzk7SZoRtFjKlVeUofQwp30oE8N42
RKp2OXCrowcsm84v5V7xUMw94hI44o5p5CEnSjN7IQHbYQmc4pADc5vhdwAVsyyY
BWp/PBR0FliVfCtrAf+08yFkNWxMTQh5juPgJnYTLhjACTjM8dfjzc/5rj9g4V3A
v6P06Cbq+VFoiEp+tNDAza4j2fwil/wC31yzuu03y1yh2b1xUvQp9LNGevMcQ7Qo
axxupSw7gheyuOZYKwCikAeCFwSPSBDa/f2DkLZb2wGH/lOOEGkAgKWbda3M/6l+
z7RiEdhBXq3tVbhwiL8Adae8a0hb3uz4P5j7RSLO87QkQcNhJnCRkr8KrMOtZx8L
IrS+oEwAWKUT1w675EGs3oG/CYULDnNHzJGAviE/p9tDCzj6fxmmH0EzPvuQ49uf
2sN+JDOQz8+/iOIHGwv44+5U+aF1I6ex1d6heKooQP0t10vBuTn+0JJRSpspUY+C
U/Yo25A1tdLtMg+lPssRmrm1rN9SVunJ1wyWBflZlNtW0qiWlAKLzZcyRuIhZLFz
wDoJTaF+3i+Tra+6bSCBG9bBb7ZNntWxc+0b8h0q9Uua1gqGfLSWRKj3m65n0kI8
TnIjpjRAYLJlXWDCrPoKVdZS6HB7TAuOsYRSQYJjTOYfimshD5cWdKyvFRYC5mHG
glm2dfv6xKKWnvYXlT9Zza+XBcdgZduplxMKBknANZsKG01bPkvzqOYce/lbizA4
qes372CuK/tdN1vDypNBrfoHUgoQsC4jpuqVjHzLeM6gl6VrXu9k0Bmni+/dVvv8
4ctaw5GScXIievYtzzObwHUDMFU7K2iogPAXTa/NwrzJPJprEGpp5sdl4JJ06e6/
yAk3WWD6dcsI3QNUOsfJ4n1Rh3oYOx/EEExX06wKSko8HztXHuDhP4zcWbzOgguY
yvq/tvibwobVbj6BWtbPrQZsdorC5nqOsiEU1RzrR+sfnUTBSebmGNukytIEgaN6
G82AhiukqKTPTtPtYj6aHdePZIp7IeaLHY2Vc96s5JLr/bSUIz06c63fCcDx92zw
BVlcW6+BFUXwNbyKfyTaHoQ0oyHA69Y2eyIQSo7/pUP3zSaEzdED9v4zNs7PPTR/
/qbwwo5uPrjwDMljQzBepYZl8h4DhOK0qMBmvnkKnFBaNWyaL3nm83gZPljq7jUr
jcHtF6Mmq9Tp/jSUXP3+muFb1kMDfKtD4/m9dZ+YjrePQ9uWBBzNCezR6G3jn07T
qXmMsodSG3Jb5wuC+TYMmcoFH02NBTSPdcvg1JsFCMVp1BRMQMi4QpAHnAfW/aXK
8Pg27uJkb0UzFZLsaU70rUeGTxVAH+ZJZw6zGV0ugiARxLECnvOo9Al8Hjit8uKL
NrYf+iSulTKoplbyopIBNtO1MpSEB8buYoIFEcG80neUxvIqpD4Y/iWH+EFs45Jb
k5+3ld3X7pGzZW3njN760cJCBxWN6p6XkCFPj+3/PeFNUcQ1dabKjNxyGfZK69jm
07TfrOachfLz/hFYckdYBK003EkFS0EDSaYNGgjWcqTDicoJV+YElKDFPhdxH1zv
VR/r3iARZ7Tdryr/0blEnTrKI9wGlrzUqP1+dvNc1MP+VZOiFMKwmqvpVqK80DTy
Ddp2pjXC+upSXetlUCzcyKcDf/04Ve9vbho3cmlYD1TRRNAzK7hhAukiwIaE7y14
Trapl1H9vXcNS3WyFrEQnt8hD3IFl4Y6HFAKLk8ChwRgjfYBprbx3/rOCkQmRSze
ajaWWBvitPNuprFsNKdITKEaEOEqEK4j72pJGHa7PJdlLk1LSdzW7eFSpcYc8RgD
8p4Seb63w20W3Zy64cem2QzW/WKOhtmqlMToT2rcIn72+OhcD+LbM6ObGBbBHh5Y
W2g+JezAY416NhNebNsLgtuTB7ep+GsoswOaEdUMmJKlVMaONNtfEys8Z3ChVNuK
LkNTqoeeD+MT5C1RmDwMFa1mGHL8kqTws32iy7X3XASfUMUro5oc+jJey08fs4OM
KtGGYRDNihRzGiHw2/4YqsHOUEdPKzKopiqpMYy5Zy6INPJdRa8Xn2GbaC0VMnX/
YlMnT0hbBAtO+Rq9CT0OHWOYT1Z8SmVHkOgnwZA0UHphYkuAQK5dze7zK774BlKf
sVE3HiBhFdaLF7LmeSzJATmIy5cTBTho0b0L9H0i7/FgbIlqJ4du04fsLRAleLIk
U13owd/hD7vt2Cir3vbYkVc76/4aCd8afIk9DG1IqSMBakmj/putLz7jPm1YxVKX
I/c0bAVz0NJcUuj0AMLB21QLkgIoA2Ca0L+nCWHYmQ/JDCCVpRwwa5mEZpznW04z
bwCe8HwcZCFu09he00qo35FIfiZ6DYu+yzM030aoGdlnVwVzaOjFdKNQaR5+AqHj
y1Np1d5/bObQi+AKcptSCN8hAhgMfOOVRGVK9UpbBBUYvlfSsU3+j16zy4gAoZm3
t6Y1Yv19Z81hW003dv5ygYZn5NLb+5M40fMDiC9Dto3Am99JTZeWg2vB2VhbSMLy
N/74ArpIBWVbM8dvvy/2NIa9CzL2Withf7E5o3No0VZAds7k06iL0cJuT0HhikN1
7c8vDz/Y8K+sTBbtne47R0D7U53Xe7Nu9CtuREpxbZassiscsxAIgYzhmOGG1aB2
oEMsAkZ+KstmtFaRv6J2TExOnUML3EGbERUwstSIn+l84ijVt0tNoHSHQvTlJ/zs
p97YSq/ruWHSEPCR2fF7x19MsZMbjb6qKxFl/0LMRhYa+FU4aLOUDGcm1pLCOOng
HgW9FFyNN1nfJBpCD8gs6WIYSQaGVtdSrkIPZcvG6LYe+Y3WUl//9FabhplvlE4q
kVP4Ny59sySaxes5twsMfDfg0jnIprXw8z34uz65t8M4KLg39WXKrAu8Cr3sJEuP
Wf1v1d3KWr/SU+NtSuvxxltoM+Y/ey5jQ++1180IQ0h8ZlCrgZq+9Q6evbVdpj7n
PXGxBLG0ANntvt0W3EuIxm+rXHma4Whrs73i64MEfa6aaN/UC4jjztq2jiOEr0qa
Nbb1oq253LYRgIvO1tdFX+kfgyMomiYyaxnSxTdvsvz8AcAwxJZE15/GkodKWiHp
fZWjh9GnCuEVj4pGox+qbfunkwFLVbIRAvCuXgyyWgP23WvCSQLmEsQRUxqbD01e
qW5SjdZj/UADjdN5bbysTC2VAlFJEtWA2x8ogAFdijCPnt1mlcUun+GLcR5CqEb/
C4Y2EVIsQ2eoYot8B6X9QnsbANBb5i2swgS8F0N6BrGEvvDW3AGWzZwiILeQLxSK
BmA4XIpRblcAG/Uazu+G3XLCUPJYi1s5nW9L+TkiCASy8ac1XERPxiatogMYCh12
s8notZ0WnnQh3xeROJqLE0hFS/Yk0aoY/duEHh84N50iD+VglYMN6P9yOWuntLEb
g7MmZLq6wNitLHIJflrxJtGS6RX5ydNf9oE5LbE7m+hq2gDXywboAV8uLliyIDGz
h1Pz16MMrQrHXb4iV03zYwtRZQs8d4JVx1vgQcZr86dzCmzNCGb9JShvTFzKnWA/
KJ+hlHVNbXqril9794lj2NnA/sk6DaOmcJy8sQ8dsCuZq0crb8roViyK9eSZIbeX
kH3UIViEfKLNX8/g/I/V95eUeOIFmaQeICA5PrazA4yzvhiZqPW7ltTld43en3GQ
PYl/8NJDkdKwe55EwpVYQFFKvGNQco37hM0t7iBKM4gsNnbN0GOO9VX5m8f3+wVT
ZI7fUxKRaI0iplLLZM0j3B9LdmGr+51nNypE5tGnyqc9MMhEEvP6sg2B3DxdJscj
pp68cTOXjbcmJn3MV4BMxouo84A4Tk9xlj7DkaJNaN3fuFrTjZJTnwHWTGSC4U1D
mf7Kdhv6n2A+zO1JTVzwm/Ln7xroOGFXoUML+EqoItthHANKOkfDKiRQIpV0ULZw
abiHq/8L0agAArObyl26zMA4YEdTCAA2kqKN2wmaguHaZqvBcBL7UnQzXt8TBVxx
4JhWuRWx9YhSOUe0mNgfNKbq1H30QZM1Nmj4UPW1aUsObmYQ1Qf8c3upCda58KdK
ATDunbdfd3jgwIlesWHW6sOWc0h7eAHOdDHXCKCyyQkcbFOlIYR4kVofD67y33Ez
rFxQSPaRtcrxdeL7jyqXq8yGBcbMXapHrVw9Tu9Z2s7l8kqZ8/1WyIa2GqYILia7
nw02Y1T0k+Uql2H/XKQIGyDTZRkA915OUcNP3CN/7qgw7fNlk8ZO8E04UdMz5r+9
7Ua82jrp0sjR97cblIMup7M2QgPzeT/4ZdzPvSnxnoAJPQnpg17Urv7gXVxExTIO
x9ZEmGD/lP1+Ype2jEYwXQvS3X9UDsdRt6M8dcb1oiLGzM9UzRB/KQQHA8Nqg2Ro
kwb3k/uiLQvJW51ErzTrTyDX7WFHQ4RPUEnuG/41K6B6NNaADid+7Pe0f8LGqgMS
6CHAjnKp2sVxeI5WtKKKgYKyS571BBb09X+nFDUfBqTvAsr/PiAJkdroA26B/QMu
KOx3livBtGtHHRC3lLu21qVVcys4Y7yFB8IUjGPRrzyEgrYQQKcBIXjkZshP+led
iHu40o+1btJJz6zZgOTcYqK9QFTPL4yZ78cv8g8SfAAJGhTds4+MlHeUxVKXz71F
Ow81i6Rc7KwIWqP0rBYfDeRC/6lakvdgNZ7PqfZ3XB3vPHWU3HflAAMbX4a45WYl
hsjmCIoA0scR4a70ETdi6NO3ZvTUpVbCWixXbm+dNtNTmeMxhiAfK7vjscqbgKe9
qSpR4Z0+wYnnE2vD0ZUJG3C4Qx06dmZTLwYnBDDevXNnZdWHWAILHSbMG6Fg6Hlu
qjnXJFHySKBqgVdieRu1haxKjOxiXSSZWCxBEg+igNDGC1/04Tl5REs/HeNZX9BK
cD5XBmZnn/ujEiB30F1HoLumnVhvZhyKfONh6EzXNJfFZKge6sbRF+L59Zze7N0F
iXMo+ts4mfk6kMYEZzlHgqSOED6thdw4kfEi2VSNSJirJ0hW5euCPstsxiWM7JCN
w13Ju93+0iGT97NsHu9BPMCDEr8nMbuU6SPtSY6GcGXixoA4IgXPr1flvB9MIrVq
5C8Tr2rcQVAQ8APuxJriSSZBT16xLdvLuApEcULNe13Jbww42yNalV7IEKS4CKwa
gOhem/3qZeRLGOD1eJjtednoLk1lvgitDF7oJdfimFVF4Lj724c6/hrlRFSIFXUI
OAQr6+hI23gdNz/pfWsrQiY14doK5Ruhxs89AHVbwNgH71daLhu98tRfo3vo65+N
e+xv5TJWcXCzzhIBPYFviVdEdSJFwY7IVxWDcqP0UOryfWO2qmgXmnwL4/dGDUNA
bp6OcBGJq/n6LUS8tpg0UnXFC0lFdFXL7yWQXpOGryXm0Opl/HV3/mFZH9257l+i
5gSJ+rTgOahNEgQ3oU3sAU4HZLFzNgdM22JpHNWcaLdchHWBS2ky7HA+/mecAlOb
wqY//t24zhFhF3LmANME/qkkIgyxsieUHPTADdqmPkBRIx/CJYAjK8wk+n/uqrGb
XPSwzxWS4VLr/RSKx20cdkyyhm9+c5w9BrYldUSoekm5tM5D+BwRDtuPaPFBbXVI
1YrPsmxKlgIEi2VX2XLHclFtEpCn/cawcVYHowmQgAhbw4APDysWA3bNKHfaeIDA
MVEc/xFnzIJoBGoFRxQ4OYFcqxoMp5ur7E+Arark8mxZ9WY/tji0zywj3N4AQ4il
155xKzDXolfptBMRLWz73IOZ7EiYRhV3SpjLKZvc0/TYm9HvyTOyk2GSx3TW+jR/
/eMKh5J5Seq04JtjnJuFZutnGBb17XFNOKCeTQ/Xq4Dlc1WGHcEn7KSCd3wlNvf/
cKfL4DOxUfUYhMQ9cZVaEPvHcZe4LHQAtf+DqoGiZB+jZdV/Rs4iRwJunFVGM1Mm
IVAexFJ2GS7EY3AkPX/tNH3rlqgOVbQr4YaGg+aTB/A/Ct25QWdNAUhToXFLfVFv
fBNu8EfNxxbrq8lH7/fFumruPCi/ON/V4OABHzZpoC9y1AlNr7G8T3wrFCeb5S5F
vAQLDq4psVFgfPOrRdPRUFu/TO6R7uxIDsgeua/AHEYc3C9azqA5QazKBaw3747N
DC+q9wJ1jSmFsadpRnzKdHX/S7JXlmIU+MREWDRu1Rn4WroUPpsNs6bhkvH/qMTR
+OolZJBXtUrahOYW9JncyBCR0fb/dLkJ9qHP86g1sglkqiq89j9Lyz/1XKOr3n+Z
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nU5MREBP2v1Qc71LgZbg4AimEs6/2/NDIsZRpncN9XeD8ZMGSZ6MZhK/X9d/sBhQ
3Kks+rfbpVmZRtd5/qHs7oFYLpHRDbE/xMBb9PyDquV4CKSH0NfMcVbFABdOPLcX
RoVGOWJpRJXLWf30xBg8MTJEryTzgchvbix9+v8lpXj8NN5nm1CRDNzGT9qQnbqp
1l3T6oJesiNMCw+3KKTwUHyh3SmpgBEk9qGLyFdlQwQ4EcCelLCtKg2bzmJjW6it
RTR0Jt/vpLPN3GkHXGv7EBZDlD3sgD2FlBW4oSUxlW5kTqXufuIYgumIJXGjUBPT
zg3iVMRsxJR8Sic6fSXsNMokXXjjk6xKSw19Re99NOvu8elGAe8Tg/ySSebmOBfa
tbgaBUnpfaTnY/4xzXca7MpMhs6fBZU+vcesRPcMjZyzRkw/3MqvLsldPTnKtGKU
rTAc1p+oNj7WrDhdkGcXwWhuJ1U6qdS1bCjPjt+Q/5rNDDZVFKI4bV1PqPC4fAtq
CW90ex2MydGc99HH1xmLwVFp45eU+IfRloX3W2bgPFEN+ltexvKpT+lXZMQaQKEN
JbvE5CObRlpeHt4iqvZ0U4LhO7NWVtXJLneW1JYD3fhVdSdI/EdDmFtx+Pdq2n+O
wXgU0qStrNfXkWF54NoAeAhwu2hIAqaQA34OHVjR8YO3ZHPcFlk0+jr8NN0AS0aY
PH3Lb5P8IZxDLB+cijV2YO1w9raQA8y9b+ko95F9ojrt1xwSGV1T9shI2WfIHWGX
ibEfZq6ZRXn57b4P/voepm5qFr+Wj4bZuuJBmJ63hkcWmi9J+Y5rvB3D9yfErreB
YCxUqBug+0xwxWheZ/gJbTLB8+5NoxxjlJdkjbduhZlyfbVC5vhD6BoOW7NHHIjz
MsV9tyNf9Z7YwyFt1gnnM7mDUFT1HfAOhmZZDQkpYPmUfn2ptk2J+ub0st+YnJFU
QxZ8MAtV/ZHAXwtb/61pCWypbh2TdFkZ3fHhUIEa2w+XSIedA+KxBg4UnpIe544u
3Xz0BCYncUqnMTTOLhR4duowmEoN7aoZtHh16jlbg20Z1aMKoOAxebSSy77ZSvK2
yA38V79ESjr4WqRqGwgPZwfxj9uQ9rrf0AIWjToE5XpadsZLfUm96q7cw2Paamjx
bvJikj/c+3OVeucDAAjiUWn3IPbCR8us6uDyKW+guc+Cf6L9SdaLU5MM6+U4Nvub
pRLqGDtf0f43R31jSwDT3IQLezKR1IkGKNGCyNcc1lEP7OO1hmpLkabFWuAaWASO
iFegL2e2e8aBwc0y4+tjnbOXGnEwdzIeCJ3EipxRc+KMXLOdzK4BFQFfvz1ogHuk
oATg/kkIZMZhadijTylJoZ+HsV3YPEid3+Ll6PoXOiH2M5sXEFdX5tZtRMPP2RQX
VFscihJ4YjCAek0J5kT41SuqBoDlULkTSRcoTj7XMhXsEmjXNBH5m1lsJimHQhWD
dE6GxyRg64/QlLPzSnddB5slrWe9vajcRl40yEMZSezWBYhZvrZZ1EUNaYAMigE8
FIRk9Utsbag6BYOxGKv5AvDoEUQaHrf65AUHpGmtjqFsdmvm+uqGmoCCK8VYW0y4
+ZBtkLW4R8GmL2kML+ARkvrBD7M7qLhFcXJhM2mrB3OC0M+bUShigY+pLJ1DxOzi
uWaeJYsbbzV0cU9vYEqx/hsmijahqwRbgWs8AYxZQUYm/v+plG3aLmMTobBdzdki
tlsmCCvU59DoJ+NTWA1Q4tAXS0ousaXOjyzF46Z8Gi+/rqqmyYhxdwipw/9Vq8P6
+ZLUZxmLHkHybRV3RgP1FuChVeamLAA8kmGtgN5l9WSgatLOP2IK/vfs5Pe7tjt5
UYqOcutxXC/2CJgjvOUsgswh7ulM7jp1imIScVMWAJgY2oQC5UUoKJklfG3Xv/Da
QYPJekn3z8yxnEGeXTMmcsl6wXDG2FR8rcf9+EfHUMU8MSfgZwe+OLakWRckk/Yt
2sFE6Y5QjHLPgfrjJlIAKNxGhgj0Ipw4QZZamvH8xLSI22bYV4WO7alqL7G1kbnW
Y3PQ88pgQBpnbR9IZHqT/kE+ITIejf3rFT7CCLy+lcjKVcNIG4JI8tR2tOsjiiJz
0d+1d6jBAd1nnoMC5BAn1RpaCQJ97pVkwpFkxPpn3i9OKJhOg4NDuoyCLuOLgwtE
xz18MabREtq0uHTUBxK8cfPxOhEjoFcB12N+jaxSsufABtl8fMot+OYB0CO/AgNB
25SejhGOSrgV4hmKPZKfkybkZc12Kl/msdFPSXxdLdKF5ANfi5Obc0tE4DAzA1MW
Ou2dje5qwn4nkSz+g59KwkSzNiloFiQ0vyUBGh+UVVXmwV5X8Td3Ot2x7mcRkU9N
NEvw4xdp+RvLQaBv2NudnvEycgVxH9gXx+hyIJ9XmJTDydtHH2I7YXxZvfTdnED6
qDd0EZIn1/u6/lSl59G0hqYxttaGp5ODrwmcfcPwcyWTgguwxuWZoegrbj6QjEuI
72kdmtXKhTIt/dXFP8269I4MBiIRg/Jss5F4Dd4l2ebkNQtFHiOcv3uLvpdYGAHk
SOYdfBPS+QNBTALT3jKyFyBOn3ebPmPB63NSAqvDxV0pwSwr5pZEnKwkvTCZwISb
Dd+BsqYzg2j6gim6ETnXU2k3jlEmnmlRnCtH9YVKu6KYHqny0Te3xsQbKGKQ2hkp
mIgE3R3Vr/urDalQGl3zwTbV7vuRQGQRlIywapcGMmmp21C88dg8iHLqdfoSegP8
kPPvTr5K/faYphyxVg5NWugdTrCNHEefnSB9ps4498nrz0jI8XmFJQ5R34fTAl1D
qXTlE6WqenwxbW6A7OF0jLzmVuAwXHMXCX/hjJyQRZiB3vFegkyIyhTFHQKxJ0Jg
nSuNEapZ9OICfs6bPMvdIAA6jQjCyyaMqFqrp81KAs5SlALJJObeFENSW257hXAe
G6jQ+XXPhng/A3r5nsUpVUIgVITyYCmrw+x/rOyTvZgWfCHZol/yhfdJ//ReA4dy
r4DOcvzrULnYNgB93yloFhJwrg2aj7VYzSKE1Ue/gtl2G6a6okS+6/2SSrvtmKSw
M/b8q9AsEEPUyWLBD3B4Qa5Flvw0HAtEp4R7rydU8CVzQPIZsoeepqWLMQsQXk+B
pApL1tySSmD6re63mlR91eQK2qYi2Qscodf/ahXkNO1tcStgPYTPEdWJ0DAzrlbi
6qiYkNf2sZJQzEjVS3trX2cjAMhovEpsH7G+RGnn058uty5RFESmTS0hRWCTn9R6
eHI2BC5YVvt3VU53s1RA3AvzSTdwJqBE6MreHi5eSmP8v+xLLgqblOiGxrN5XsXO
PykXGZ8iJT89/P00loP9wf6v3GCtlL12999ocMI79m7h8L/Fra7ABjw3A4x12RBQ
xXmxV1EhHKhf7wpy8tTk8F+EVkRjb8ikP7TMyyP4EGpkru+1g1wsMyKAsMrZbNN5
RtF0WhnIEGxQ/E0K05GLrSLq6QbN2oKxolRZW35GvgvAGLNs6HyOpOU7caVQnWYw
Nr65svJegnOOZs7Pp001zPkpZqoQNMLEw7mkt9TJljbDXkV5lReOYBlNQVIca64s
5pLGQM8BOBXZBgo07Npv8Iyui9V221cCqZvgL8EUpMvOB4jclSeKZr/j9uXjRLQI
yy6aJjrWPX4Jn5COTT4aopBewWqx00Bo3vX5nUtbY+T0V+JkNEMGWItBpB1buqP4
ZFzW5YEjBbqMBnYVo/i0ciW0K4WA/3cV/bYRwypcwusxzPLvHO1YOK1mRUjW0m/h
jOTxDoGT+RlF7R8dEHjmciYJ38Roqkxsc+aJMHmtfFaVzcpO3mF8WAWaNO6U2soP
6Q0JcTUCWqBoLoGXNMcO3uXsr1KX6abA8xS5HRKH91MIlGN3LjHLWkjYnaWJqscB
P5/6ATPWgkh3PPUbUCSmdvIErNEihqm1foy84+b/2MqV5PJjqFDbh8PTOnu0wlGk
8MhmpV74cuIwDKbhemJDA7q8afYrE1ycNoDVtHryqwI=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htIm4rN7oAzR/KuMgC1zb3vh1ImDew6hgkC9ZUod/gBLvTju8I/0qfsZirL6O8lK
qPv9DdVb8ZxNBGe8h1ezWwEyjAoY5Ap4goWZxECHmPhLyUew/3frHCfIOK8sfgD5
2BP+wgMUQd5AGXNt98EYkkUphnVyME9esIIkqb6bZ3f60Z7gUxMMetkId3hxNj/d
F8HelZQ4ROIzLvHLSTuKkbaA4NSzSqVRAcHVPaDh2KENZfwBqxtwHVKzDfxs0hOW
cNc2PDtE0jWswC4IrrDNAcoy7P91PWoFFe5vr1/wGOoypnyeDro/mXvXI0k/K9oA
dpMW1CBqVyRG1NCiUn+uPau0m/pzhBOoCvW8w7RanB5WbZOWcO37Cai9UwIql2dk
RdkmDmcTZi4R06r8MFaxgHgdhDPQduGC4N//ZXCJB8loobIGgsMd0xV1rOPb+YvI
R5bbHNTBsA6fnN6+kBBUjaJUgFJ7FieuaLcBhbyrPdm4N1z8zewVY3w4vAegVEu1
pAidhwlCr1Ed/GY8C+HXtSb71gy6rAanqHXVrK7hha9BzmB4ieXaU/OdEkXa5Tgw
DHTffD/zAWINr02rdnFsnxZ2yO/uTYSLgrGF9sT2voMhwBNOTg/Oy+mzp9Nlqa/K
+yuBcpcKlDIK+GO8zXOJb9y76/shqEt//bOn/e4t2ud81TDmR/AAfzvnuw56yrNy
yFckk05U88u11Bfxm32LQJosPHLP7rT/7j7nIZRI0EAoN+PIR/uu1Y2ztke9aunq
/p26hcWSqtokTbxTubXmBolZ6qZyj1pU/ohro2ycm9nNqPVHPc6ID2z/FzTzSjlD
MlyUnpr7E4NCaIloxa1/slhAYUA3vh0gtDd+HCKGomsz+3Zi08zrxAaiXnbyDof2
+LDUc/fuo5mHv+312coj5kJu1gInL1BgzN8qhwKsm6F9GJb/W+VVAb/yk6VW4JHA
iPEMz5odvpC5l5pKsmQFdjapunWORGsHuZI2/rWmXrCQD5naRQZkmyb/nAiyJEkF
pMYcHrwxofiXrR8t/tu3DaKR9qp/pPKpgBCFkQQDT8D3ae+uIoObmeUPJZ58BH69
tO8kai0iXNqHsJJJ7st5fWfZCgYFk7BIUcUGBF42hbX3np1FfwNpMlWA71BsHDoT
nUYPjr+IRNxUjEnsyTMiKno/ezPmeWHoDnZlzdkevMRgUzMojD/smKwai9M7A0R7
7Trm4LdKK4cycnidEE7Qi5WcJj3ZXJ2qixub+m21cVQ9OaJUsWytPXNVzkk8EoLd
DjbCXCI7N1jc2PtIX9evQjrlMlq7XsUlQd2YDuvFvpitgP++wkcGwGkCcM/gEM6U
S+1CP1GxPfIHTZql2ema5xhOdMPPqGAZL0AJqX9cBIcok6d/4suT5cU2AxGCC/R5
bLJ7sZjijnqf/GV9CsmXQJHKxOQi4Yp6IwDlMvOH3vGbAW7LdfGWnhWzJ6fH0ceG
LwyVR72vHlu3AUmU6V49XWETEseQPLt4yUPtDREHdyGPf2WeF6VYumvU3hz05l4r
N9ZRPPttVrU0M8fsFYWzTS3snNIhlzWZBrHLhAir/Yf4QNTlEbO4kmBOqh8Jtmym
3LCRRDQNIjMYyC1I/GR/7v71ZR5fCyomDW6mb41gMXd1sBfzF+Y98dETiJJZ8Pks
EeAcGkTfDwD5yqxjA+UMmeDSw5DVwJA3rdDQorLjIrBQ5RBUJQkyXmNLtzOR0bcy
Fb9m7KGJYAp1KxMuBKCBeGEzL1CP/ytHbji8G5yPYQ89wq+iaqcA14hXat+78d3E
p0wiWOhscAaXbsZKUQugj1DblsptjViGegN4VVq+txFwjBHMaedPNpo+7OqH8KiK
jrrTkoLWsHE3yvPaiQaLzbFCTgAgmY27ZftackSuADR8URMwAoKrM8+nx065Uhn/
a8NZ7jwyAnB/TSlkTA5gLlrgaVhVjTBMkqj8315JJ617mN8eORu2diYvmt2GCZZz
yghlLSq7Q77RypQAeoflEXzqFvVubD2ziEsUQv8oiv64j3N9X832/sBEH5OhBtWj
TO83klmetmuOUM4wQM8yktLfpBtcTV3ZuPV1ulkuYh79p2tfBZhJGOvHE3RAQ/uF
0P1DNDW7p2eyVJGHDLOUrBZIxu1Wj2GFiZLvvBfhwds3fy3XfXREFKC7SsjOAh4k
apFakb04K7ABo3SyqF8xjLLFzC9qbyGdmzBr8XFWhglbSAf+2yKCXQKeaJTvvdEJ
1pOeTOxsiuOhBKxibeWoW/X9f7w+FnBX/k1DdhQ3RV7qXSdWR7OEZHh6RvP1ZKUb
Ajyyn0tNjd52C/saC9bS0ZBYU0uKdPdw/qyBstt/1v7cCvunpO+MYhNHW5hl+nav
7LJY4e1DBu8x7HZSY7S5CNPxb+e/urw6auyMwvpFgjE+stWDoXoKWn5bate5+Joh
MSeIStOT1i9B4YMAmb6lD4LRRFjoI1aPjaEvLDrwabepMaW7bO/9x3/zhv8s422x
TZEm4U40mlnoSuMoycGT6hnHoal1jLpvC2bZkJA+63q4BGymGXL7mYeGex5EQ7XW
yExn846r2fZvnok0BPO4be4RvJLSCGZwjDf7vvUyTQVRh7QgApGwEayIRqcIN3VB
COeu9cJJTJaOULOoYmNL0FeU1sK+eIxveMD6obxbMmmHfhP2Ij57rMaKal9rpqpS
Yu+XtDhzkqDo/Le2rdTTHJuYhX1wJNM9Ftyxn3GcOVzMMVFa2IOAX9MZ3kk26fFD
XK/Aufmdubhr6ONIy+XAtAc7QV04CyPkQzluXvPvDbAdgdQ/Gi92g2PoaOlvJbQW
9cAC6HYW0KbvmxZt5FHKjEF8udioQgGxRdrP5DXv00NcszPEGCNT2SHjYvj/2/R9
uhOa+W3wkovZOBjPWGcFR/CsOs87lB1jYkPL4hCg0sCc/WraJzogeavCnG4HUvtK
BLRKSeYVKT1XxOsam+rGbIo2YEUn3pwwRYMPxeThlC1ZWISzfyEwidsrQuB9rSA3
u9jXwmeDEICKo0kMSbcc/MepfYoWh/9yxlyD78r5VXqLQIXV2WIbFd0ZJBtAfAKA
ZO6950DDzRzUlyXtU1tt99IGag6SxCMmg0Ln/SDfNHz/RYkDdlfNTFZr257qJa9z
RBzjKRywADVy0rpcuFcHrKqNHiI7RjzvYolkD4wmgqXhGAipPFx+eqgYmjQaYos3
F9s1h6exLKUdI29f0tvXUrmVSvtF7yOz4TdK3QnMe6F96TVOCSID91w6j5zpT7fj
pjoleZQkOgVnp5XynTJttCXqC25zdfUZCY8C/+uVfu4H/XOjZM5cg5J9GWJFyyH7
KCWsPaIVcBV7m5ukmFYA3emFmOZXaa1OfPvTqF9czw9GyjEScgZaQ7vN7y+8otT7
9eTrlglNjiNWGgH13HWRlwlMqOPjutcmtWZkupPkkMMfjpwHfsNI503fzkGctfG1
Rz+WdxA45we4qtyb2wNhLnW2YB/nhW33VlA9fzh4mrN2Nx+Hy6Ju5nMaWbHfnIDK
QcaDVXvqt36UtdhB+s3q7ih1p6g7/ibGjnEMpGWiFmhxx3IHzWdrCuL+a5E1m5nN
gsIihF5zRhOAgOC66xzhFd3ULo3AxsnZ78Hx5bB3r6al7gPMNtmpUrj3IS8cerNT
YS/5ELZ42PpL6EB+B1DLIxWuz2kRjhIUbENZnphze6d9hbpKNDQpDAKqDnzRPnco
JTaFVP3RVtnN2rh7UonUdKILeYY0xO7lKLDCo2mAc892KSBqvhRx6WF3csp1sePi
f7YV97YniaqNPKhoYIyjuUvmngLWbROKS5vdIAq6AHN8CG7hqLgqDNdefIAWewSQ
yhOOmmDBHUKmp7LeHkMTkTWJ6SJrvz2Lgdvh+hKnLV9nMFQ3zCQZQKCPPv7ceGfg
vH+nDdm5YvjGQSBhX+i+OH4PsmwboSZCjZ5feRqUZnhepl+Gvvb+Z461MhVEh+kb
q5MPtwAtJM9tX6HIjsNGdwQUJyuA0NlXVI0+tsWAn7KOAU00C6s2NpAU3Xf7mWU7
H+J2U6MyOfTYeN2rTtd0jbK1nIeRvQRrXmjnS9ykeo1JjQDq8w3rRUpkkWxCr5N1
uBofUfNxUIv0yX3pNciJhojJPXRGc3kvwsQtrF7amYE9fJ7+aUoTk2F8DdtNjT8Q
M5YHW7AZfaDIIhTZLrEWhju6VA5NlO4gYGEushdxNzEFjgPcPOcOAOWxFQbHiNfG
wcmjj4XJtElO48MRFYDfNznv5IdKPrHp7IA8PS5PkKB9nvcQOTHW4MnYXdxWrHpX
/SpNzB8BKOe7nUtPZ8IxHVU2xJcd18uKCf4j58fzVorBrPwT5OyoJb9rJ8LNugqv
5TuCkMLu5f+Bb6S9yqmd+6FRDQEGJ9HfN4MCqQfRHMcDWU6IFL+eKH7HyqBMEZBp
vN88rQlVaLt1vfDF07urDcsw4aGqStOtC556wNHFWuSPTusSSOMwvIz5Df8fCmVN
2VzTEcRP7oKzreRMHmGZaL8S6lXaLHyxenoCRJhwIqyyiMw5KfGwNyktMMOk0U2G
pjV6oCeFBVmeH8YlLvovWgN8NQsS0PyX+YtIJaH3azEaMh+cZ0yxPeKv18uc9dHJ
6t2l6RAoa8YMlDmpqKgur4RqRXZ8UsvA5ZoxGXHyOK12JWz7C1y0rzbeAPxuKYUp
/4IO0T24D+GgNH/GD0y/U1hMxCYoCc4OjMv4DJxRANoMceMFVr3YzVw0HQjwZQRs
FswcdpE3Oqe8/kE4ukIry+Ax7J3kzLkdgcQH+YFGq08EwtfCknu7S+lmcBhZTi/4
i9PiejO7I7jFHxNxX0f1dGX6Fc1N4rNzPaYX5mGBLD3FNN9CpAdQni3BMOdPytAG
uRL7FB7bebr2NIq0aWobQDpI6nYO5zW7bQolnguQJWV6YZRhJDMc1TF5RUNIED+8
z9x5AUyxPMMYjy54d3zVTrv9bbv2PufYuETGAg9VtFCI3RYpkERzUPShwFQlExw5
XOFbcgLxOiIpZL+Kz17B8Jg4888KB7tSsmFN76VrVMvPYpaJrAunIwcqqYxnM19L
V96McnoixYoqWogwMTDS+rqkPfFW/ffAfVWTHiUvBFSevPnRV0GDw3elcVc1808Q
btbQ0bMobRil/Q246dWttijz5x7y2IIHQyICk/Nixofu4Dd/qyJzUCh1tI85lun3
yppor36UZqNmBx/a1GBwNCZUaZSAkfefeliA9yjfaxPWwRltXu5M3JS/DrU96JQm
CYgkK0SCKIVqxMWCfA40OPp8EgfqxQlTb6GPUbcrOM59ci9lOojWLLscmbbE//15
oixHYIkiuWghuYON6QPa87ne8vglRf1EfIlia83xCOB8MUWx9/0lIzYUO8zoJGOM
L4NyGnY09HiaXboOPTcywN5aauRnlP8g7K1zuW/GIVwYFFVNlyX8pQnXPZ89yPO7
RrJSlPVsh/MHMV5FVDN2SGPihNKjZMKZuf5PQ7jIr9WPrY4PGBoFFRLMsQ4ZgmEa
jfcP5bYUuj0lALTBFmG3XLs/7nXAG4c4n/i7A67XLMPBxbExqSKhXUZwn19Kzonc
6mB2XJk13r9/nO8fTl9RpZPs6c9StXnjGnqHWNfyoeW38y02fiQ7Gb9bOFao/R/e
uZi/g0kRQjPl8vTt7HTpQF2+X8b6Y1ohLGxi3CJjot0PB7wugGryhrgMxBeSve/4
5DdRUFJ3eTY93FLfwm8MD0p8H1HHm6nm93dKrksvMC41mrf23Ke5fctuIDt1H+Gk
LmeweYxOjsBoQWezIN/YQkSOVP6x62cKJlZ9f4/Jtynmc7xV3rquF0lhwTnWz3Dg
pyhu7jtvix6tbXCTyhXjymz51M24XB4XbeoZBVBI7oGwbQHwFVElSnWjIoLrAdTr
YBnYDVzuZ3K572HFnrvdgoYhkpSaN3CkzamBwAxgZVyvqahrYA8XSNlg/oaeSZul
4cFXEzrxxMlLuyp6yHJGdMTVxKm9V1RZx7ELVnZoXuyXli8nRSyhqHtZfOeS+5tX
ZXBRIM/JkL0SFNMsaeLR8gf85WVHch+nzdma5q/T/wbcIIQIO9zinVQHPAhAZKG8
zzIzJzOJ1jAR1lwDnNc06hmLI9Tm004nzwRHeMmt6MMVjPgU8KqwTod0DKlAYw4f
t4ihYl9lH+5fAeYyxAGWy+L7IbqE3flxLSfy0qgUMN7YVM655ZPRmP/n5exk+gs6
7Cy9FuuU3uTqCQYEvDpzQPlEAHa5HFeh6FMk4wb+gqk3ngbpFChPvl6RBkqBcRuy
rRecwukmhLMJtM3zmHI6Fav6X0SMVlTTcjBk/MZNaBzdqmNPClz/asNTO1m7h/pi
GKo4RqdnZom2oJUiln5jmHJ6wMVd2ylsUPGA97T50YQ8r4AAA+I72bwZqbJlxk1Y
/xZpdqrE/dFtfWH5I42oBAKSB6Tu1AE3shZf7kJmuLZ3xdEa2YmWHT6Y8eROOH9G
G3y+fHDylKJif/EEBrhMAQLQ95J+OqQkTiPhWtjhu3z1KX9avfc1it8A+zUSwhFW
NM/F2FYXHRTJxmgHueNGKGheX1Idew9kdftV0aL/8LxBDC7qjoBKyWlvbXzJiLz6
0nYOTZBNyP209wcTpnQqP1TZk/3wSBPp4Yt4DAwRe/k+jg7Yi+CbHGBpyrM00PTL
TmU8m3UdYutoPjvZ+V3E9YbHkdbEgofnYepXahG23vbp6oG/m0BKJPpQy/TStwlc
bXrbNcYzZ2WKOWHwR+p7vjXIPOm3vK8ulF0E0yxD0Y+BruCo6n6BtRavZiru5cDT
hveuqiGatfLG5Yf6o59jZFoOMmqQdW3eSqtbY2Dp1zwPBpYrQ5Mr1taS5zm3dbzA
A1Stzjq54vLegGCltArXjNRZS6PcOM1keVUY3e79Y16mzPPHCvdiySUAzWtKt5wj
+KFKW7aC1n/vWwhhaz4guEgR8EKCSMgbJ5JC/akHzwaSLuCRJzKb631l4JyybYwZ
aruB5S7vwXJpST0QTIRQeEo2TLay1/qMKO9YAb0+3K4oBVbzWQaNqoF76y9WunK6
tH489m7ngxEog2GS1e9fbMw9zw/bHY/MBAiX/pMZg9V3RMpSKndnkbQXesiJEDC9
e/tf/vbCMMis1fFiww8cPj//qeZoKcEtZnWBfyIYhM8KE6gSk9XiTrQfCXJtktuk
w8qnmN1ErFYSkStQIlpPtpUgQjlnKqrvSQXWm1vP6VdN020olQOFu3FKWBKXpCc5
qfOjPUofB8PM8DoYY2vH0kPfECgt4f5WNTuZIx5DwFhJsbL3UbBfJdDU4/BJeEkW
0MrOBIUBZPi27tzNCAjCXHgpes+mlG6cZQRGtJVIuaWsJEAp0evgz5dfghUyvGXV
uSPOLCuFky6HQfk3slCxqw/jRL+t5n4P2mn46ur54Htes2aklXhyqu4C3IGg9UMT
DGWl8OUilcsA1pnGxI4AY9UzTWkkdVuEEAUWM/ARombZRYtFR/fveKH79ND7o7HF
xb4ZAR7fgNrZji1t76hcIfYyUxfripz+BopzvCdijDNrOQv74Lh4qBKXvuljArmc
g536Pe4/cDikR1UM+QqWwkfw5NvAq4R5WwZWTIr/al9oiPA8JAwDuGqniX3MSGXI
AH6NKyddj6PXMKKOZgY27WKx4sbgN5VnwFkt1H2mzkZNqOhXcT2PShkC+zvb78kD
WpNTkJZRJcd7Gjn1gKD8mvPEAlvw12KPLPxS5YuscI50IzwDxDuZQToaO2CCQL9E
P5tUYiw42Y5JHYwa3DrCy4Hllp9r3eNZDIe/yBVs6UwYKZQAPsBCIjpD67OmEMxe
f8M7d5kLDzLX9gDHW0pljfQgvnO/RBy1ww1nfys9oDM=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4whXUBvJAPQR+1XEx9LkQz5C2cLsbs3EdZvPpipd85I4hInHJ/741PZH1hsM+L9
XqG4BTcEqmlumoxYQzTm2acquDXhZkPowW+gdZLaqOlbesxwHsrpbknONB68okxl
EWcGn/QKVtBxT7c8O7YIcEDiW0xi+mjKEl0+/EDy7yhSyDOb+iH5YAcPJ5K8iP77
YBg4cG6YdGGBLmHkL07BzRKb8MncWbkei1G3tIzQTzCXQnYYWPIZBZUZ9iJoSyIe
k8ktpqkSoGAW+aMg19uxaTX6pq2cMyDk165XyrKIlFIFefvq4Oilx+V0GuBruRG6
ufETQYZhbE6/z5WfqZzK9qx5bfgGxBZqjyApn3lmm4sJpppvVAl5jogPGoe7XmVM
ztn/QbbeNuWSUO+dUILFY6ETV8BM1E7DE01Lxl7W0ivJrQx09kbiOfHry8Kee2ON
1B9A6n6yuoArTJUB34TA4qrKqdrBakmOmaAqj4FGeH+6Cd6AnLsT4Frlex0nR+Iv
fLW7L28u7SbaB3kf/9PVAONfd/ipIA3DZ+navd8KR/+cNHCQ6+ZGQxD/tyWrnceb
oIHAo/w2S56F/mjs70WahL9wAEEnw8lf7UFEXk/rbAIralKj20wd8QW3c/FWyygh
6umtlqNIphGtRl6vdLlkoeQGqnu/sY4We9ABt3I5BB65iPVT/XVLBSVbeyagkJkY
qOMW72iV88BGjJpUk8bAkJd4ljICzgpqFXDDj6A79CbD0thM7mh64FL98x38KcNy
PT5IltaJELPzWaABMdE7yNfI55wsUCF8/wBnqgvgPcEn6ujcpVpzNH4pIflb03jD
Ms8Y4ht+Ni0y1oh1JywRuh8g2Nfi7Gw7jq9CydY/giS/B8ezkuVcLOJxwom6dgsG
hxaq2J9IB5L8kwpvEKJx9TLOLkbdqUpTBkRgmrkK8t5wnxB44ERBUdgfJKHCRhzb
O8NuHjwAjKDHWEMDlqW1PHqzl8SluBZrC55vBrU6euYMzC3ksH+SsjMFyQamkX+x
K/dur8iuoeKR7hA2I8dHbUTc8CkF/MAqQXW+09SfWXf0Bztrf/nVhP+uT2jUNW39
pUDGWBfhm1pCuwW70EPP5NAf5LU14O0PCS1mj/eXnSlvxD/mt3zlgtM2S30VXveT
o+CsiDMJF8YfL4p0EAcrH/RB87SYb3T6tXSVVQneiGTSY5ZoB2+aqLLqwCjfLvo+
jhhuATlZf57FC7KDOLVLjCKSf2Rxg5UKsf1Cn6nUY98KXm9qfqp4GdKJHTdm6KCh
Psbtb+Eviyn/Uy4L7RdiFodHe+4OkDZOsQFHFvQ4+Ks=
`protect END_PROTECTED

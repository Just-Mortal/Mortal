`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SotI5qdavsxi2VRpXXWhcCnQx2Ral+ciMWloVvMskpb1FXU7j5slzJN4eVgPATS4
6ct2WtScNaIOUJ4QI7PMhyG8gBETHtmM2TFurYt56oltpW57c2ff0mWdEJaZgtg3
fHLYRaO4TPXUln2Gl8pNyxQT25F1WEsiEVTC7BIk2ocl9ioUVMV+sD30U8/dfr+k
+rFXaqiJJUUNMytqcCKd9f2BbnQ1x/yK0oJzhGtH39XiJqTBbpDnWJa7LkZZAIu+
6/mVlqjiACQE/7EsiHgSSMhvIiNpfcmrh1XOBewThEXsXCWDEgt80ulqbu+MXb4O
mFRt/NRkIh8r8i+K7NKEoS1e/Rb2bgyoBtbdy5MZbWgAZVRa5+4KmXdqS2MwAOwx
PyJDllS7O0w0I8/dJlgmURX5eRyLJ4F1iZnX6ESwK2XqAZL3HI2xhqHpC+KwQnHD
7u1xVh2PpnnSkkhV/EXqYWIt/fxiEXOfq2TK3rUE10afarRatVGrGxey1Phhll3X
doZhSGmCsByiMpaX6PBBMcDDHxSsLHqXIK16UQBV1Ezo5On0kgpmRKGXAByjED+V
DXnvuKyyW64Wf4X0IQJIx5B76/6cMe9+sNFaQZwUFNdhowkph/HUMeRX3Pi9fhFV
u5nN300AJDYvrffmEU4CVy5Dk7/xw33SEKjW/x7rKU7VozDXTtSy1srMix/vMlHk
aWq69VZFLDEvEwQ/4hguSc3A//bKMZ8E4e39zx+b6Px7lzF0s5FzrjAxTA0DSHho
cMyEvUt8JrVFcM/23VIuX8PYoFRytYWbrgC8rzgdrb1v3iIqJtJ66kw7m1Imolr4
`protect END_PROTECTED

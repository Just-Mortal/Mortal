`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UISgD+3CRRqe4SVnijIHKwpMw47ZQeRibycSaYTnUGc39G9KpV9XxdW+VLWyj5gn
uKk3e9WEQ0eD8ON8CZ7kW4ggjRH99O5DC2g5cdYAPp+t7WQtIEzdOfV9s7tDLI0x
E7hvRaepRVyo8SU8cKnfSTYc5c1yQwxScZc5kgsRS6GA7nUKerjvaigj/p1ftfIe
Y+n8354qlKfk/cYkV/RuU1bW/Eq0bHkIphVuabxtom91OtR0hj4shEQwFX9Zx3pJ
6rtYSkPDjdE7goW+geukB11DkuGv0H/U7mCBSHXoJ//IXf+u7YDh+ykj0i3P1qZ4
HfmF7P1922HtYX/WRCUwKCTIwOLbm2bfuHd18WhtGvlpHQhGCuKyJ8BXfgDslk8O
TOHENF9vSs9C+MRrQNKg4rO+yq30f7M9iRWDvYSOrGXwcoKkUD3M3NETXMBA245g
jTRRQVIp6wL0HylN7bb7F7tFc/sVMQykFpvLqmG08eFlRfu5Juh/io6Gh6RHXQ1J
QnzeGRCEWKVL47KKP64E6k68C7RCAZKpyTIoM7BQbuKuCe1ra+lJnpVbq+ebtR2f
G49CTF86KE3ZPuIFrikVG/UFJTP3x51FSI6PbBZ3iz47pSJv/PGXUx/tgFUHsWwB
9p1fPmS+g1m1EjqqylYucH3Ynav0DtMK5gWka91ZKBGPIutLrMkqHAmozQKY1U98
RZLzWLJqZydEsYu17DXd5QqE4JDi0PhAvfCibfUn5P4Jaosf/67OWGdOln2R08pK
IiAITKbk8/9YUZFztOLjiL4jqAk4gDl977z2mlwDrg6ML6aPDrq/PPQdHp/QH/mv
w+M42XTcqnVtjZIwgbDizbQUb/fbXpKrEermftEp1InylDNEPaOXFAMTxr6zyknq
P1Oi7uBOHVdALhFxCNOdMye/LYfAyMVkWohYn0N0q5g1p0k0h2Bspuca2wr6uMOp
g1lkiBI7XgerJmZNQSgReSTSXXx97w9RvBaNiEnd7cUKlOyE6kuHlx23pVDfFT2w
FS3+1dvSrMGAIlIMflS6rHfxXe72vpAVYttGV8e7VZOPnZbMEgZXPwhnnMkhgeaj
RH6xdTGXq24tFV1USHajMqe/UmCMsSU+K6wRhmARS1bTW6yMsF3noFQj7NKX4+HE
WrgmwsddGzGPd4lks2UeOuLEePWjf0SAhA0t3cgOnYezv3Vl2B+aqYJcECpFMxv0
8QhFZ+uIrMvT1PF9NtcfyTwnbfwCHvNCcCS+eijBmvo=
`protect END_PROTECTED

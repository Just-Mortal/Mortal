`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aw57J55s3aAu9mYmlQQnTkO6XyZEOqlBqm07WcBb1pibdIiuzmxj8j0iNnqbIUJg
RlX9ARE1+SF2mVQ52AfhcNONJ0sllr16GtlnItuyssp7NTR298aPbrczpAzjdGfV
Gc+sEf+kSeGwPlgLVIWRitzqmpMelah0/Lie5UquDisXFU+NsL+j8hE8F9kN/c1k
qfXDw6dzR9DuKw00B+9+Pnot47KMYVXa27JxNi7L2enk1LjCNl9XBBlSC05OfSNc
43XUIxU1cIoy0/4HKphdQ8gj6i6VEFMWIUnC+AM5fAcHfWV56fAkvWwcnicNVvap
KyWPDKmMHmqfFFMYOfRdXN/8AiAL9cFZX50X+w9lPjtYD+6jRH96aZXmKOf5rERh
B+X7EZVZcZuq9t/Cu1d5SvHSEfO8w/tBb/N7f1WyVdn0viJRqby/Dfd7CDoxcoWS
thRiKj8rr6ID/aCTjTP5lOAXlVYZKSmmUkr+owNQFt1fCqgcXnPwQ6ekfWSMvGN3
ZLHBoEgSLTrV631g5ijmpF1ra8HuhWR8Ek5G+HlVmNS+1Xt7YHe6NtA5MQITz4IN
gjhqOZgv+PIy2hT5KpkSWVhoMIJRdq+wAG13Gdztevuf/OTEZcS8Cs+7k7AhqQBi
XsWttLs3HRROUPElH6mkZJVZTDG73N5dTkAEgknrGIKmBR3F42wk4a0zitWHvWWC
o5iTlXD86SKdYoSpMy663Os6MdewA+4llY6eyMjQyvwt20kL6vwb0HhUJ52co+u7
SQHPgfM4KXXT0BuPBlhDvF1wBup+JEtuMF6JOw652rU2GS4kjUGN7t7xnFK17HNq
Ym5IXxKvTRT6T33KZ0whPZ8r/Mlf/ctLNf15E2rMHZvNQUXccIEsawCJH/dgpHAF
1dmADQJdyLlZjsjB/b8Q7netOrbmds65fAIOXqDoz3MkpSReLZibfU3eYT5xQfEy
Kq4o306axQa1gx2LSWhoB8i2xSkWw5tEPsE9ZWZzPar1GwHLMCMT9Cyd1pVwQJnK
O/d8j4ZziB2PWsQ+aqYf2E0zu8IkrpJxNA9lO+PclN49nn3HRr72etvXCNQHpmpf
83d/uBjysVbqcw18l4NYzcgTp8e9BUcb/5g3ZQ2q3hd0YBRZb6SvfEh39mPbBI4T
HCwiAJYrvmM37fqQSl9+mz1MZyQ6mtqYV1MFdyfQRLPo9N4DA2s/vDCdBf6kzUgw
zJW78er0ERqzQkO6+Ar3nIZZp1M6dQVRhYhEDMr6xCBxzPoF1nxBuyg2sJbBHVR7
pcRnmqZFpmAJVxrlySNHUeeocquZCVUi/nQ6gefQmlAl2ip6DE/yE+KiHCyQMTjy
cdieDC2u43yq7A084JcfZajZ5996Cs9h5PDSJmVWJ5PXQcLVDvfMQcVXwQ+vKEuo
lxHEyfpXLwNKMZm3NsJHaKBLRKjf//hgivTxOjArvltueKawX8QSDw13V9xYRpHH
zNLZJ6lqetx9d6bw1MMGCD8mmawC3bMuqUehZW/acBpFliUNv69lLzdhH4jrogFi
5i58HQMieAlJemOaX7Pg5arBWYOnoNTAIIjjZtv6a5WPYL9+FGY7z6B2CvIfJf1s
EAbeQzcAKRFZ5njWZy/iOWSOhdZTSAhZ5OgbLCLb/xW58mJYQYqWGZhnTdhrMeof
KRve8PucOiaL9ozbRxI5GhqZgEAAR7suGOgLWDRLWgkipjJSLpHLdAjqeWgYbbbN
+YnCWFA7/jvsv6fRWI/0NXlEWROkBFPlK6NihbcDz3t9aWuPc5++TrpB9rvE78dY
DBMkDqgYFr/U4NkbgiO8px1b/iEgxZrOcspQFrqbZqA6Hd1qkhJzN1BPtl6sGSwE
CQ3RXMBwqfX4eKE+QCSGiGiWRmPDewIVCMe3BZeXKIGgw4nV4ytWmEUHUmMx/ZuL
V2yDswwAJ4n+9QpN01davlAVs7w6bRSLYc59Ni5Jyjsx7Ks8YzE0yWt3zLO8dSzx
jTkSUffGb3OPYmu2tOIlGpWhJZundSaC0kxJQQEfi6FyIZg2hLqRgg+SWmMt0SEt
FtwPmOkC9PCy6D4j99EUQ9erLRoumGhtOP6kxoMpWEsuKItOv47Y4e/nfXDU43Te
eY/TreCU69aQ2kVe2SHlsRE0S2bAAxYGVLIfgs7kB73ZMbPquJoySyQ0T8xTmVU1
5EuJ8Dka4V1sg0vUsLSriMnr9mka3sVGBSmBfxByjf9uJzMC1T6KDUm9uNFnzBDo
Eptzsriu5sY+yCn2BB8MQmMvmyewPyxe2XxtuijCsLmP56iCBi+O3rzcTzyZqQwe
o9T4w3E8YCx7ftia3LYsOA==
`protect END_PROTECTED

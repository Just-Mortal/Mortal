`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bAiDt3++ryosDNAaJBixcSXPmux4sFTPioKONRHtvajwFJp+vYBGIUDZPIKbSNEP
bnBbHJJnd5lCYMzIuGKfXsD/5aXnGiYAEaZkwvtm6c2HPhN8GPkKCMPh3DkRR6hM
1nDu0RTeRJTl/eMOlWyIdYoJSsZ5AmLH0+O8ApkqHIhnx7CdZSMfHfpD/kl2oks+
32DAvL55tuf8PnWlMGQU9JGkL9yz800vRbC6CRFS4mLVBhxlyp556P0drKa92IW4
+A0zcQj30vso59+Nle3qXx8WlwNfrnDI2HW1mI822CrHKiuI9GSiHvHQRsWd3qGJ
vvcBKfOxH9QBhBpXgJI+m/rJHLSVxixa5tfmxnPbCK51m+pIhi/Ozo8mGCj93euL
dZOiZL/T2gDC+zp4DWSLEkUcaKQpV0DiW+vSwtdWrlIA7QL5TIW9oWwLtAY7LEWp
2DaDwa7U+3vxezV3NNiib85BNAKRsirDpP7r2I+bPS2oq7JMjYQelCIBlBsQwP7n
FON6nlm0DkGxLGTxCwZKW4tW2WqdiO/ur+tQV6dG+Aj5M9IJMAyzikuYoQYGAN5d
z3p3LdGCcB1etVILe0meeHIhuDWTc4kZB+GR7JDSy64QeXuttNkeTP6JkRoqjipb
P15Lms9nCrDkLTEPg9khKOqPeAArmaSgAtGk2nFqiHiWbSUscDIbW2XzU0zUv64B
lmIvvNZjD65XL69Ifl7La+gm/cWS7egenxzDQIxvMwg9jTr5ZyK0TFQ54Y6Ws+Sh
nm0uEv33bx15UMZgqDjI8EiXZEhfjfDpysSE8yaeunlb9aoL2f/IEkLpAZ+7LAKT
IN1kWedqRUl1eets3L6ZrPoUtU6ffVS5GqwyX+WcpWwjcF2p5n1i5Y9KuZfOZHhK
7HbRqPEMozZaUZPy7FU87GCyK9fQGeS3hLCfy8m5lKXReEIBwJjXrw4qbQKNXEpD
VgfZYrhv84zCpLjcE97GKuY+dQf2UUj3zGxqW3M4zrJkyanC9LAwb8FAxH1f89mA
z2lqRsIgMnYrmJdxkEIh2S4ZvKGnoqNRbkA7k8wKC4SkftnnWwm88jEI7QHzsSdM
26kZ/8PD6UcDo8rlrePJO3f9EWZAwOyZgMTm8jzBv7XDrn6+edXAME09yKx61Zvo
z13VdRpWVitMbwNLeWNIOSmy+3kI+RtLFBvJn9TD53VTNyKw9EJj6BQIx159Gy/U
FjNH98d0roh8Pu7Ym1ZgxgUyK6mP8J4pcKSbwicJDH86YQImCE8wi5JdzZG+Lkma
7UkN8dcl+mG7l+saEGsFuOWCOGdwGe+RxZmXOwlNmqfoRVm59akGYNl0sjFyeuHU
kLya3q7rzumc/U8a0BQiGy4t3Gmve/zCUFoJmgOp0BI=
`protect END_PROTECTED

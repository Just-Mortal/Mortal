`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJo9O9uVrsM3XRsUIO49VDQowYO5qqg0PLOHR4mYxYImhLqarPw6tqt3KWVzccol
Q1ctjvXMiVdI0/tNM3uuh2kD/JCszQgiFHSbjMBn41VTomfsI8EMsFwv3otp1R79
E6Kasge94cuB4Sh9ql4IbhyyzArn3Opxh4jiDmZDOSFVP3omCjwuI4wcbWhD6UAj
8f1M5SO3/yIrFilUlzUjb+68P5gLU42v3KaGe8+0CTBa3A7dKCQ6hm9gv4hXcI1M
NVswfl8lckT99BgCqp1iM+FIMWGy/4m3nazCJuaeXShDMflgSyXvRMEmwoj/0R0U
38Ba9Qd1RQAXlC3HWQh0iOWZe3+LsnIj6OuHFYWHAmINs3ZtI3yZt6W8e6n90u08
Y4uxG8tOg5FipU9LByKX/TmdJqXWcFdQ/veTEZ4ZF8M0NIkb8vTnEDeQxzChw6bO
eYtj++VNBxjlmeHKwpbR0tHQ6eRqnZ91jgW5piD4C2DCiNJ1I6ZSCjuTd9ZIiuU7
OrWHnuE4GX2V80/0D4kG0gT3ooBYSmUEa/xAvFJI0BmepugvrtHxO7JcD+8XPZxI
nnfpNPYgm+oAqykk1/pzp9e7ZBkyRh9A1WAqITwNl3QPBlgEHLF7eto1LRJ0CCob
L2CeVAyasNzwPWfPkaDs8CpF7c9XUIpRHtk4htn7M1PRr99dwy5HaMmNPtpCN/jY
FzdWvLna1lg2YwFHf0CyTwv27O8kPL2Lj3umpnGnkiuUWApyoYBf3ebj+GBoNJnv
wtHBSBjUP7oVqKimVGLSi+8KXLflDFokrz7W9rr4wnAqkveakKb6i+wCYSCNm0r/
eqWbvOzjGCHmTOZMS2QOoFdKMGZpc8ZOwe+uucyglVUF72D26T8fTGYD2dipNWft
ccRUrzwE5qRymGdFl4ZbNBfY18dfazuh4R2cgwLFSj4uYIoTdszlQgq3VZIogjLY
XG7+X2iA94iFa3TpnAGJ3lvxv3rfJkxTWCAjw4XQ6pjj693ZAuhy3avZ3mbURwMO
VTMwrw099V6OGGspW7i3Kwgn9jOp/a/FBuXDEMBl54oY10BAnwLfQjha/AeQxtO1
TQqDBp47mjLlFT/QbsRTelB7EUFlx1+SnBg0EI1Ozslc3hRwnKPigSYPGFH4tF8d
Bj3q5X3u9Ft2Pz19SwXtBjUAlIqSRqy5eUoECqUG0yrKZ/xel+oIn8dwG6xuLyTx
XqWXMpK6mqrYyLDr51RmXAy6rIqNmrPE++oBcKFeiLrme/uZwMQhsPN+uN5me+U/
WJTyZxKjkmWG+GSpIsS5sGPRgzs/nVbdv75fXZYVHyYUmUB9aXoOv/NaDmuIG4SE
785zNr99Cp4BHezM5Bp37zS2ToBaYp9K898FPEa0eWFjrzLLD0Z/NQKazBufi3A7
cO+vFTYICL/5M+OIuL18eoh07RyddMGBuQ0rKV5FayRd3UL6TGAIW0ghs8+14o9B
JVZ6YF8MEr4JanDJCnyVak7feMcZfq33nrlzDf4+LigOF/9lybaROsY4uQPuMCIr
jeDGAMzi8x8l4px+05lTqMQoBTRcAcPoc5K3XzUkLvfLfEt6iC4iRpU/nnUC7gu+
Lb9WPKaZVTskJZfNv6AYwTdOBg0ImHwJzC92ZqwwSTJW59W6CJzIfbHFIPJCGSR+
LNS62MC06Kv5Ly2T7fGZulafW0twytBgKmLLCahiHea4CvR/i1pfLrap0qmSgKrp
rcG1+qZX+bfwvq680uC6gKBQfgqqdjKe/Hme1V7ambjLpsLEmGw9gbJnc1/+uiTM
Ed6XqgKt5H03bmc42LOANUdKD71R0kDZkozY+z1PimWUuTTmATurqgzod/oI98bd
Hf2vP2zzLeC1JKhowEJIwuI+4u/6cSmosKTUFpdvcvVpLipYMmGV2gZy9Q18Y6/u
dpWwWgsD9ZPnacg27K15wWMdHS4axKW03q6sJ7brk7DLI9an7aXv7tzsyzZBvJM4
27IGqtMfpFxPmlMEntgjHhsswdk05D7Hopt4HvbE5WHE7zHtna0JsfvybSnhZ0OB
8+0JhuaIr/+0pJ/2ZWiNwOIzjzhQD21ixNWasrk/MmGRc+LPAGZBBafwKWkTAEHC
4/XD6yMCLTT7dQ1xJq+Qo+WJ7C54TXLrSTWz7Put9pZ1yN0+B1/c8V3ylD3g+k/0
RdDoWBrJXAgvp6PlYOCIGr8aNLVYguG/7lfahLQD9TLj6UupscGlcztwGNzkaUvJ
kG9XqGVSqJyt6ugO9cN9bJhpXxEFW5uMmLE/ezRwiw2WLy0H4jiFsNkEVDjtZMa+
2UpfXfjuQanS3F8tjm39iB6hlOwGON7OR9sdZifrcbNSHW/vwaDfaCAJANviUYzW
iR/a8VC8EWqOZCcFvHJtGjvMo7WIEdN/RJEOLj6gyDUlSCxUdlZLSneUKKbRHuoj
51380pJBftUyFi22OW5+H8dCu60+M6FNf4ep02omnJEqb7BoNgS3X3hciMhioVDl
HtBdjWB75hVpTjd+Qn3j2f+ogOo022e7JaQXqX66MX57Sira/UEt7dKG8x2wQw9z
eIN2tkD8lqUBehaIXe60EYPezpxqx4yoKIi2xwt7qxm4CQohAKamjahZMbKvyfeB
szbLgbdHPrlTmLsfH/qHZmiu9zrOZINJnlop3HFqpFx+5ZjnYaDWveN6ODgd6YYl
ztZ5xtjyJllTJAOChS4g5IbADtwyDdEHpacawkDBPgxslI7rMAxuY++RGHPXrhs3
P0GW78+p0BqO+5vtfoqNbj8+4BCf4qjHCBwOKoKNVlNoynBqKtQmIte9B71z+NIE
qLA7hz+2Il9SrbFxW+Jd+3xtyAu5+oBe7+SExzgONpY4mSU/7XFgZzj88gSwMeFT
wXAqUV0Uj3weYMeY3p/opq7lxc8xOHTJiPf4qP7F1wqJXFsKD5hrDH8bl/Wb88rj
0ZgV6dNp2UZJOiYnf7vN96lnkgciiAwl9/oxw/ea8ru/j6eYcFbYwPGeB9AoG55g
0pBaPxBk9tJZTuL8WP/2pfQHw3pTGh23cj6KeFwmrS5/vSjk3MVw2unkpGqyIOHq
qvE8tsT8f6+noipNtDM9L3ueYOL6G+Xnp0bqyLU+YQQhhR6qP7p495IRpaPhLJ41
61j8uSabwrZPpuhIAeAKUS6dQp34EkGjaMvaDEROO7NITfOsINwofGclCnplKyXK
eBokfNTbDKox5TdrUWBn0/4x1Bb0S2YW3itArPRsW4h31QrNaAiq/sBZdAmyFW2x
U8GHPUYj/7srN9DIXMx5yue2BsW3ycqfOYUQiKoplLT8ShDcraR0CKy8YOEGXyGQ
1mfyw2zCjABQrWM3CjxzUWgakpswz8JN15Ydwu1+3lmBWGm2Z05yB+metfUoW5iH
L51/IifYjEbjSZ2CBuOXlnnqfP4GA3DaxjKPCe+VrLurGuYJCrlB/UzlbEduco/Q
q7AhRzTlhfusRvC7fOpsyKdT5HqqCOp/H4RQNL0L/Ps0M52TC7rSCO9pb+aMj77h
lJ1HDvYGReUrDA/GHXp3ZP5glrPQxI5i1e7JIspOnpDyzt29yRKlQe8A8KbkkZ4j
tW8IMspFxceQ4mlQeouAPFX84oUq5QfGWRBt3vVLTyw0go6Jc97QDRjkxN7tQ9ZG
Aq6eF7HQY0GEwmDr3DgCMcPQHrdrLefD7RqhePxQMMSwsmdsRiyN42IacaT8lde3
n3jajT9deewyLHGu59Io0sSGQgWBKX3l1aGC9Hn9a3s4dSPKPPeE/vQoBVmWdiOc
tH0MRkXTfFfVLo3xrYYXZ0Hk1uE/SrIwKE/+JaNj7y82c8zvlNLP9YbEh967kdsU
kK19om0WqeEYKqjGH1+VImnu5dVD0fwsZx5c1ZVlvuglW4C5EA7QZl+xYaT59GyS
YyNsb3O5YB1iBXfyZFeLcMfnah4Q5coVm3xDP9i3+dgkunL2XxAUZatHF3vjRg+f
UWc20Q97Z/ev2KcN1B3+QInT8Z+gK4IMqochxNCx8pZDtvEUYwvZQ+xwJrlKXjrZ
IhbXK24f0fIlEGuz73IykBxwI39Urd23N9VKL9vGx9ANaEZQVZDM6Y/8Dj3Nl8jq
bFwW3Hwt6NP8JwL38PSywjl9MoIBNL+H2pjNxTOhGRT8cfDFdbb3cvvfrXmdYfIG
8Floqdy0wqQcuGYhaG3N/qkiaF2H339Xz9z3qDXZ0m+Inocl0znv8XQo7Jtq4Sdk
QVLqbxkmWygmR8wQ8PcIMLxUHGhCkbtYNH3uIlYkL4LdGqTZebGf9lS9Aip+rNHk
zOVpHCctohN7KKwsiKXo0e0VV1yQF3hjIaKr9xMhG2FZ9fwxmxr9OTH5m8Ik45+z
gmBXy2r+azcarIPZ2JI+F2UOyqchKtSUyBrAx32SGhzTGQHHdv5WDmivN2JSg8Jm
GJnAamrcPzf0o8w6zLpYh4eo1wBu9vEBRPuOGKWbWRyApGso6qa9XI8F3R/PNIJg
xPDmE97LeiX9C/A73wj8nGciA94mn5XqtQsXsbgNnxgA2gn0za/FXidzmzJR7xhT
/Hwb+BDISy33hqVMgCD7e8aeXT1WXxV469PGHVLB3EYezDbd9JyC+86AIyCMJ60L
AQnzOGTeXNpeyIF+QSuwQpHsKrYxCyVfakHNN8fb0iCf848IJMXetpjOzjOr4HDp
/qnwJP5TyCLCDeK5/3N4zGzQzyjFXYT/gjKLduOCucVsWLvJ9MVawTMemdVzpv9m
XEFci8369K86EduzNgtIyellE9a4U+Fwy2m2dmV8h5yayaOc6K+8Mq1uBD1VdeYA
B/Q2lKnVTXE0sBAPfddMXsp9ToCDsHg3Kok18k+U0G2tpORC+mSnztUEC0q3go7B
yXJIQLTvDpsrtRWdWPJtAM0SortdbJ45yvDL/WX50MP2CL8oz/z6tZMNiGNVRN7e
vjUxupCZ9dYdqUR9tJjnrEs3Yc4Y9eUWnEeA/AZQq4YU9cqYqsORN5aJGMyqcOX6
0oq7NvdSFEF+1i/x+scoecuMu7zwHVSx4EHI1f8YgNwxAgVC8tbMkN95BCXgNQXg
YRDUxSq54Cgvc+aM7qAqEFkp5mo3oHpjmWgY4EGOMM9h/9Inndl0TVP3otlQQWrl
QBvUmFJERjkh+M61s7j6o0NzR7xR+r2/LpmRPs5a7XiE+f1mENRSRCrUoCD836/1
rGjwqLou+MlihyY9FJWFgBrJA5nIS76nbFyP0HNnDdtCeC5PjH34RNsMwnD5mVn+
jiJdPL6poF7uRUdBRYCGsvclPTddFQnyZb+CdhCJPSCBfAfttj3NuQxdH6w8GuhC
u0GW4xGG26NFVJc7/csoUzZB4f/rewNQr4t49cfNZ+U/hVGHs9eTrt1RydSUY5Nq
u7ROSQXCfierY4kWOrKrt1Aog8HT++6Dyj8bsureSs0krJRO29QzWcpjjGdoXuMT
bRq8qsBKlhQS8UbJhR9VBLw7s12I8A9Gj71zi5TqnZBcVVRSyDDfnU6mdMxS23IC
BbXg56T1k/W2ZkTrmRf/LD233+CH9ahl6439L/O3GLpc9mjdsDHBERx8AQ8RM3zP
Hfj8tQ4g7+syz182hy6CCIzP1IoMmkO5RQMKurL2j0hz+DxkXPQkbHbyKGA0RPjE
gdfJtEKNw13eLajP/dw0nqboS/T84K0yugaM8uaQ17Awl+7tGlmuf92ZBT33hOVm
9BZ7vQAolsSS+Pvspcu4NwLRNmiStAfeo3MZJTcMYBAN2kiu2XOCn02/rdaY/7Oh
KM7nh8ub9phB+lu36qMFrqPwgAxnPDbRxWHilT1msYNx/5yHt1PxYyP7UHrxuDov
0ExXdyYpSvCsVaa0oO87YYEfvU9MFNJ0WFRnavY+AHkybo6EOzmrPbE7Cn2jwcjd
SFRn7aK6toTNzMr/YSExyv24C2CrCyeD8VOYo8WmCaRaCIh3MIWxnUqBbWmS19Dp
XW2lpud+mUyltNyeUJ0MME01I0rTT98jVdeSx7KW+5aaiPTQCPDFwxr9RLYGgFRn
ImZzafdxaWAge2ExsUIH3R9OjmMlrQpuXxkaU0r7vlwKaagFhXDm2SI4wTpV+qcx
7fhtBWol4nrjTJvtduvbhcA/NZGp4V6RXIutkbRJkYYa6Ul1fUytfg03XuuUxO6N
9uiMC4Pi+g2B3pdId3s0JmatMmLKQE8kBUsnwuFDmBLJk/lm5MXg9Tdvee7fVZun
nVpXGOjL0DMlo8HkrpxsvxDIZrxLX0QGvSEzFn7z5RLypMfJWfvWKbAyuxWuh864
qjZB/WKfOjziTNg6T/jbMkSSvGnYRnFIUEbIn9Kkc9GuAwXxHAUGUgKG5DIGbImA
g2o72hLJE1BlQsLYYj4x859Kt9vtzcAsSeFTfcvTTRZLCYYLrYbOa/r2fFMY/X6l
+rLeIzbm9NqSZDGJNeyqdBNgs1idMErwmUpYXKMihPjVNDMyl/DaZ/nN1H6ff3Ul
WoHc9cCDBhULK4FBZYNHOpLZSo1Hvc/7jk1nnEJZTohMu5S0ctp2J5Yvl12+UgAW
Caii45YJQq0GFQXDQZgmiSi9LgLTfqIbDghMrId9upTDaQ4wVkuMG1bh52Q/U6ME
3eH5hny/0M0ZvZIXRxIUw+Wmdy3dvjjDybT6yfPGnB/nMGDraw18ialL5PXX8Wb/
7rnclOmS21cbaI71G59sY4xn8Pjj2EWAv9OfM+v9RHxdaugT/0CqfZcdM9AfD8vv
F4rMYBlNYMzJTXjuioxJCR82X/k1drOWOWabghViSpoZD2I9EDCN5BpnUkbc3iBm
RKBwgTydTsyjzgqohg/KTiStjZ4OcUkCXK9/pqjNHBCXX7zAHAkABAXlhcx5K2RI
DR8j0/AnWnIr6KwGU9aVwYGsABMwa8G2DRIVRKCebkL5cgzdd25H/LgcWjo46mTA
zJESXw8nLHxly7tzfDbj5OlT12O/OJFdilH7ponRyekHRU9Lc3GORvoi79nEupjx
eMP7LdkeLeVa9f0HthjbKederb1Zef6erEiW5Yxv99hdR/z5keYeyqLiVx8dBQLc
7dYt+7OAxvQXuidLb6ETlb/xNnjsJx0ZeGw+I1TIuod+ChuIFQ+UAm8fb4rNLEk6
10C6S6goCS0zZbgGZip3iPNliJGc4UveuS1zo2rxy25zzb1WB0LA8TpG/BF4z/bI
DGGBL9YqFBubjGx3ldvJsVyKw2932gD9wQ4qG4IrdVoo+asDQkdi8o5xtY9YSHfG
OfXmdo0oBopdgcVDoqv9z7AHVoNgWfQPdtE2GD5TyM9+W5HFpAepIS/BioDvWhUb
Rz1a/uGJdlx6JtP5YJ4yaq/JecyLvz4gu9xvNwsqUz4sRd5WY6YKHGb+6XkRZxsI
J3psyb0VH7XBHGTrkEqfucpDG08VJ3sUYFsWicK7rkM+axj8kvI++Xa0/ECrkCMM
VxNSPaNSJ7UMqu93A83bDKJPkzbsAH2NO/Ifl3sD1YkYcFp42RnPRMal32966NL4
FItgljKKalDshZ11RfpVWoIguPMusl9x0Q/BH2O8IpObGVik2KZKSRjUP3YrJ6lo
T+aY7py5S9tS8xVpWa10+asD+LOSMriFYAn5EFu2T8QH69ZlxzOpMKEX9GxoiEcT
qw0Z/LYHpeOy6Of+wLCD53i2MZNVEPu2O/fjjH0hFA3aAwaQrhDNnHnIovCpaB1b
GR5MX1tNslE9PFBIl2Kt6fimKA9OzIOkkJkZ0qbZH/hi3pJYGtK/kwLSP6oVAWRo
lMEQ1ncusgzNlSqXSw2CZb7f8woQo55OdKyhMspkyZVmnGGNKRgZbOSdxiTld6x3
sWVwhfR9bYcqaxfI29bgDz2vkN17nTQA3+h4f96fY8mHGzTURVTkgj5YpcsE6PDF
AiUhcS2qNyOTghHCWrOyJkaP73LnE5Jse+RciPc8BpEqxn/yEN1C57Z5FwBLXkJ2
n9BOTLRgjdsJS7OnkWzej8appGh00fR/xeoM8wQfGtiMZ8PUiR62REUah2jT5g6a
yXN8LuiIb5+BGm88F+1AmESziWng954QEifD+SLtK8B/q9H2wixySNZHvZuKFj/L
XB21JDNV3P9299wXTYAtK2g/OOGjXpVPgYh9TbF8hyeRrMvthGtQq6RAZAeczePA
rllXasS2R/QT7HaxbH9N0iI0BkDH8swPx1jhJmHCVunLjdBZulZBsOOBd5YADjLT
+iExmgSxK8V3+ThWFHfX4HixWiRKSs984to9gzhEgKHZYfDC35q7e/aCUvwxZvlc
xvyIUXVAiUVfKVDNhJhu7rMYX+uCUXv1ULnhCGnwzYIcSeGvHlNQgGRo+P+TOd/7
rX3SK7a4D2J3K4BH4DhFnN76TtZOJsg+j/ac+wxZ6RB6SYvR6RPbdSv/Q2rqWI0a
h/x0J3I4UvqiC0v6fjPrWh5JsqX/wv0m4UxgCeMS+yBtO0L8I517EZANJ76/ZaRR
CuWihZhYzYonCFt7XgyF7+HW53EWMUbkhk8HLMJqX7eqIgmCsqH2mCtappY9gevU
6Ct2cAqGLqAycFPoFkAUSObngqZ6fhtYD5+X5B5VXS8pyDS1w3Deu8agDEjkyK1J
Y1Nsmh7a6XcdSHMTttVyyiOkfxlvUbzpmWgHIZI/8Bpu0zMHZXBI5nYhkh6+3bFO
eP3zPPqv8fHbMIVDFfgusJJtqRkiHDrzLcLRICIXnIftpvOQqbeTljpPF6jkR/Md
L5BGh54wxOM4Z/ssiJ4L6DC/2dJjy8sj5sB26QMBQHODGFfRphufbZyTm4ksx87G
fb3CSpdyjYHh8RFWJ2SJk4ze0cJLo8JrdTHZwfNGnoAJ2JJw2YhkWmGDW1UOv/pJ
R4z7FYFy9j/++EjzUCFU95hUmYJtIcjB2KupTvY48il+0zt0hvEwOwveQvQ9TsY4
4eyC8wzGpspAoNBjOH4WXzUrbIXvt61QyU87uckxrE9YCgW3iQqjce4S4NHn8ALx
rr2tC7+Wqtdgyd2lv3Be9OAaINJP16BtXbjV2Flb4nZH9QJooAXbKCC58t7m9+N1
wj0GO9c8AHlxKi55ut3Cvab4H72b9C27EciiM3W2vObXgRPQhqyUOvsq5RXeHKsv
yonEwRxKQus6LzBrLSf8WSkgDmCUZ3ycWsTRgO+lpeGtzzYbxri2Sp3heLK1xOE7
qSKWArNmGoZgYWKnNVdMkWTGsm1xTKBh9Sa5ssIAaRuNwZWARZ+AcAMOrlZMQkyA
LysnNiEQUXiXkIjmaaicLd10abXd5ZWWg9pc645PAK02K6liPxih9adT2rgN2KxW
EmOnfo7Lz1x7LfQtOS5ATivjojezXvOZVUcQkE3f8bcBdtnauPJ/EDRLMpovi5co
2LRXxHJDYrPTC6pr5VBZbMtAPGAy+gJP5RwQB0qlYG5yARfBkpHwpvGmmeXv2CLq
hujmY7JZ4Pd8LoLlc2dgCd+P29HAueGDE9t2PXN7DoudWSFqJ5aaURCy8XmUdzSD
wAkXs/S+zkHfdJARnT8pkw/k9HPL7FOpXof1maaCNDPp7Yft/GinRj27FEqYnPBX
Wv3Cao7THVvplTOyaIkuksWwAdmgIzPn9uTu9f/ggH+o4CKR5hm2jHQWvEoTiHpH
76OM/ccDQhm9GeymGUXHvLARXrBZlaDe4nCvvEgPuyM2JaVYeyDzsDFCS+wOAasx
tISso9DsVC4w/iDAWeaHNl8P9eXKsRaThc7nT6a/XE/0juVeQx0Y/3CE/vGOlfWR
1TFLw0BTndDdog798cyM19bH6YfZPtp9vv8X7F8KNOuGlm7RCAMJrHY4vzQFw5yT
+J1KMYNh4/kB+jTOZjdbd38s7V6sqrwn6ts9SGOQEyZ9sg4LOdltF08taxu0/WWm
xOgs2nrT3waMR2RjeAUlMs1tT3xEQbc249I1TZUknVe+2fUK+Ue5dgL1dh3XVaeB
5cf/d2TH8hzfA4JmrttuXy6ws/OpZVWdm7gTiaJrWGiAPsDxDziqpPGTXRu9PDfp
fBm+405EQkDCvcS8ql+GpQpUdhcuDhlp3GH+ZRlBC0EHg4D9LVCnCvvfDy1X8U5v
LN0GYO8vkmV3I+mCS8HAhBtD4p5kJLsQfphDCYTIn+/kOzFYs+aX/uVaihq4HR6C
SY7hXolBalcalFSliYZdIqmloW9YAOPXC9wQd++zQVeN+x7/MfJqwN27/gAcfw68
O3E5hqlNQ922jh42/WJRzz9aRvtbaAhrQvNO14zOD23QFX0c5oMEO6YseT8turEF
OEI/WgEHKzOQM8Bpc05hMMms6AR9Y2AIzPovtMQkYv7ip9Dq6ZxtdeLp27N7+9dL
5DyHHtk2tVomAKmWLutiAdcH0v7Qipgo7rmoGsrhMv31RICGKdTjZJbZsndmWl9M
K63vivqOJrwJ8p74vV5DVtnUKFpUlNP0XpVJVcUjNkS67dHL+nR8tJrL6UTi/1mV
73f+/ZmsRuT9lzoBJ6m6lO0dEz9G2d7kyUPcNoTWLJ4EJ1QVvjarj+wFZ3r8BJ/H
4ht16oKEBU1+VVu9VNAkZaWmEe73QroeIhR1XbU5yvEvmnYJt7dIp63zB/UR+Y7W
7Wp8wMw8/rZTGJOatpQm96hzwwTLXANNXW3umrIcwSB4G8UHHrkr2pKCOXbmD1DG
KzfqgDnQYnJneXz43FWkJz9N6OAxRCbwSr11yWCfuBWOq8vx3V0ZRJq3Ly2MfAnH
9f7F43WOzbKgmUloP6+I1NlAW9VEhftG4sqVVBuEMH/8EBTQHQSmeWiLSImk/j7l
r3snJNZkV4pIQXpSJcGaXWjNLbFqxmyex9QL6r0bYP5JP1PWX0PEzp6Tf8+PBoxY
2+tyCSQZgx6cXJ2ITnVmgIkCFJiYde+ow10Yc/Jo4fykN3pq33S0l2oEUk7tHMBu
i2JO5JrxZV8dkvG2omOV/0KJTFTE8JaodGsC2Ky+W2zxMnfkqglmEZ6bzQQ9jsTf
vY3tMj++UWTg0rtf7febVZVukfLsbiTux3WKMuMMGtEASlm5aO9aGmx0O+cX08SB
RDzihox3x26GDssIAP/QUEXcN2hs201P3BCCIrdrWbz8i5jB8r7tRnlL1PlwDU16
6eGdkxcWqOKicM/5j1PELgjzC+H5MwKd/XHk3ijSoVoKAqecL2jr60zyiOg95wM1
vuTLwXlAB6QuDD/Mu1hZLabKPXmxk95+7mIjRonS/WBSFcI20zvPtcdeqDIyYg26
DOF2+WpPAJULTTSx1s8LjMjaNjX20/yyHUGD7NR0dyepGkiZrwPrh+VO3qvspxZI
bOCuUKReiB0hF3Zy6WQx/RqXX0kDeBw8W6QuxHh5OeHFuG/qoi8FVZ+iWh95L4bw
yx4KjF+5clRuM3/az4fjTULQnAt4l/rslQ8cM0zM/V9tiX4e+vieRbuMyiLGJa3M
lK6TWy2/xKyZo5G0Mi95STc9moHqR2LvAG2J8yjMPUGiAYuP9eUHgw+kuqRw1kKA
JImsWM7hxTQbUh9yqnVudzhMyQQu1Qf0UZ2Z3HH3hEqx6/R0H3cS3ZOtznKJMvCh
5E7+qjpHPQo0riFm7Gyj3JybOECju5KoO4PKTEOkg5HaG3zNog2eUBdyvlFPItKS
WX3Okm+2C7XiPKWz3z8eTL9KHcv7wk0648ASHVlUBBBGqMY/XdTTLVb3dTm5FSRB
K8XKSOLpOmTFuOmwM88iA989kR2EUvGpo68uqnQL29Dg0skTmIwZ4PdkehGdyJL7
J6F1gBva2Q859kjp5tZVIqFDfmFJWTQdSmhB7K2ai2FYYZRlGhKr4+BhbxYZWVhw
bpTimnrpRhJvThvMZheAncg/wtDvOfLGkGQfqQLoH9M7gas8b4a8fRK9J3y30GWD
HyU14aCdtVAyDfYY+hZHUhG9gw2WIJAn5TPW013LtmUI2Lw59d0yhXlSBn2nzxMJ
E1it+xyaqh3PXvNXHHwfK3oesfX14BHCmWNAR5ZgRBovcQeBiF3/EDcpPnTvwTZs
2USWyJcv9TGMnAd3rA5zxlNsDW6lJ2BpTWN7uJ/ZMZAXzSBxcPMtOWXfMb9rvm9c
PGNNdNZnRl7dR2DO4iCzbzlRhCNFf8N6qGZRjng38TBJxJt9n1NUFAqMRm483Rr4
zJr5GYkOlY2oLo/QGhKQiWMDmKhdBBUC84xZQnn7kF5kmcJNK1yCbkKx3hmKnAD4
W/ae+6TJUmbwn9yvRAZr5n3KIzMFga/6b0rv2wTYpAUzdlwSaQNT3ZCe3LLyg2eu
FLaHVtNOIaHa+U9dFoy/gTa5coXBTW7my+QEvx7gkgYStSOxS8hqoRZpVek6veLc
fnTFgP8ZQ/Tm+r5SpHEY9DGQoopHAJKYldCZwDQ4Q5/zzoWMnUt33TReE1ciWx+v
hqhgjI1vAhNyhMe/VJc+6MZDcVnz/lzezFu12VdgflvtI3r1t7hn1ptyyJ3HRJjv
yzcgtE/mcb+m+mg1DZaDSSsgIZcyrFua1WDUQSTqFALYoLwDJpA0fzwwQ1C0wHEy
2jQKz3dKi+/DNiOuhcaGRIksadLtSlGytrJr3tHrc7/i6cf0h7qrnLciSWLVO/O1
2qbgW2EAku7Y6XApWgB9e6OqQ0YkzaLi8Bugrc1lj82KcAzLOs8A/TNMktLuwPxQ
6ZWE0Pp/ssRHZ3HQElMjV+hWdfCyd92NXJr/07i5+Zt1cbb78szRQfRs+UQzBVOu
TL6BNy/Mkil+It/giJwMm4/PnQPXw5fOJKi3PzJfFj/6RyQ8j/xg/rsH/9N+1xK6
DnWIVFTAg6uwVV9A8Vc6WPXt/WVozrYIQDExwdBqC7tP7rfL1gX4xus3btRRWl0e
lkKwsTHd2g4Cpc/NT3yYlWMX7n3/OVZhNpeGxZQrzXlfpRlC/xZEn8xi8iJax3Rv
3PgOmDxYjonHN6o3imcgLue2O6c5/EXp19T6ZNmfPLhEqAi1CDhAOmuh85gIMaxi
v2dfXtaLR6fG/fjwOHxnFK09GtzGdjJzPtBqErhMqgQcSok6rlDQ5SM0liV0wtST
6MJq+bMHlcZWDe5+ojSQx+DT069kwUuROOjVdtrENf+9zc2g38dB3+9G0SCEiTy+
3kfFwzi2MM+7rYwF37+q6IqiFCaU87I2lyeMCItQQHsmydgx4EiuEzHzGmBtp0/S
/iPOzmGb8pPqNyAc/ZApvlEmwkO4bGIqpv4mgIv6psBzz7giVIslZoBUq1jpYAQv
ZDnuEn+X8SkvWEPlj6QKeoSHWO/8wXg+rjF/p5WAjmm9Sa3F6ax1guoHQ6fimrHu
xDuc+5hxv91sHdQ/fiYFVN5BtGVClnc/J5hlZAAum45qmaipc/XYlujNao8VrawW
CtO7vh2fTGrX6UEDxyNbRjFGMl0U0RyC6I7sgVv+Ddi5gk8PNAWJdb/fIDwlRejM
ka+7Mnm2swUiPJR2NMlQnGYaw/b531TI/QRLZFi2BNBp1+Yjx3MpU1pqpm1+TS70
j+nzxBXkcSoz5dcLrpD7pYeYLmEDeurhBbqr2Soh0xNiko2bCSuKU9BQRoSWcFGt
Fpodvp6g5KTJAumfCmXXwHRQyHvGsvpeYHkzfZ7g3QwQ7RbmsNA1aqiZgGpE1vjJ
PRxzpBJfsFEPC7biViY41wLT/t3mTN97BZ5Y5SgjIeP/qD+dZy/PXEtSYRe4kI/t
Js+XINy8bZ4Rg5hm+m2X3lMZNJXjT+77GnwGlXUvw7gZBgKiBhGC6rQwZmEng+d8
NNQ3CalzOsVmxVlLu0po8/lopbZZDkXxzDzhRYow2KnnzazA7F/kohGopNsi9FmO
DahzpFxnu0quZw7aqy8GxZY41jSpy8HfVPE8PhDU5PKH/z3Eumwfk4pHi5kaWmnF
ZMiTly6MxQhAU8AW8pYSbkxrQkYawhKvHJghoAXHY4DQ73VcTDzZMeOyJu4ydXzp
NflajRcpIqb+QKPYOB4PIl95ktF6NHoXA3KLJHIfHUJaUDdHy2GURW9NVUQc6/pU
hGLbXsaxMgEKuNX2/saYcHIOThb2FYhJN69OADL1S9vIrAtZoUJwf6EpgE8QSjtF
ojObietN/I5e408lefw/UOZw99A5qwZ/TCLkClKanBwXdPk5DLu622OMqpQFgCpV
UaErxnqGqPRChrjXv/rsZppInyMqXPgP8hE1kPMfYLJ97wdQDxnwWOyQzmJ1OYqJ
0vkoG9N0DBoHw1HkJgANlFDsILUxh1i1wik/pbQS5Vh8RaJCUEAh67s85albB+oC
u6sy8FnJnQtQg4Ihe1vIMvPq3PCSBwg1pzQjmtGupgfyhKXU9srr2feq9u79gg9c
TbRhPBcom680UrleFWGu2vSlHik+vqV8iynGF/vrLr89xBKYvcBQfcSTTHcoWs7y
x/ZZ/vu3r94rKRqtrk2neWvI3gSZ4vrEvxMKwMTd84oVk1vpSaCmJeKnA9vmjSPF
Li3Yf7IIzAuwPltiQ7TvQ/TQx6uZxW0a538IEMeQICeNYJ1HwkjFzwMAngIaod4u
82NNcKhdMu2u8XX8qXfYaFFJxCRqnFsuis+ATkjHDtapEz2j9/hMFd7Rvfjbsoy9
fHxpnrYROJnsanmMYZahSjDWbDZZ7h+MvCVkGng0IJxj6cb0adbNOgKKdZ6JZge7
CqaTzCUGyI4aDj8vKS9g0KT6SICanML+FFAbtVS33Z4pypsHaIZZMv0lK8QkR6Nz
vwp+4nttPcesRxN0lWwlMobFSuUzBLEw+myxKN2yZAHJxqEP/cBfmowwn0YhW3ho
WfEOcmbA1b3z3SpPTFnlPyh6xuXTj7H0dKtdZA9rdxR6nWkEScCqWS7mj1ZEOZl0
LD6UIrdwMycTiMF1DrVsiiFu7tHA21cnaGLoOaLOqs4Rxh+qr/7ef+klQ5og8NLF
fIDAyh1M1MBrndLxyZUDQapJR6SXwJmAWZ5pp2Qd/UAyVLWuJc3FfYk+D3nULZJz
vVfZ9O9JxIGrxU3TJoZe8aTevGesONg/4QwpaAY+Rmu8kGxQSR2c4DLBCI4RTOve
kUQ2DuxLVZyNdpKjZZn5iYbEOfvdHMH0SPzq1J1ZDdnoB9Xeo3nWtZLVX5kZAGZs
ZjXc2evyia+4xWA0tNv19V/yDuir0dO5WmlaLwDnQnAGttI3l0jEtEhrgSPQQbHE
DCa1F5hqxIIwilV5UXxr16l5bTIXldjVFeLXh/PY02848hycAM4WYO9uLN56B6a2
w+APtaSZ+tAcq3GJMUkcTAVcUFJQIUX1w4Kof4Ub5aSr/3yLvh0KYDWGFaWGrwaw
U3tkdye1YJabq/AyeeO37lDyEtRWhgLdgKEDXxZH2mYn9615XeaYxV2S7TjTzrL0
7CDXJsNCnb4V/1HcvwkklnOF4DyO5awtkwdD7FX0vK9FbjzX+N8ZkIO+iZ7//0js
dfpDEcHz74ovqElwcxTRCrPJhCbQIvZGLNU/b5vc428K2S+z6yIRnSwGaO3XJONK
sLEWQbSVNdZuPlAiVlWWdOuenri+ncT7NBSzGFsLVUJJAw/uLQPeXTKM3AzM6gWh
/0l15YgTST0ihYqWkeA9eGZjhPoX5iQA47GA2M/hWw6+SpNkIIL+OmjPm6xa0RyA
jO/a8WspOg8SH0rhoqoetbO7S7XcdqyaFlPcPdoAHSLkXgeKkN9sy+Jm4meCGjes
ttJHRibUtDBLW8NyHgNrWFFh5nzmithMX6FZYZvi6UaTFm5QmtCG2+w+yJAkB7rk
EZlayfOr9k25YY0pTnvXuwTSJ7Gp2Scg+I8ajU5VHH2CK1dOVNff4NroI6g82HKb
+JBNrudefxfcFJYlgVq1k1/rA96I9P8fDVNW16l1mLtRIHC0erxQBwpeRpDze7nK
s2ilh9h0Eis1PwaMjws7o9NCQcTNeoF28yWGRUU98abTxf9ZXdnMVDdIun4/WrKg
MSok9CN6ai7DJ7vkenFpr2cHrQFtTWhw4apOdhI4fc1Zj9Tb17t/3x5PNOlJ6+2d
SRNjXrmmxw27LRXeoewbdasm5+Qz//qTEYOWpIVDXzU80ixGpOu89FPU2Wt9Jx32
7SmEUFWzsiacslXD3TiJB1JpaRWtvZAATdSDfUCT+gwbeGj4AxiNU6sEnfNnExqA
KgntixWUA6JOQdUPqhKppp/RkuursfBiaqio1wBQ9RsY4R/ifxz24SL0ftKeTSZ5
vSP2gsxTrHigFwq+4FoyP7A6noHE6GDxwhgHdLEX17OTGr5oUzIEXKaPEgVurho5
L1TAfyId1FdCJqwhRvPKe/sWgND/RviH+jSzDGQ9BmDeo6agZWHZgVQB6+lvWdjs
KIQL3fDVGcGyvtdaS7Goim1OqSZtoLO7ZdgInxdsAlKKwXfJZ5bjvDKE517U3fRd
RMCCLMU+xbw4dd+I5T9TDBoa3UIa5j77uI4/cjNAHvpLEFe0QWIdiehdTVx1oKqe
nRzXSwYL7Cfi+NygLpgp/UzLl4TCqMrKXlsn23UJQ5sFfso9GxoaZMieshNTez13
2pvmqDtTGQj48nWiYfwlcqDPFDrFaJ5VrFSgn/b8sQp0ouSRPNE4uBZ4NLAEESQi
aQJPvjKHgGyedI9IIPbMrd2ZA/sj5RAtLdubpjg0ORMuq8HZxfimTsSP9dexq6xb
yEQFTDFKZ4atyME7H2/OKLO536OkIkTIRTkOKes78vmn+9Ipa6Y5ICll4SF+NT45
jGtMK6PUD91OgX1vRZXoUbtrZ4ReCRjSt946rkyJcpiGBB+cUtKm9aFl0s6iLmBg
U720CdMQ3yU2OhpAx6TekIGRfDof+T8NCN1NGJ2cZdTomelnpp9Wd59+wNNN3mX+
kcIklwjCh8r5msaS0L/Kahys07kfnCq0xOixKPr9YGQ2mECTm4U+lTggcVx9yt2q
65TkjdhBOkQnt8pLWKrKZQgfslfoPuYEUA6EYmoxj9j501B2YO5rwC1ZYls+g0kw
DIZHdme01SIRZcjrDjP7i7CEvqGlko/D5lWbLaWpPYyO8NHYq6h7HXD8kSIc1C8+
/HW5HCxGIFknB/hsjUm0Xg6Q+ghlbaLRfgR8CnMfCFWbQv5peiJEkV5E4q+Ve4KW
ilLNzIRPYhSZFXy8WPZhyAZsnsNp6Qse93UzBrrP511r5EUEc2c25WlDm/rpkL4w
DgGRUDQGR+hyhmPX+TMpg7vtwrk/vTrMP9ry6gnUaKRBvtuZhFzNqY2J4+fFoxxO
QTwxjP74H5cipUY9Ft80yE46YmE1CLI3eVJ2EC6qKt3SI8ZPDeiSYI9jQBeM+aQN
G7t0RDDtGXoRMoIj59kk522OFFHEl4ntR9l3TMNBIU+vFmYbOJnyYJ3SqHq5BLIK
d0UbmasTyelu0FL/ID0gRt7ghipz6YLG+8/AxktKIQ6RGVmOVJInu7tTBOSc0lYp
USy9o9OPcZYeIhKNh1iShJzet/6TngmGHlurJMXvEjDbIH2XYd/CL1Q+V93aeQnx
CTWBRAVQxQX9FJxKAt5YzmXJF1aXtlgaz0W+X3u5FeNyuzoDiDjtRj/JwAc+gEzN
BorZXnMc6X7ykQ7c2gwv9NJPkpkq3MzuYbYpSbUljounp7cFtvB+HaeEgoheVRK9
OlmkeY2oEGbNL4muA7yqv3lkw30A9QqDufWg+DPk1dHfC7u/+u47PeEglmoUqoHW
nl006pZu6xrjbPYdcjubzMREGMVhaZpsKo3l9mpfxJA2rKkcJ9mgk62ppr6PoV8t
79Nifsw+6+92qJEV4+iF+Tg1xhIGCHZ/tjWD1zxWMFWXNq48bjJ7CviehW/Bg3N6
oNCzeWG5CxadxyZj96IudYsiTzC/aR55oi5HGgufTZ6hYb7LnB/E6l8ZMubN2U8O
7xV/h3WLpv1NVBY17oMQmzcJrM3UgTCHjYv1/07szBOkT8Lvzct99vAUMjbYZBEP
/xfoLMtyqiyT4GngipkWNBwonY6PmU6weC14S5PgAQ8srJzu0IlFB7znYVF1/BIq
WdX1nH0lNqf+a/S/aDGl8kWFpgelIlUMYGPLOKS6diaL9Wztn2XyOIAbBMe8edqV
woWqt1w9j9AQm7f6Ds659yaRz0CkHTHHIhlFgu/8Fv1ZNrYAZm770DGRVUCIf0mH
EaFWNwZQ9ZdlvOr8C/g3UU6ReMJO5GlZxHHJE27w/NQQMn2JQUQ7qwGPctZsdoMu
9TIsKllk4CgnQPQM3TTe2ypnVhnWhffoze81q6StREoXy5Ri0x6xevco7Nn7/9mn
DuJSNN8xt3H6bWnoE5Mkqfq4kVm7yhIjL49t7mI8v8hSNdqEZbL9uNRRhc/+YloN
9QLsmepm6QszCl8zb8gxPmRx9dMTWCSfGEiBfSE5yoxYrN+6It6WiNTWe4j54yR4
elTbBuhS3/mDf4ABHv73GoYtD5GBcQbbGDpTsgO3hImb+kIyRCoXuzbf5e5Ae37D
Bo8e8tONf/Cmm/miittX0XKegHLIF2asQd1ukLXKrrlu1FS47SgxMtVyu+hUc1/J
xB8jgMoHQoafj6B9y0rRchvsdhi3bZi4mWXGAgc4SP2xoVmGS8rxdo8WS3e8efTG
Dltbvaj2rO1Hf1GLt7WXfub1FE3bsToBOznisUmANuQaLPxwANAEmsMSAwVWYbOD
U9u6snzRFeM9q2ZAamrmSv9ZlVaY3QxLyhNxI43eWsAUZGa/pP0X5TmOTzacl+wy
WNWcKJBLb0eDCxKBifmVRr80ZIFX+EtFE6thGuwPwEKZqyTeF0i4VdnLPQ/khP9G
PxPkQwtTYjdcfKBxOsmzR+Hhc3yuxS4vEH0QiT4kZA7SrCiKq5eqHkIXP/Iz9PjY
8M2MVQQN4dZ/39L/p8Du+ilxZeKy8L4AYZhaAdPHF7WVfCgJavLKjfcBGZScYEGf
pzmnw2w0qxd0W4BpSLd6sh0wW+bH17hA/9B3u9Jucj7FAKnuKOtl4w1a5lGDOcn8
cgI6uYbPIFrGRlsT1xLil+1XR4JGICnOpCFriyhzQ7pp264sIUTOnKDD3HhA7uGH
JOxQOo6Z0K42GXUM/lM/2IpIdbLzc3sJPEGrNKUop4StsLDs1VIPON0PLI19tl/b
WJYla0AG6jzcgZ0GQvFqS7kOOE+hFr36R2nFui1I/Rj0NqdCDiqHxfR7e5YqtJqw
e/G1rSUK1sJ/PfI3WcMAruvotuXdhjJHCqmRhfgjpRpxYqBkoS78yxDYLZRcF34y
d1HN+X84ltCUyF3AFR97F7G+vm6Rn8Xwk+vio9McR6YEkfAF5j+xdUhTEwOrkYzo
e33kagfp5mJ93M/Uy1O4+1LCxgE2Py1eWQ1giGeKH+TiHUS5YfXp6yg1f1qG0/LR
v+RavetbqvjU/1zSWAW1lL7dbfU/zvmHyVMmBNhz950/vSapnqCiQOS5xkPVX5GQ
EFcReJDx7eqb30rR7maa1YtUVApPn0hwlgtsrx2qhwkv6yq1lzlE6fcQUABPOMoh
/mB5e+DUxV+cLbOv1ATLV45z//p/I/vbIOClFl8QhPDlgYJFllZ/+lb4ucgHiJni
eFvSgqZ9ax7MVi6RGGLssoK4rD+x6Gr/53WEY3n123H/vBx0L9kpTh+Z3yEbtf/d
qCYPQ4Lp1pgD1HZQSU8Doaf3Q6FRub0tapqBGsNlAgoz/WUbDKYFR2XL+zymPLuk
bp8NdqmAK3npa93AlglrPgqV6gDqO6r7VeIMBPoBsJirtMk/8hRe466ocUk0M0X5
EsoX3IcQou6Cy4AF3q5UPw0uU6eO+Z95l5YimhoEa68tN/qzePXWoEPOLAI7MpPO
bNBBZhesdlvX4MedFl5f3FNVZN5AGMZwPd34570zCIwa1O6MtOBp2knAplS1uGwz
rZPWcjyqJbl+trtabIxXQBsbHbgOeQ05Umj8iHJczJpgkHxTOVBF1rtEbfu/yk8W
ek4Kmuhm3oFjg+RLlpgPuRVFi6EUHvEm4yVIA/u+VOPGD+u4vAJmMNzax4QFHF2h
YUxLYpHhtqRIu4Rju9/rItad4zqYcRCJY1Mrh9S6rpF0HECv4vktfV3PKPGVXEdJ
2jVA2oeYbkvMhrAh+YGhr2O7yYWMXhenkTwNfOD30CYrRlCER5kj87RtwR4NqNwX
zdW6DbqAPd+bzCFznOCPNjeRGhWjUR90S6K32WJaPDp7dnnaZorHyNm89AZzEdIx
qSUypRYDvSBHGfxVdWoDBtTs9A6E5HRUURQfvggRuaGZBxc36MKbLLavsgvaNAsR
AOvokk4et3HFw6fI/BE+V6ZnqP+N7014O+05GZibnpMkWUEMI2sxw0eqNkuj4wwg
kUs/G0TY+1+APOkHkUroG7K40DlBdHCD6CnIXmTWQRK5gf9Cnz5hPWXuPh9oMGaj
r3ndu9QDtcyFOea5du+FlbPyFjIpAWqP6ADyDviN1HDQY1jKM7aKyGUD8N5QCl03
bBgn6Lk4h32SRVfNO+cQIAlxEJ9n9pVZ4uRpxo831HV5g7FCbGk4RwFi2PjKFi80
4bA8gVDqYHtJqQsl9+pniVS9J4G7fgt9YaPZYGb3mWMF/68dZWKtDqUpohZ8Mnob
6yQw4zx+VQ4q2vBKIeh9EH9u9P1EHmKVmBDGj1xDLIMzF8KFvrDy7FxBq0D+MAA/
pk6FjFvCExNyN6z88Qmbd/ajd2NNDu6ieUyd0P5YJHatU4p+KK2X4TeVPNdTJjPg
e75pHrfUkAH1BG8u6AZyVuiTVrpOWH2j3M+qzY+Dr/szNYHbQ0cZXoHDsWYVqJom
g08dFv4DYa75Kgmf3nnU3v8JcS9ma7YXYPabK8n9gJLaIAsh75pHm2zwrRsNnibX
wzKjU8zOeTkAcZni7SwVaRYHQbhGmdBA887Petfq3ly3pIWQc4ZS6vPY+hFeM7iH
MH4AN3JO+/oHdP57ua3r/JNG6fgJMEDExlIo4f4XHZ2puGYo7ilDWZRTWKA7KKAG
Its5jmogVHl/0EmwRfeOQ+tSKE5VPm2jAKG6GEpvvUuFC+6vR2K6VjVMqTHoUy9+
GjPeu0y/s2TYqUTKVxamB0DX/RroEv9ENL+TzogJ5TW1JMXhsbiwY+sjTSOdDb0O
t2MDEHQi//Ch69nP3BPOr52pvusY59xTeLwhZWJCla9LaBL2oiFr6xS7M7lRSMLg
p2cuQKXrsz4nQbyPyr2zVYQL4nDxkNuJsfvDdXsBgfezDbP/7QUk+dBb2tQexpJg
IGA/LN0MQGzdFBycfvMs87JXB6ILNOwlq2AzwxaGMUcs5ShU/YjXhLhAuK6QUmy1
qy7JU54aHEezUDpIvbktflOISz3yMqmw7EpO4BBowuDKfucH/8mI/fOLB41ccNC4
NgvnY60XJDNF3qn31L9col7VKrnIZ4Rodxn1pWvS1aO6T52ZDl4kXrV6bpwIcrph
N2jDYlMxj8nre0DNFtfTMnXUN7O+6fWAWCc4nXyhdLu2WyJJ02jFhYFJGQM6WCCs
DjeKIg9mzB89nvzoVAmQ6uTgUm+MQK6ZVxanTw2sRVS4utlhyF9xhqGgZB3gE/xR
bQ4PJQv6PdHgzuGa8mwOYgULMHT+PgLW4fEa9bpRHht/6RH3aghhEk2e/oUB8JN4
pypHS2cCR5CZvcwBCi7IbuQai7v6DyLqSH7SicqJIVyE68paYCw7Lt73RZxpEAAD
BEk/3qz5Fo9FjCTtHn6BCoFbGd/aIZcWvrfXe9EkVxI6tzqO+UpPZPj2iqxBSWKs
m4+MmCI7YAqF500t/TdhP6LGeIivXQsA//RD3PcNNvDvrILEmq9nB/yrXI9VR01Q
dDO08T51ea72aD0Ls8FMkboa3TwBnlQO23qqhYCknVwzQowzeydJnssBO9YWsI0v
Cm/h7YnU8LKiiHQW6AZjgqoy7WOlmu3p/sodf4qAJaLPW1RsEaknAUzQYd8TseEE
UGuJ0a59UVve24ntXGQvR5YdLHP61qPRd5TgqOj+ynglg+lpu1geD8Vt7lkWk++0
+okpLftaAt8MqjJg7F7v/eZLxI/vE5MfSDxtmslJRmLoik9nHSK//sPk7iveAqHn
tNdKYquqBbbcAz2dFqdmG2kTsNbhps0MODa3DqKcH5L3nnq8x4/Dbi0/nV/YFJFM
D/lKUrKudvFfy2qz8+Vg2GPjP9KQLCmrkQkGqOGBwOLQnZU+iuZNX9pQFXFFORuY
7bKqt7DJJ9Nb6MwrlYI2iO9Uu/uYQP2RUzAH1QJyuLv/v6E4m3rZ+vfEMoquEk1l
XLC475jppgk0uN1CjNcPpPiguuNtgKXMO39K6zFmp9uZAyzRanKikB5+jCI7UhJt
3ufDwmlYN3fNcckXp6vYzRK0S9+bLEnnYDNNQBdhaor23Xf9a3QRMBviIo+gofQW
cUIclRISyH9VoMsP8C+kHHF58d3mZYfJ9pPywYfHgHnePIfiueYEIWXtoGsabrBT
/sOe7aKN4Xuie2jA8xB2O93vKRzCPGSp/pXoZNjdZEM0Mvmpz1NW+a/INDw3th7g
DVVuOC6EQSZ3tmv9TgOyKpg8/6WNdMMIsbHQ0xay2NuA4aS8OeMNblhR47csn/Fw
2Q7FAcUKWzKa+JTHjqRmKs/St/2rHZQTiz7bXDKATs2Ww0Ll9tS0g0AcX1spoFQb
JUlMkMMCAezYhvQJakupWvYDXhksc7ZtWX8Y/gyFWN5k2FM3bEDg4NxB0cNQGzNO
2033h9eExILu3jLkN/FXttWo3B0QzZRWS9msuXJOrBfiAVwSYZexM+jdTowuwkYB
EhdVtxHK+DJ2WM1GesjL6XB5LgwPNUD5lWx3OSrXrTYYgt0euVSLLwjKPathc9Er
tmfliF1K7zFfHHfNLHUwhDxTOsZSAFDwSOwlTf7M7MTl7NulwAVtEDtswbngzMj0
Sy7dGm1fahOnnpEn6bRNLfHMgHUIUwnMZwIdJ5pCEMEDz1btihEhlMG3/A4YDeN0
li3XjKucbK4MONxiT+UV7Z5icrffYw1admZvqsKG8HfOS9nVQY0ev5ac2MRCm0Ru
UIzXC+SEBri59GAHF7EVMn87593cqKQBGVGbBzI8HSeBsScZsCq6tbWEoDWek6kQ
cz/ZLx5oWvg918DK+QAX4+DoL3TRWu890nGzkBhKh8tixy5ceiPIFoUj7q/ux5fV
nykFG0iUs8T9P+Bkg6yPUpaKYsM4rWURYjOaL+iTxkly2awHSSUML7E5KzxwfkA3
FmI+IF4uqbmADCmDI+g4QXnNWw02h1wo/iYSPIWxBkVYa3762nASyLz5KrAdiaa5
eZe9nCacZ9vpTlUIflEdiDX4vdkQ9lELuqznnBIfTh+GY4jYOMz5DP8VEVeVvTp1
l4eOe8m3OpYuUP9llViKAcxtwU7dk03Id+gh1RnVu22HOxm9jP/9Fk8HlPEy/99e
AGhDcIFlApGBMy0i0VWqqkMwTHvWsJ2VggFVoyaqA30AmMegZofrBR7M0BMJqmbJ
gi6tOFPtUH7aUw0Kyf5HMVGvTjsRfVz/7lrejbanyZhHvOVMB4GClseJdhPhZusy
23NZpdaaQrAC98rP3jmw0RqiQ2Q3Thrtmz/Pu3CFpdjVWDAzOOLWe18gzvf6/baL
VvLWFqIMp34BqYtRX6drFYRY8LD+7ThPyOYkovIWNMqC5vGV3cDy229rUOAddcKB
2pl1u+PaWct0skFgc+LT8p1oWdVy1Vri5AiyHY2ncG/PBvOnHQU707Bszw11W19M
s8CKAvi3l1eroUsSAvkUW5SHqpc20UN9wY8lrosVZmsx5HoQiW/MZSgyDH5cGBWX
m4Tq7kqmcInDQEIA+b+QlRzmgLhihGTLM6DO0y/oq71UKted4RiegMRXtTUMmTnC
01piXKWby5N2zE5IIZIjdrnlqvKHXwhv2+J5a3G0BR4T8rZhT3WfwEJmxPdAJSIs
4iBfKWNi+LY4KTx67JAA0WkMZuhv3jFMHMIf6BAbJao0OBuYm4FU4JirCVoHTIZe
SLheG6mzOI0/ovAqqSOCR0431fZFgpEMt7J1zD73USVtAkoMDMFvcM2H52x6KRbG
H0xQsVpJ5Nj871PJ9Yd4WnIIJizxgTNW6sMEA49V2QaFbFYnWP5w/ThUYDbqHOPg
OGAViIq4GY0iAgcS7QwuPtdPfLI0iVDn+F3yEGCdN5LeHkmtzty0Xy8woZT4TT/E
DhWu4R8W062ulbMYqT1gyJ8dopwTP2214vR4aMwyBGgUTPLkdOcp8VyjAhRczq0k
wQL7+UiPUvGIHE7HlrDnJzD+lhjm4Hs7JSAa9s0pzIevny4iAAQ2PcUQRIwSzFPJ
NtKZGbznt/2qV2L+DPen/rgqkGqrJ5mmByyNFRbRY5NvR6405YBpbm1+jKvPYsdn
SgXqeb+IRK2NI0mRUKeZpBQOs6YpsAWcqF/edOSETOVfgDuOdAZIYO3jtv5DPJ7u
KO8SiSIV+xOJ/9zqaPXza852cRwuiZkykHgzSZPW6OmQprVclf/vwzqF+yFCcNYw
6A3iG1N+vr3uFk1q0Q0KUOeVlLgd3xzicCEqy0JKbal3QC2jBJRdRUqfhhV+8M5w
cRJQ/CdHF5Pu1qf1CzXI/9eRRdKfUjW5zTbjhKiK8NfhlqMs+7r3WGA5MiWlHTQw
5CjJH+pgrDYARuJ4waaU5NgjN9cKgZY4N6u5HW2TsS//f5UUAGM1BYOIfWbapJw3
lhVSoFSMD9KtHVZXmrV7/IMfpvgnEr1PcbHeQyrpByKaz6kM1kotj4dYFFXCq7+u
lPoETxypvR7TI5sJobfrrLLwd8XNkAqhdodSOsTdocoUXJclTNamkPtNoU0AdVCj
Nhtg9GXT3c/R1GCSsJKyBDbl0e78P18OOBwpxpguea5gePL/k5Y5KVOwCx6BjdwG
b2/PTYfrVLB+unpvqVq7hvFQyqxP4eLSACWm9RB1N5fbcw9ESIO+bjBQr+4DLvW4
/5FVvWkmRn9ZasDLTBSG5ECLQP1jHcpG9/Y7QkKGcWBtU2XVYWLjT/m/PllhBWh+
uzRWAKom2e8if6Ga7r9yBMfrl++xhSiRidZKdcvVG24MWFOcaOaxIXgOpfHPYes4
RF40eLBtWY2Js+zN8bo2cLfBz6Jlqb2dgZV9JjYLs8IBNsocO2HVvPbkGxlpdklq
3E919A9O19ZnKKhRpf7FBzaZKJz2Hc5GtJZeEKXafM6diHIbVtDS7fg60ylbIncF
a1mPApUGVn2h7oWc0EzrOOOaIKX79VHimJCdtFVizunKyoU1VU4Conf6R9bx/qkL
Xgi83Tz6oQo7bfBlJCfVU4JahTmQsGlJT2vjgZYrIUSxDBN3lCIy2hjLDpKemC1v
lWHrckTe/SP8uvKJDrtXwtwMZ4929m3G7T/qqvTqAIkX6KWk5Ut69okwM4dnKRWW
MeDHNvvhJjGJ+J9i+ynb9ZUg50f4mmHrRrBg8etpsgEU92TkolgNRXpq5uI3ZIUd
2QWZIFiVy7JzUCsWdNTGtqGnkx5OamON+mSot2xLFg77odt6K5DxJdjo056emNTF
ntuRMzKyuKGC8lNBVXLuyyjgd+sHyl7AdW2kVX/SJcdfeT/gbSozI9VnXDmk4gcc
Z3JjqF2UBkj1DawTEwO93+/mGuqefMoH04qRrAsXG7qLXe3ky2i87lGundGxzRjo
v6AAQ72xMqF2SvJ0nuVYmBfGD5nxAa/HBLZnPWFzCySuZUXi7A9eiDYZC33bydqJ
jFJ/fVmJBgKBz28NBCQVvxq0qXhedYecA7LXr3nXBwChkmJtSh5qvpSYGMtxeJBM
WHUIRpLkV6w5mIjH1p94JZ4bQoJjwPkZE9z2402vFsbCDPg5KCLscQaeyL8g2tDu
hZoY46raryfj/fZDDoEnch8QQP8hOWQ40OSS4Dref7RqSsMydRqIihptEjgPOadR
sN5QQHXNhcmtBbFiaj2nozIC8xOu1mnMlioXpiA5kRwjqZDMBBeOFvUfh5o7eM7O
PVlXxjsZAn8mTB+HgwFi8J8NvJaAhn9SM7mRJBQGrhgvicX9vebWD9cLLiL90sjt
dfeHXzge/VrJlzBigkH5GKUoEcal0d1lOXcOP9APVBZ/GACgk45Y9u6fKXu+DEGE
oyqTh5mVYiRm6mydwmuawO67mF4gbKr1MbcIJYK4BCzArdurWqWtvTjUxzKPoGiK
Lh/SbViAt4KkSYWnWmzwXcIrlDORIPplqOGqqpOuiNlD8+snACUJX5eCEr4MCNdk
UM0xzeYzFlF+p3ORIcdGFVPa8v/QWGHUQfMPmUFpf4ZEydSyh+HTNK4drmq/0Qbf
26+/CcQkuIoSzFZpPf8LZJgKrgiej5dhppW9zoTJwLBza946YUyjuh9VxbXtS5Xj
zUvJIxzz84TzQ2wc87i6aNhqX2eJnWLTb6kKr5BxWkX0Cg4hkvu4mTFGspVRY8oK
plTZ7m54QwqDXttHSIYJoYdLsQLwVEUQcN9bsoQHqvkWmC0uhq4Bl6h70Ww4qUl+
LSezycNVaaQfm7q64RuYQjo6PdkDcSnFP8fiFXLrqcecho2RvDTWliaX/oAZml0q
KtvS1O4P6TFMnVpuSlYW+bkHblD0Vmc7NCRlyxIDNmEL5rKSFYe2gr8a85uxB3ec
gO6EyUDwxJ5/a2T0J0aNPBN0UInIbRg1bqsIT5X4MbBzPUYZ2UhZQG7T0IRz5AIe
G0g+hgqN7qezs3b+WY/mu6to8RT8p9iAAcKNwqkQejZiLp/py53DC4wEnFhCnjVJ
h9Dk89/zGmtagLKsct7KcWhjhCPTFM6h363ktUUpt5dFwW+rmBJFHalyOKowZ6AX
z4d/O14eeFTwn2G/+qbYGGyIQ+sn1qnroaemi7feJpNMmllvS0dP1O+6jGlEYy8U
OtWkvB8BV06VtDWpzRbO7kuO6xgj5XSpTAKJI+tgnPByR72xuBpnVTu7ODuKwD4n
llK2al76SiOHmp8ItOzAHprZZoc3PnO2fY0lLTnHM5C1e3GHcSjqigICky3YYu5+
QRlJ9EKXfvGWVkbXV7uAgiKG4avPAU3HRSD2nTqHB8CRbXlpqRwbVH+WQIcqBPNf
LM28J7QZLMCXP1ukxoT8YnS5KQazOH9AyB1TbkiUGJU+aEM1XYPKVG2rALp7qZrL
GUcDuKIaybNUHzUgbXIxM14fjH1v9BQrktZUeqHEJVqKllSYSBxU1umbbNlszU9v
2yYoP+cBt3V+rqdKmJnKOSkvIuN4IoJtIbHDkIZdQthXcidUt9AlXxIC1Fz6lrwh
a9VksLSKzkiqHfwdtMgG2lIAFrPgSwwVTkccDXL/70Rd0NsP1uVyeKjEPBAO7o5C
z5NzhE7RE+ojix09ytVYrgG2UP0a/DHHSnrNfobu2bXFSFdA4swauoRbbgtbfEuq
YFnoTDDDcB7WGeDNH18uHO7yo1L8jX5ET22YqlHiAzz7fiKJiYac+0KfIBL0WXNY
0ZnHml3LOeyNLltRUjNUaV17Z9JN8nYmTTer/UG69q/O5d4NwJmz0jZoJ/OcjSim
weCe2+zYsWKJ5F06EiDXmSiMdqfhDamIaUW7sVMe2hs38mNjVcMF9JEx/Yc6pITK
Mi3GkFHphLYot0JAARzzPN4asfNRkjw/YPq+BV1YV0gpV/KDiCp4KWvU55kPU+gT
6WkYAK6/7y8XGPd8Oi6qzgW+AdBY9HRQFLsIpZQ3ZLUfiLfTCbRUogqcotVfC973
qpDwDMd4bNbkTKwNbeMihpk6eIps0zk1dpGzfKnGac8bctCbmIwvKFZwzUXUA1fF
Wl2MAkzrYAJRrWGotkgtXf6NYz4hEwSWM5a1mTsU7YMTKFRnB9XXRrBR8gxBpHaH
9TuMsLDK9GkfgJIIXZKaSIabMHH/ZBvRgFFtXGKwoVx0lcfDuGpD//NlcwsR0RXR
5FUgjiYqCptfwb0iQoqagF8W0CnlgSMpUHP0VHAxzL9oqINB+XqQlba/+/V8WLxc
dh9weM3f1kdCx/wNlLWIRqQyP7fQixrY+aKaaMGTZTqUh00McoLRL2lg7CpIPvHo
XCd8rvWyTebbCAwwTH1b+mvs9uo0DLFX3Ten4sbCN4s+IVM4frfmtdc9IBM7urAI
WmWusgah6y1C2uVJ9oBKsS6BlF6B7k/r/u5lH+JYi+6CYNVrP9iD3RLDuZRXcWPu
KbTJDTXAHQqNOfLysrzIeFx+GRMcM9EDmzzAhkegJgd44ewKKOBzeOqx0ErogL9T
vrEm51N+/n8L+nrG6ox68kHP5E/8wPgswWJABDEV4d0b0ZGcbU7RoYxZXMlJ3muk
O2/URoN+Q9ofR6bfAl6sFnspZrXNWdJmP4bRUhknCGIoOSpWtvSAA4Ex52A7s3J0
qh7/WWGu6So2dYMl38RgFoytXNwAzCUcXS4hwvG1EtlbCWrOFueCHvpyNkG2c+Tr
YA8zPfgwaDyqRl9IZq6Q+HDXSUaAjy0XHJ6ng+R5ZeZWSvY+amY+QPH9excx9KU1
LbqoXczFaqw8Tmsd6LimCxwRF5GyCcGesVf99H7PY8hXvxlgX7E7VrMB7yM8397O
sYVS03Y+9FcTRjFSZl2hTSI7O84jYGXkYdslgB9fisTT1aJZnM8c9m/DaQBqPGUa
TaUOpv0YNvB7a/hgRUTYu2h+nwEULamRRAPMCFl1ijDWF+bdk6n7UXB0Dd+MZw0K
enpg+ezl5QxJ034nYxeIrO80LqmAnBazQxfToLm0yoWWVavYbs1O6OiexCv8R4GA
qj4K4qkMoWYUiHBrK9cm5iRQmtu3BZEBYCAm2anTIpVfVhuV4FL5P2Y7lcRlmxGA
1qY63Yc5f3eD12a1QU5lTByp27+oK5TZ2By0sfyMrQCsufm7w3oNijW52yy2UH0M
jsDMv2IKIC9inEfAmbw+t7YhGnrYC/IVl13WTeJ4GWv+KGbwfR0HiORWWQ26FckS
EVzlEROj2BnBpkVg7x16iIb6Qxy9XqGYrwbhgxCPDwXSyzO6vciKMtOafQ3kFBFE
8xBcVd+QAtSphBOZ3j74kMAk2T9CBu8UiGoRfGVxwgL9/zBLb+zS1uv/TMjDkFks
V+13DuJynVmgxzMhRACgQnBVtc3/rs2MG9Kva0A6th9jaNX3aqpbD7h8dB+koCjq
LSOEEVmzI7roj0TSoiaLSa+nNgtVkS1TMH8L1xMqN3chTOnL+dnoKZSdgWwrnzC8
JdlfvZZVN8fELHylJH9XQ/lVOXXgk6I53O3VOWmbKLOmS7gx+aZXcrby3FqqXFcu
7f/y9onA/U9ROumyDhvHCgVyPfOPVX+xK0PSNowAczM51Czrab41YcEYiKw8YpEO
a9LLveBD66vNjkSnDa5bKpFb4sBDOiC6IvfPaWH7tfR9/svdczocUOFc2Hi++Fjy
eTzBskS+O45JgI7WwX3n58CcyNQkBHk+vkB97on4Uw50SqGahKo/cx417WQ/Bl93
oGk3YYcHmeRyB54gYbWlfHL0BcGfuij+zbrB8AUrtxcYiXbgKuVhm9fwlbXcxxdV
G/WJSDl7X4VrhoPsYnYFhpzWYmYJELCdVnYhmHrW7hWt/wFHtDZoAlqvzYhSjcvG
/3jPTZjQyXeARE+m1aCQrDtK+30FuLCdjjiw6TrUhv64Bwj9isSj3vD5to/ZOajh
FymE0h+EGLHatPzbp+cemlnZOOZVcBF2RoonnH/MpJTy3cYAaZc88XtNFkhRzTQ9
pPpz+uMoRWNizjg1OuMG6swx2gmDV3nYrUjLXGmvU5p8ISNI1cs856YTQqytM2Hc
k2n0btkwHof8hWSJxIzgEizHN3w9YJsmZnUw+oaELoYQoKghHTRGWpXmm8vaqBKW
41/ThyfHzeAjhiVipY2lSxqOj3mdTSPlmVjVLgoInE26lmym9WgnZx1tAuXYggg+
QPC4FN6zv7phMAqeh7MHh9HjX964bS97E1+2SDs8QCKL5N8OEn9je6Bl6hMV0xvf
Zp8fSsoGMSu5pYlVxiDAHbogxTq0wuz6Y/9GMw0nxwXN425upwySYqO96YfJwSls
JxD11nav8TzPhh/VXdHUFUD57x+J1c38xg1tOeUeqGZU1f5Nqn/HShDWAUDfHGZ0
nwpPih0kNp0vnCLjN2CxSPm3YTwGrvfn9lTvNtHKiaHi3CtvwLrQ+GgWmbJTihjg
dNwE3Lasy1WPHT6qT8bqkvD2Zk+NfVu6XTygQ64xR7fN5ml4I0pRTeuPjkdJUF0R
jCvlPMwU3pRc+2jwDeYsrFiqX9nOaAsqqvayBdpSrotABJusLpXfURgSjd/YJLi7
ydMubSosD3soYqEaBNTx1UYMuIWCyoBXQO+KivVYUV6nn1ymlGMqNxXaAkAdFBxm
s9eApb9x8swenKivaCkpp+8chctoC7dleL1wUKFEx2EMe0JSfwNeLdwy1gZLrUqO
s2Es5tK67ttTSwk9sTuFv2lJR5CgJDsR5AcHUQG4TAWNIYmMVXx2A+1A7+s3l75H
J0+820MiciqwHTkzgF1eQSSRMltCJjsczktJwAz8MnpUPsKQSX3b1296PBmuqQvq
j5bbro2mF48/k9CCo87UH9XHiYMzshiuxFh6D6UZC+5sLxppvENeMPg+O1vWcnLp
Mx3ZlddWteaBy6lvBGmgLZq5oYekaXaTgh3+gnxvkfn5svW6CxXzSvXWG5J4mZL1
Qpts0qKO3zFtYRENUm8G5YHjCIKn9HFG7UYsIDpEcuAY9t1tWqD5he54JebASTzk
PvZin+jc8+9sMbeqiOi16jpqRzUsFwwgD2vEFVbTdu/U4ex3IMNTUrmmGILGbAXF
suSHTtE3DtNX9yJpHzElXsisJgNJGu0LZ/hJVIVd76szjQXIawJ9Y9Eojwcw5lov
sZqtd82o5m+fXyNEkIrdu5DbfSz8PioPvVMH2aYmzB1H0NiRVRgFQppOZjyIg5+U
991jCcHW47757ATbMn8znkT2qveR2gtbQtOZU/RK+L5tV6gThuiOZVllhzeXg3LF
5BIRZxFZcbArJ+w8MCKwZ6wPooIAcTBYridDqf/A2dZ7uTIl9XTQYSan9gn9CiR5
ZK5Kj55zFjp94wvIKo5FN8Wrb9QtgkcfHgrEec1dYOBAB/VB08drEnauyPF4fIBD
Lsds5gPOyXXp0ZF9W9StIUxUcPu91fWLtqo0pF5v0ZhfXdv/zTzJSi+JebbxBH2B
ToHV2G/NHDeBzVClHxwqZpe//3CEdZCePWbqJk2M9xodgkWpPVJKf5/mjuHWPaWD
jqZBAXjzkcTwH/ixdlnxTNzdYa9EI0FziIKAn5yzMchap4fhBJ7mCYn9mtKSKza/
G5Rhg2GYC1gDFu6oRN5IjMKKRsCxcCQFmlWZduONTuA7MdHotuoFMoW9fSunsRI7
WhnTh6E1U1WqrdlgFWYHlBQzgMYLE/QwhuCYfxULkCeEAhkYayqx0Rlx9lbas2X0
jgSBZBGcXK5/pK5WJhyTrvNzd7rJt/D7ef7z3NrcM0NEk/cElH3ZMvxXknXb/Moy
Wd/7v6gN8pF8ZqH8wdlqhKPCcS61H+v4rUvEkNc42spYNwUAe+e5QekoQjdbjKoV
zgUFapBMMEhJ8sackHKvEXpidWJIYBZrCoWZdzbt6MhmYbghcbRMPWa3lBP7S17B
Fy3fF1T9RFHpJqsObWhwMuF19PAC8UZCWwDlSf008pjNnPP8V9WO8cH4ZTMsTIIm
q14BCeQz5r4FHaDhymfFOhyfmtyFVrsdX9qMDrMlsxc485WbZo8LmvxgpeUq3Sie
pi3aQIXaobuSWMcUfwr1Qw8cUvAq855ur7LWWmI6HsxdrWKW62aUGJsF6xYmdTTa
4WHGro/Ol1uInBEhOV/Oc5fBCBfQA/4xTzyxDF22Zpjci8L6OgWuLgywZ0od0hnD
F18UqRT4kuvDK5vExYnfVDVmXfPkz+1WU8y00GCiFOybfrtLtgQQ5Ro0ih94pAei
VcCKjsUyV4VVcGpnvwS3rrr8SPj+QfFWHKzDHSbp9wi4fCOkcrsX3ak/ZvTnD8io
l/yaFLIvwF6yNHpN2H8CMvvWAV+4mOBeJ7lQ+9deNEnBWuZK2fc1JEf62iD2hybS
RuxaSdA3hy4NHJ8lLagsHYfxgdrSPjsht45tnStk8LLKd90TlE9RqZXrlwbJB4Fm
kMrmAyxhfu9wDwr5YmvaAKckEABW0k2n+Hos8UmDdpLrfOn0KlkuqKCu95iORzvT
Dd8oxOhSQiD70FLo8WPi+bXNExk8YmZczTt6dACGVpZ4T7uKooMnopTB+LHUXaQ/
4twYQb98KFuE0mIzxTKlZy+1v7ajs45wjYipfB51H59K+KQYyRgv0pu2SCDkZ4kL
VEUHhsUSo3AnFUnKy6uktjWAxPyxFEhRRq0nDhfcoju6TyzoLSjfsh3QCoHyo2fE
PWxSR96a102GMXyvHAk+7q0HEJXdMCFPNVnmmhr5qCuaG7p9yWOSjZOHtWEiuXH6
RbiBzS5FE46fj6VJOJUIPEpLkbaWPWzpNsNdwBiB27M79Jfr9ZRKZVulHM5RsF90
xcWygCQ3YIjc6wvOIcghvZbKS/LGdrDh6JWRBuWlIoD+J8Oj98QXXs4Xm1b81dEP
4s/KuVg83xkvj9Mu3R5RekARObxJYSg8jxVEZEYUIec0vsxRO2TRCT/mxBeuHTB1
OzZ7UajSMsV4uzmmwkuHZHGdjHiwFxznZ4J7FyD7xqA03leraRAp4AeoSCApgjw6
ZEQLFMWhOfzA42P+V5Txt8PUq745jJXg8oBC6G5x9hB17+JnGtkWG3ZJGIY3+cNI
jN65VMRmZHTfVzlV/qJnSeHgHEA5oLqVRsWseTrnxBr4A1yFSBnFQCdF4hi1C+9H
KAQOEcWnpeNbmx6go0yn/1fxGRGYsgFfkh4XE5wMOm3mdQyhbX8nlJ2sc+Ao1oum
MNiSBpXlHZFwYC9qZTwdX8JWOE/IDijlv1nHnZmROIXb5gpPTjK35Ef8EQN1iOjV
RlSZAlHpmjpwKQNguTpc/KE5EieWAjPBSMfT12DEI+9Kycr81zkYaNmK720TdDs3
G7Y5cO2QMBNjBU/bxJTheHak6rm4kstgtiOALwZVAUcodmeE15uQFFAVR6zPIL3q
LMAhWwA9HogpxWhr/2CmB2+czl/e526WJ1XDCuSQKJlgqlwZF2eiQenf7Ft+RRu1
3CGbfPoqNs24p4f7yITiLE3LSUDUGhIbsFQT+JUVFStYcSG6zgPO9fQAloUOX2mC
RlufVUy7lPOi/5fhkK9VI3bf1oEeofLumEWPq7gUXe0LyG0l5mu8BaXh5r0Keb+X
rzY4bmSUmlZ5wG9/PYhmmjkss885kbljQ4VHvUSudlEdorgFjiVJtn7qRCvtFhh4
fQ9w8uPCYjNg/NFLWOHUtdCS+1KCL5dJXBfA62QDJzWHastvfXSOHV3zZ5y8nWPl
bQFOKOp3PnxHXhduhkSKYAkhHhHPRwFxjPaFqvSrw5jC0D5i2r79SowRmIlg0DPn
j/KiSaygyWmDKDdkQs2HJWbVzgfdC5LGF85pbFbyZCPEWv+e6Suqbl4aBOcusDLd
l0PYBnsr/SnxwSRmlG5WuujaFLE29SEQY3AFWVWbvRC5udq04H16Wr7SxgnvBH3C
RC6jgQFse/lK+QvCcPktuKRcHhJoMGdlK4MtFIU9bN6RbSpbYgKPKkQ4AhRUx8SR
QkCIagOgEdaIijN80cei6H3KTKDe3g4ddbEGL3OYnzkz8sVjIw9wZ5l1OiE2jOIl
LDq7mKTAAOoA1xRyQ7Ri98MoHNolJnlZIRP1jKVrj3h/Nx0mgJi3druUtWod8HfU
EfKoXsIPW6Da9tRX16kacedmfqm7eoYwj/vQ1DYEV8otmqvc95hQyXzXz0pudGF8
5/X5Sn21lNLNS83hmWtF8yPn+9GwxlC/v4bUrTDsXBend1aVygW0u2AGXfkJ7cdU
IsVyKjuIJit7iFXtamtAuMd93FpqFlpXyhKRXBBuJSsVQG8FNLrYxKFFbouYYZay
N8xIsYoKRlm3kRP+7weuzoYhUE2OfZNXg0lbQoDKyMgos244xgxqiIzfUS7boZKv
LPdR7sZB8VsWoBjqjzLyI5TNUgCrAVdOVimNUJU5e5CZL3Sa6cuUWCeV6ZtB2qAn
A5q2BKMAhTNgxt/PUzXj5vED1kRuzX7ZJQiozN3cqg6dLZjm7NAYTnBh7vWNjD2g
fukjoWLb3ZLhNagdCtUqcPiqE+RuOpaExGDQZ/lzlpxGrR5KmJQflSvgctvCWJuN
N5Ho0M45CP2PTYi6THmD6xXOm9U4alEp3cjKAEzjRlwS6iH51IilBp3yMIwHl5rb
RPEza0cPWsmRwgQMpZsX1BxDYgQoZGXqeGn+WYxpky3KehOrMJL8jUTDmqLZu4VO
zNoc9yTwUa7ZsaqqeJ/+K/A/aqSdmpGXtVNvMajRra+GRxmbVEWbUYW4eRUgVeuj
RUEC7dmCia3lIlkXjypfRcupI1iM7XzQGEauQzVHD+YSFcaJApNnf2sGxmU6hG5b
rmx2sL4aToF2b9b+UMCHwsh79gOpRfVfFOB/IsA0FFR9Un7NI4OX3O6R+LrV77WD
goP7sg54YGnmHTl7UFRAOQ4M0S4j7dwPAsVskbg+9gnoPjWfdpaAT+JJavxxxtlP
fESDzWW4mNtob5tnmpdRdQEyT++0L/8MEeHQq/hlvdAoCjtU/5jhrIOU4i+i9SZj
zrUsJJmWms/eFog+3p5rRbtBIHX4v/swRUMGw3CaCUL+j1Nll5yEQrlC+acnb2W5
nwtD8MQ2spHmVcSxHNBaAXhUGwqVvNsWp3pUCX8bkLA972fCqUonNh91hJ5tHbem
SsY5u45qHzSvTZAh+s+tV63/0Svz9xDcmUDTW+pMPzUkY4OPK9nKLbx5emW3RZzr
TyxQNh0OKtevaoE9YAzMXAX/Wg+rLu/q4/YeH3DDq93wC3VlrOXNXWhmao/WUdu5
vRHCibB8LJiANLULRTr/jZiPDcNuvthPt0M4w66SVPpvPGhy32AnykekhRIVdZgj
fmIBNpdtrAqBW0VkK2GjIaRkiQxboevruf3KxwN0JAE9CefAIw10+hN4mzDcrnYI
plFStCzATVGwIsk6mrPDwcBtwZISeuPARiRXvCLXxW0oVp+Tpu9v0ZEEiH2VYble
0wGPjuVrMdr20duLKhWqlY3RQeznE/r846cTSg84eQ3lU4Q5hnsupSqAbVxbvFX6
Ms4I2qttRXU0CsgSD3kJz36rFk0p7/O+djuUsq1er/6HK81ZRxFX1awxp3Uionjz
XkCKwvfsVCT47BFCcgJ9pO1syVk8Em3mwl9OoGDbczOSdE7cm+o5ybItWwlwCD9M
inQE9W7knA9L8J+hBIC4I9jhLf8p6pLbruzjwuJt2bDUFNkTN9+jKqzX3KZQnenk
kB+ldpZb11PxnRe0Z6o3b3osGSxRN+KIMcZxLbmGv1q+EvQm/w1plpfr+IvuG6Ar
8jMIcwujovFG6qmVQ4lrDn+/cryLZYcnw4VcQaxTEByhUuY5M1YsWSePcqK8rntE
V0eURq//5PKzOkiK9ggxoRXf4aS0cdC660ShjzuY+2O9uPxwBTfH9g/+ETUs0FPt
4vCfNP5CbHvsAZFkEnOKj2ahOBBUDYWdE9kNQXkaZF7nlyuvwhQh+TphGiK5e9at
+e71+rve9QlPduodmDxgTrbElGAlZNrzIKecmRoykW6xQ4CBvTllZgJ5qGCijaX7
2Ai8riAfBqtnge4N+YQOdBvy+k+EF25kTzIGi2+aI8UN2NuUDiWGdwpowHwffCdz
cEOovO0gLElN1tPw26XjbggtiaGPs4MCNLorKXds4WmmiLSXZXpdNrOoMtlIoDSj
pYNQuuIDS0R/8i+a2c59OoIkCH9EEspjtxHMk803fzcPMLi1yymKn2ahVxFcAp0Z
bTTw0XaMp6ikk/4i+JXlyLZXP7hwzRn+dkCuYaomrrnsddmqkwn30T6/UvJfpqUn
1ReTGGZv24ZOAu2ehi4CInGwy0QDppIhyhUKk+HqXNKZbc6UyJlUpB5/PsxIg8FB
NWDbbA1Y+Wq3u6xHUDseuiSCu0T6uxCwhnXtNFC8wtI99uLtqV+X32UkXdWHGMJ/
k9tlfzoHdPRkuRPexCNNI+7HTn2bC3Y7ZUYX4ibe09NBOtVMwnHgN8QIbvilzSe2
gESSkLIuPe6nNt/DR10KzLKKG9z6qxiN+oOoZQ8wfDaS8+oj41iwcQSB5FSkv+kK
mof2Dq2no40P782RUuK6f2Kwr5j5NWMGOq6JdA1LY5BwHCw8+jKJgABDywGhl7ke
rfmnO7MYepKE2rp1WVIeippgHrJSatUut0MFwr+L9mep2/Lw83dKjjwiygxCNwyv
UItUILco8oHPEobYG0o2tK5k9RbIgsJh9AZzgYRVmWQv2+p++kXs1e5tZ2LFCf4p
1hHIcn8NPsedLI8tyVYtWjSa8DlGbXfTueRcXl3gZa9ir7uCLiO94VRPzTMFJdA/
rsSqSSLUYfGUwGvpDrK5D1p2TuymHY5qCeNZfxS+lJ+f4v/tC7twKFhLHH4oGSMS
pBgR7ICRwpJHQkZZ+/eti8RD43gK2nLVruirvBUsv6h1TxjOwb8vktLMWS6JAsBX
mKPSFo4svxQqTGsdGYApZBPHd9LP0KaCWlNFo1rPZ+IzfPYEeAyiZ7sJZQQJRyY+
nBU9Hz2UvPiE+RbTIfMkJmohHa2cE1iwOG9BgiXGVKYeeEcckSq/Rjt+fms23wVG
O4Q5td4xuCxLTTuPwr23/piDFwQrgcAnTbMzhfsOKYiouJDELw0wvTGrO6tvg5iL
swVNrvttBayIUh5FtedN6SPywJJ0N0cOkqn1dW3U+mc6gzM0x+AWOACCzlAfjIlx
MBjeaKNopTcvyvytP08krFHvuvixXuls0zvAXeEXJnuEbr5JXwMW1gPPC9v4wkm4
O/JaL4Drfr67MPKdItv6r6xETa243saUhGFXX4Urz6maBV+1IqtD8YKxQTRwt1yp
xNY5fuOERw2lWG5YmnC/KPv4tHOaEKBk77oVyXVChUva3NaKA8ogcl4tPswR0qgW
SWTdGCO5g0FZt6y/W1VgC4j1DSmfgCOp2mS1w2c7hYwi6epARNjp2nGqFOV4fKPh
SeVqL4ykrCtkUGOpPoYzf/jTu143T6ZE0Xk8tf0pS1HOJP4t8mrPZ9J6iysk7A9C
IhirwmUeLNZMMlmf7l6r/p9Bsnc+vXadOfIj0OIoJlp8u6SuEIVT+t2/c8Zr4pC0
Ls51lqA/O7whWT70MiIuyWGOxGkhkBOg367bGZJGK1Z60ZoElUndlsixZ+q83XmN
8PRDymU9t6zv2rqRoTbJenWquLfcHyZxHY2hDtWY1vkybdujiI5vQ6GuRqer+fk0
vcyVofLsBBQGXAc6AF10IhKfAG+q2F8HnbXf7eJdElmadX51gLIiRhyQysyjezLw
Ui3u+s8MELttcKpzuK+BjMAqcTnNyzTwXpPy2F4yaXC+Op7K3PA7aztlyxPxRsOH
6fIx+e1aeOjUFqA7mdfvqvfCKlqoMIXxusHoukHAS+VWBzuOo+Ww3s9mrFbox3Do
8pc+1MfOrk3WCpqj9rj28bHUyf0vkoTtF3Aci7Rhqz8BXjBXcKlJE9HPtd1ocjVC
jHQ+0jKWzkaJSRj2+zTkD2dm/qU8l1eqOcRhpRSKeKSvgVFP64YZesFlCfY8sO6F
HLPJVK/doXVXQIouUWlyK15Q5VPbiGsafuIT/rA0k9GMZKnW9cWNOPcXuhA1Xkx5
IhZuabF8O45bHE3l8WMPudkpaErsUlRIfqA4aVPZ9ZHQWFHqfqaI1ufRmaxHn8rE
JZaddL9zI5DRba/Wlgb9QhxDHEiLMuKUSfDwZ6Cr624JXnTKU5GVGeykumxQfIq4
W/2sheP8OWTlPE8WdlC/gnGNkl18DARq/9YDOYUlgjIDLoJ+yi89rYOYJvJSj7Go
x1m8LrK53CU3TqlsEb09sakqnseLh9OksJBMuGCac0JpEilpz70Ifa5Yv7Li2CFi
vh+Qrv3pffAspQh6rCXyAMwAMs0h/p0/sVSQksknmrN+jhSbjjT3Elz5pCcITmNN
oXfDCysAIquDzSgoVOZ2J02wnO/uusKasrs9w0BofiSyCJqzkhk2oi2BYmgtdWH+
txV+Fk1GucIJUqz8t4VLbi+oZlthHHkTVMhAYzpIXhuAetuB34degQCmw8oH+gsb
OUJPpop9Tr06lR59NtLpFxaTPjOAZ3sL67WwJW5pls68VbfR9MhZSd5xIj9PCumI
C+19nCCPLvmvgcPX4T4Z0lSwalRl2uRJXqa8W9vkO1AOrh/GZcl2mKd1QvmPS7ro
RE367R8Dq4gMe7ey2aH86MfcXZkcYnL0e+AxioZgTs8KBJxZKb3+Urf+rOtlNYKr
/DXDCzOYmBZddnO7ITCye8wu3yhgtp2eqMi5na2unZaIyPwEejQwvnH6gbJ+DXM9
CB5dq8IuHEsGvowBR/Urxu1iN4pp5bULaB95Xl2dShsYsSgOhwZ1/fzIDwgvU2LB
ILIZChN9VKgQ9b/e18EegFPgRwr5ajqknTapKBO7G2q+beko3D3qCl7d8w64PaL4
KJXIgZR0i93anaQ0dvq9CtUls608q7x11SnzW2DaVX+ivlSewQnc/ucEaUJSByUI
pHwJ1+NSqo+FuMIyTohA469MksJc53qnHOaLW6gx39PgY1tyHRQqSmoqOnlB+vKW
MpZdDMuHFNP7OwSK6la+lGl+SRLSfR1mtoNB/g/tJ1dSRgcOEat17shG3Td2OZBL
4Tx2nrLLCFI8GiYHY70W84ahEk2JZA2X8z6edBdsoNAU+ONt/JqR+3PGxMnibPye
vUe/gEGDv1Xau9+EMPivYkEWAUPKcNzkRWvpMdzbILNbIwp5KvH4aQoO9eGF0Ici
PTcnRWCndE8TqUhUVfFrGyQDorivO7CMRS+T+8ykZHKtYDIxt0lvOUK6HhO5Mvun
cUtik+9XaCoO1HAzWMZyC2jaZGxFPyWVdUkYDTp/4ZCdp4u1c5Hsq3wkewnB5PCt
LJaVf5tcBxOStCbYm/oYoK+r4ZMGNyHELgImGZMn5XZrqoLpF0tu2P0hnbKTRleq
Rcl+JJBT0A2JVqnkOsNU3/BVCpycS/vnWzK2Gw9chFGF24oxUQoIBEWKKhnW+RBA
7gId2X+25F+WQiGWbK4vYnqKr3HJzWN6qxOH/CeOYOJisefHOH0tgDag40SCEIgG
PTmvb8445K8qtpYXmWYQiuzcT533V08r1muVpX0P9JfC+WFe00EHXMsMWYT6T1yD
ru+VuuAc10zsqZUFuU/EG0lY1P48s5ppuy2Sa2atRPPgxKERDC/+A60swak4RCan
SQiaLvlNYQAvPq+7Ijzbl3U3zwkaTdgxcrizFydEfbzbt5PMjx1yt6Zo9YxOXxoY
Yky4ExbeB97Oj0rnhVscGb+Qol9YLJvTsBBwdhlcVgBZ06Yec8pW/Kmi9lctaQBp
smScN9cins5mOYyWsu9rWA+xBg1xrPVb1Ziu7GQdshVEk84zyibBfk2z/rozTQgW
50kWMux/5PjPuJ4xaJSNppn2fOGqCdicXBmJNOIXd7tuU2MhKsTGtLE4Ob5Xt0a/
eY++WOymiBXLTlxxWyUznfqV9fZrMfQvks3gkw1zJUJVyiIB8n7mDD6Yt1M4sba8
xb5qImMrXMTeB80aUfYGo9FykSk6OaiDqaZJYzeMuC5wKYJSoUZS2SbG1zgrB/rw
w6MrHlXEiWNLbHd77mxsO8apltSWUD9wuD1lDtiSAWRdk3980MbKdlN5IvU+Pvrv
r0mfDK24BOoP0kX5TO5MIbLPCSc1kHqX6g/BduXJLWjZDfkWCWV22lbim/OF2yRL
H4pELD1vLaVdkHvLi/yMgYnM4ymozmKwBhdevjErnImmuWOVP7LqZYf/ypAKjASw
LxkLHT3xNL7JUkWcEgru/xB9JuLqPMuoZIn7YMuX+0H+Szn26v7akU2ld30KFTIP
RGG4G+CNUel65FOUk1GGvm4Un9djZtNJX2Q4O/yPicgoUYIFhpzeX/CNzmaXuVPM
+ynFR9kThpYmB4ycUr3CSNOA4N6GfxJq8u2+0da5i/kZvoYxSjz6ppYUnEC48d8E
abccNBLcG411quPqxW/4f9hsUC8x6NMAxfXK++tnT6jouF5LhINZ2rXE7DWqIdau
pJzN3IqqQWZfHV7y9c+1TB14aHf4EMV9oQZYN8ZNdiVGn2gDNgE6MubKvYUDuSZf
F4Q38UqkjniQ0jEd7k3z8BsF1hQcRGCot3VC9H2J15m5ImHsZLRiwDlYaVtc8Z8M
gr4HTxgZj7prrMP1F9u+dLu2qcjNrXS9i1W581ioB2ja0RIzdxDdi0EdVh3K2Laq
tLEHTCdBJdw9iX/EMFZ/tCql2XwSGs9sqle/ZM5LCTsjGsi1yTkaVLNFAT/GiUil
VaZce2UsOwsaH87qfmck5Ygm7efuuIttXswa39yGPQWmTp+ybYDPMQvzejoREs7u
9Wa2jmpUDxwa8UlV13JXyg34iKn+rm8X+82PBYvaAs1QNykAGTMzpFwMmqUS89s4
HCDQLIS2mePp3Z0jMN47tbE8gwZRikWTH1r46au9PMBvfpdpqyfljzKehgnY2Sga
LjXGaygrCmVx/N1mQRXxi9Aq+DRtc+0kGsnq2J1+ryl05510Rw+EzwPuJWCakbDf
1HhzPZuph9IfAgU1ObzGLjADeSwLOCqr+Zj8nrbZrRISLdZ6wmp10vGwihedxRRx
+m7m9m6V9DOO0B+UM30nc6EVT8XQlbSHj1pdE2n0ZKcwJRr6P8EaeyVMJPV13Z9E
+Qgs4zwmtjFjYpTa1mrtRlRJL9q5TRHdKlgZfu5Bs/TiYvzJG2loC2+R3rbem4cG
g93o6X75vnYHmqYpAHxwxEDf/k9/gYWjR6wHB5vGGvuxAGKitCHfAIH+ioAFiSlJ
RaHSOlxg98EWHLTK0eOl6XSxkEbOeeF/UbYFTsvNl4YrR4bDmdtgwlal95BYBNzq
NQXFEOB4uHZhu4YBQsxJI0roVJpYzCALQVOwZ53uyaaZW6+SL238YGi+PP2O07/e
aUWUxqlF+xEH/CJ/cMJvB9wmEZ1480lFScEbvyM1wZCyH3nDZL9trqlJq7sdBPTc
p7yg5BbAsYIspv3tSIskCYuDDTHzyQ94YjbY9Ga2KZpHX8OTFxdIIFpU4N+tdpdR
6n7D777E252qzXqfzMwy/HQTMrUFX7h5FpEil/YhajLwV0nMi0H4tLBRu1F74qGv
eBF7otnjlaDu8YAWZc0CUDADM3ZcIUi2M8V4nQO5ZnlIrv20+J1CM0Shv26lMl5d
XbaJhulb1QRpiLEkZuudmUH+6PdEod8fWKUc+OTw1bh2u4MCoDdexc2T+gpexNez
OExyopqs4Iu4Pfa52gpppmn60sWenW/uOzsvAdWsyz4ptBgRC7zETxkGGCsx2LLM
tuOhnMREzXpQ7vceztp+BQl1ptQcwklOGgJ6LpNYtpr7WJXYOua1kkue5uWGiQck
cudAJaYP0Ux2EsrFJ/tdeEVcgM77fJBpI6t49nmgiP0cgn03a8lfcJ/gux6Fy7k/
mQNzMdn8pPOXIR2kbYPO/MC1EGjziMp9Tr2LMZCbv5hKkIzIY8TcZ6uq6q/gPyaH
YJw/ZzmdJRMA/7PNZJl5oI5iTKnuAxlqe1IYUB175IYeVWPWxIfe1DwluNJkdF3z
WC+tliZUkYhI7jDRNavoYECOU2ngNzev2oBnlB9OB4B8oIRgoP5EsrJiPRA/+gZh
tV6OPOMhrMYmSmj2AQjlW0txH3XjX29abNcDFssHYxgvPFBf+opm7PEmPzGstUrZ
ddHgHXShJ0RsG8IZx3o8xXw0Q/galVTEpnRmzuhqEKl8qQuCrSib7S37AcaJGrUS
DPtmD2U/0ZGnNPbaNxBykuR4bKiuOAkM/ONwQEOY5T99ejhitVGkV8e9JS0PvqdD
yNSg+S3qdEN+GVWapj52iJSu2vO8GRwt+0yu/p5tPaQ028oBrnx6OdrJMHdCSCrx
6V3JJBcNJDozrTpAYiBLQCuFsmLNWqAwbiJinzUq3Y+TjqrUvG+HDBT4hpJ/rLv1
yXAySD7Ny/n4LGbJfagcNbJoO0as5fti+bMSPtpYp+tvG3jpXG3LjlYx94foGdoj
7u0fHxs/ZymTFT70JSsoTuhrJj2KYc9vJVNxWuk9P9gSj5t5EsOVCAMfNQYdRgx6
V4sXQzpysQjNXdo0vPPaY6Lw1D1y4BuPQi+jq6C7TXys/IpHCq2khSSBd5lnr6Ma
pAkoTRTejPtiyi3OB5sa0IbYlaY8bef8WdCjTUM06N5SiedLR5ZirRomMZvfHxIG
3RvHPIef3IEJzC692Zwf0PWZ9vPYVqj2wPYY8FqQu9rIO7ULrKu+Fh5k9v9cUvWm
P2zSMuLmN7Onz/1afihuO0NxoCNzIG4dtPlKhEgnRVsljleqqs8CWxagzh/MUNEq
wTmKe+2NwJLYKZPiHcNpMz3v32S2gYSfwqmLhhSLW08/alCIsnLWSkfigY9hPed3
pkabG+8CtaRTQpp35ErJ8SgU5oM3m5s+7C1yPVqAJycl9UORcRU3mSV1ZVP/IIIg
rqKa3rgKvgiIgyIFBMthaKrFOeEV0tELNzOnMxEO9y9D0dTwORvwB/ek6NKJKrTr
wxudYTwleObvbqQc5cLvd74TGCG0WuiPgkJtPniha3sw0Hxs537scx1lNldQyr9q
OO7QyozH+6ddYn2fHz6xuIHwnSPXyBYixrXNyhnr1ElHvMeg+deMu2E2jBPK4yyP
i9kp49DhTum6aYHTcVycRAYLs62QY3Oj4qeGb5qLJNIyMwNYX21v+lwVYiSuIMgn
SdrOyn5eYJynP5x4MSkgsKOZhJ1OIebskct3jh8oQn9yiBdpyxpGtNXuldCGPjtq
o2ic9TrR/A4X8k+wXe7CwCKgvkfaLTj3nV6h8fM3s849NRQ2Y0yg6t3fisKx0kO0
mHB0n1Qy+x9rlKMg9OtP9aTqkEgH5z93bphcnswrXEx3Y378WtZOMJ4RZHF33WXo
Yyr+ycIByTbdwqTpLOMDtRMbK1yT30J3g4t3UWVVugUX4YFEsi8q52lN40gIiTYC
XhmKBL+S1AArhjNtfeh7Og66SPeDA1ViSX5jnvQAPQfmHHqGZ+RI+7uvdpNu9DWT
ts8to/LcN/Abo2Hx1h4aSq7zsleCy9bGFURxUKlDZRDhuZWt2p2NDDU5z1z5jzca
37mNLOV6Ro2CiGY92vNAnfZrUQEstzYSz3TyLpr9MwD/NFr/gAKOFWM6gJNzi/ei
x5YxItHP6iY959mm0kBkEi3u9ANUYTLR0HZy9dhTsQOgzTDclR078bZoH9ovFQHh
TYqhjwRA6wA9YSfNHI3X/lsaJmTo0vQiHr9ySV4w1fwmmJCveqsw/3ZcaqfrlJlP
J1cJWyK7PfmmmKfCrrAX8vvgzMYQFBGJuTv5HVOwde4oVJK8qKa0AZNf2VyyhI7e
cJxrwvcdKBdiuPSh1EZqXfJNcjnYQSlpTXh+BJjZMnWwFPOjVDq7m7PQ286dkcn4
1BC74OnYDnLHQ7d79K9xzOnZDagTGqVlQDkv8rABpo671i2NA2n25KfHeP5+DEvi
48WFmyK1qMD/8Z3zUkzGfActtSlu7CeQlfRkYJbMmVP9zWmEpAhUbx0g6lhKOImv
GPfL43UOYKq29uGPyjyTvKyhEF7+hqNEyoHITxsDiGd+tmBzU8wUKIBsAKE2sGyr
Yq9UUq/epvqjQw/O0AVDtMqE7ZDBqRWxwytim8PMiDsvfjBz0gnUAPlyWimdoXgO
6fjx4gSDorKmFEW8gEWLBie7kk3xq59KIiA3VEctp1bHIZSvqO5Y2PL3iSKwPJ+E
JI4ngkL/zFKygHm1i9+tQldfYPMbXniN6JTlWBLwSdD5LAP3rWWjotUZ26nBnJ7I
4N0rPOylBLYS2wJ0SMHBE3WYHscZ2IP+V+x9lP7jr5lrZ03+STa/cOJovau7L7Ke
K6IFnajo4kYYMm7TMcybMU58BhnHn5AaRl69sgnjzbpfCDWzw+/YP2baAAgdza/C
oUxpLCDdu7AM2czm7hYhnfhSHRSHJh8RcUcn/llkVUKRfbyogbFMBCyDroAd68EV
tP19yri2FhuEPKJ5w6g4DXDsZyssrxYOkeJhZEWQVlDSHdQJQwvVoDWDytXO8lh8
uYOy3DRVicfIp/ZD6geAwso35e93LTx64KMkHVtrmoEZ1Ed4FwRibiERE1hwyEn/
wgNaCHyKx3HppiUQFn6+P5BUyZOR0H28wh4kCeHxVAurP9XACkuZmPdXUhIk76vm
R0AMEPj0JvCRuzavaznQ5p2oaPub0pNScuSXo9YJ4BbX5gPullfRncZVleea94S/
r+FCdnCw7yG9GHFjYWNqLLcyj6pNqh7xJp6KezQlt59/1+8Y6DCFJlSwxCe2+4SJ
X2ZLNo4krrGZNZbK6eKzjMdISTYvy2s8ew1O9QvThmxgRyeAWzGk24o7UMSnc/aP
TxNvhluJ3kUy67/IhdurpKqfHab4eX3Ous1NFUfrkTBzh1KCTMx0mblb+L6uq6mD
YgDWz3dxki7n26NEXG93O/RybLP0uuWqC3fUxb1LcEIQopqEF9ZzAjnX7C3INsn+
VdzXR5izZD0KYywdDd30d+rfbAI/UJYWcgIE+D7feqof38w9XoA2sh2vf8rR+VVU
P2gdA4yy67S9HBt710BKi5H4MmCdMrMPJQJWfIOJzJmpl5VH3E7M31mTrOEAC5Ue
9MaT3L3pJ1N+3q+FZxbFr44unV1s6XkY86pBc7v+M5VRgrnPRkAz4KbLXi0tEkKp
u/gDI0jKRQCXvPl3v6t/f/BfBH5WJ0I4D0IA/sysbcOoU5Xq4jUEuf26FhBCKCUG
zMmcsddvVbDke1k+g7QryJpc5Ax7U45ypfg62ybQBiYL/VdP5scnHSRLEpY3Pv3K
1pAe7Nhgp+eNJ2DJcMN0jvM33zMBIOI8F/+LMgEt1HLjuZE41hNQQV+sPRYsE07A
MqUDYwd3jZcIl/T167by4NeiQ3AypmH5YqSqAU6Kf7IyPAQsVQMWaOHJLbbrk9C2
0bDd8vhWuCOEdgZk1qEgHTwZKStAu3VhSijL4TbbNyt5BTYzRqkxNVyDDrk3DzVB
hIQIKEWn7hcTcO8mAkYlpYTLNcvYyJw3BpcWt0TxBmgXhiw5zGY+G/vG+mRn2Ogp
Ck6yYH12cIUhSDODga0canLFXxHCau/NQfChZtMNBp9asY4PAmoVBYSBIFtoffjz
7FXNi3SMYw6pa1MQMjDxk0Y+JnQOTgb+nLA0qiBXdRfw04l0znyRsn/2Gl2+6Ic9
X2uurnlVnAA37j1Q1Xb2ueCjwg73EdsKUMK+kLwuyyqQD3ebe+KSspkYbxJ8gqhu
w6e5lUQ3fOEjtcQyeIvVgRBzCuSJbK9AyxlgvQPZuxTSwUecV7FBlhqskfiZDx1R
XMODEMgGLp8R5uQ3ZcfCVyeiup/hLvCUPFn3m3WPFqhpXpheKZd6T2tuoYhHLLWP
3HhuTSh1TY2jywczZl0dxwx/NTHvtOCDDsACSFSs7JEMQEphkP34My3XT4APYrDO
4NMqAXwsziNfzw/D6HIOdTFS3DX6+zFqSRvBk5Ccur2s/I3r3cHy6RuQwhNMEUGk
tYb02BnPsHnD3wt5Xz9x5/QiAC1Oc5gdJO4JMhlcD2gvSBl1y1Vv+uZUkVimVBsV
LLvrzwc4UtXwQwU5rjnSDe/kbFByP/hlIPEhtP7zJXr9ZQlQw2AQC7szNNIMXJwY
8vGrapEBW8I3d/BOz0gXHvESuteQyMIzlRu9lcmuKJqGEjSSyj8uvajaVoA3pV/Q
PaEPsjN9EDbiQtp5oYG71fu7wGvrL/qv/gCJH1xXCxm9yVSuCdiU4s0bv00OQ+Rz
17ck4INHY0uCMA4JY9/jVSRdjg5YiI9yY0kVzXOuH8hbZ5foegpqDxaxhd7qGRA6
l2vt9XdqkU9HKZHEaKOAPm4aGF7zlWwPQYDI4mjvjC79E79Lk7oaT3wTWG3j2Thr
46SP+MSv9qnjYxZgvjRQ4VGRx3c2CHFn2YqVtV2M42uQNp8xQ5bAgPZDQpIfJK3l
2GGxLqoXAunJD2W5Te7C8GMa9YsnnSOk1unEGZCg8L6eM+GMO0gKrQ4yplWMmi6e
fszOJLcvnkwVsYjVWcgGIZ9yZAXFgPrhz4RY6GL2q5BhbLwLg6lmhF317VjZWI2t
DfkzMoqhqoFPW8PW6z+QK9IjC4Nfk646Lzn6lDZRDIOXRsn1zTUNpe1Sz+yHbkXw
+kfxT5/PDaY4MT1y9rpQ4dGG/vgedj5IrhKiEmzjhbVDef4KalWNZODjae3Tp2V+
keRrTl34iEcZl8XEsB0R7MogiRG4XJb8vikQh+LL3OsDpTnZUqcI1Dv5aUtBCJQH
Bp+oPmJFlqaGJQk8M0GwbGB/7L2L7DVgnPgPXTnfR5pJf8VLjWwRtNBs01/7Czn3
2E7uMwx6mQUsLzgdbq4y2Z9MRG6Shb76n23m2MpBKatLc8qL9QLn7Wo6Tyy7+rrm
W76JiV9BhdUam94fK9+cuqEvf1lnTWnsnWS4kzYH0LZUli5Mou5kwAoCCeiL0aHp
zoKkNdRe+Q0Y6PlohXI+BP6vtUaWZmPOzWmF49ZsyHwA7yzW6F7lX68c90zBY2JB
KTIrxZAhgMTG3HPEKZpZswz6j1xpnAac1GPFLwqoH/DezVt7Bk4DlzDuLPYBRxlo
ZRJ/XSfH7hHsNXRpBbVekKRZD86kSz+D554FW4IAls4EG/4K5D4GZtVlD75OzzMw
OMAi31XvnG1Xpt4nFZM1ojMKarpuRzceJIlYiHyx5mR8AJqcCICaQUmfXzGaUxwo
OKkUhrDTxaU0U9wdaw2AFUtR5dDSGb+ebuxhETAPJStX2xgk08nSlh0kWQkrQgJb
EfyYkSnZ7yR/nYkzr1OMs3PYdWmYGDn8Op7tE/UkdYqHeB0lH7dg4iHxsyNGMosi
Vrw5qnpElZTZowpLewoY4CUEBhokI9gJaZd6X0czGg5GY5EqT6DBZC4ujfQmzPr2
/ectQWaYyUKLbtGh+wg6utBtjdNhg+vuahIPmHE9R468PynCYpRHKvNFV0kl8ntV
wZL1N9tVh6KJ0uMkR0YuQif6hbNoVduMxcG6QqDOQuVffA5GX7AxNkZ4V/65spV0
6hMOMZDPALH0M+Q62ubzOXtMjKf9ykRtyoqT/jZfnTTHPXKN8y2guhBmRwhkSQjZ
zvHuHom/hc6LIlDnVCnst/rLO/WZd8SphRX84WcLrjtRc8EjpdN24G4n6M5VlS+k
LbXV49vPbHL5VyZFVeoQ5dGAmEw7kF1/iFcr626bM4ljMfA0wY3BwTNp4xt8QLEc
FhZOXQ70SucgibvVv+lS9I5uI12Bhvmb6MYV0bbdFZklxDGWKz+Ozt+4g8ACqz4M
Cv4K/Oa8COuUae+/Qor28uDwxcJPiIAeIfnzmUyLOXbOIqVqG4bOzTdhF6tuLdVa
jasK+9Bh2EjYAXNC/q5OJrCUDXQjEF4eSd3c4JqE9fipd5z42pspws57f6DYNq9B
A65lrUTPVKzdxxy7izII8T3qTAu4YNNvh/ir7DdMRX9XTDlRlARMGxo3bX2wXahf
6cHM5WzNsw9GQd8gtsEeGSG+9vrNaDPlRgnx2zfW1qj213STS78j0uMi8/eMJiLg
KErvw+2DTxfViMJmwqcGwosmKEJSV2HByGFodajodRTHSVsczZKQvZ71TatRgtl2
HDBWch1WWfYAorcuWgtbCjJn4oD5LYDJ8UKzRirotPOvZk930nf/IQj7S4iRbi5f
0Bwq0Ahy5NDlWFxawpyfzYrkLm8/QvjT+ZOVWOy2bE7jaMZBtR6COomARYZwoXQC
74UkLp0sr43+Cxoj9QapL4fT4EFi7Xy7Z63etLEzpmrSo1JR6Ozdsk2+TVSoWHqF
s38MPqL8ZKKVVlEtrOfYAUzN7s8ptf1lbzFby0w7E1bFAU9y0GIQpL3akDMvevNy
6CM5xRr7XcD0qiXgY17Tu384s/4p5KaTvlOoBCtVZEHxiSCSClLkPYyKv8pTE58q
EJKgmjsyTQt1MezNGPAXDrgZ9FCMtJzH5Gp7GETyB+i5ocHYm2n+U97f6ARUurGz
tVrNAzbMN+HVWhAhJUIBHHuTibTlCOkoMfYitphtbC9QR5Z2NYiQ2zvuFs/lhx7H
mxaYsqLaJSCyZFH/z9mtvFgCq8Ey+//LpXkAA8t+2tqFSkHgzxHGtBS7+SnlxUq4
6WCbBQM/M64UXGs/1B3sTBFG2Z4YM6NSO3OYjQnXARSCHCOYeDCSvpiBvOWpqyJn
SyecD582u2qJYTLn/ALkj8tdkVgO4Gr75hW8k3Cd2tJhvb3A5jkzPjbKEoBROEhy
58yUZoctLSmiuvFKRe2CDy0gBc3sp0zW0cFVmTFR3R0/Kuad0dR7RXtUVc6e+W2m
nQIy52oBE5nljy4zMb87JNSQvxw0vmvDR0ntA7XIst77pOUgz7f+YQ/zevmOWYnr
2svogtbfnP3aH/u6SLHth3YBMuOOUc05IKJReuvNl5/PZSJPFPvbyEVMaDtMyItT
e0f1vNkhQXiqqFwNk3zu+2RjiIuid/vrs8LbIHthP4BrnENdV2XofqOMTRtaRlh6
xGXmz0SKJV3eVABow8BLz+NtmMfbxbWSIOiqhsTPTTtzRoF6inobkoKn/Z3gPKbJ
RDlcBqSUoh2PSStRqriZ8DBJkjOjVysXqWWNFVmsL/dJ9wV7K7yh/ulvrtuTgT30
jdh7X5Uwn1ZAoyUSd1k5MwGIAguwscIpl4lHZaOkPLaufV2j15OLWC88x2AZk9Zy
V5xecfF/qcRuKO2a8M+Cw5zVZVZmqu7dCR0Tltlhh9mPBvPeB+YMbOS25Md4LyDn
37XNzoO+9wz0vVWkjZkUXiC8pADInWmKYe6Lj9pkW52D/I/SD2uUO6AASjrAsJtf
RAw01bYX2rHoalt6PAv5DDQ9FrdFNipralZxVU+3LUKHYwn40UMSX3l4FjwE7Fcm
9eEXUwk8XT1okpLIsfLb0I+QqKGLb6pjmNnta363W1HtN27X+ybCNhFtDTYRRtx4
Uq6rZ9YoF3+EXNU0177TpMRLmF/yXSClmhFxIeJMXjMW5RCySprTU7a8kbXWGu/L
GBJdAkm31SHjLxdaKCuIMx8ttFi4v1/0iejlBDhzs2TdmJVyerL+t44xCUCpavrF
COGhcnl0cjP8na5C/lMURRxWSEsf1Tdd7KHJoaJYk2On824N/QAeCSqmgJOsNmIn
cLdOOgPoHJpxC7Ckixt7HuCfA/wF9OZy2TjmKQCFtddR2Ss9nvjJx35VcEXH67YN
a3QrpjJxCBjQDOR3O22BmwrSY6++GLpDxIdgrx+FR9W2CjD5Kz/9+mT1JXusYlBF
hM05fZ+HZZTCWjk+tKASwZqSz1hVRfOeT54qafIBn+XU/oPFw6fX7WEq3wS5VhRf
cqxNpdGV+kFu9B74YXweIDoTRf1uT6im2PRu4X0pm0UyKXHQtAe0HDaChIizluRR
4R3QJFkwlZg38zEiKGjGZE2wAqUHuBkkpZIKcc6iUqSzvzd3Xas1FhzmtPOjqHlN
cMb2ycuMm2+s767vjn3NFfYE6VENdCVOk/V1R+Bk69XM5P67rYZgKbY15zErAli3
fiP1K2X5SEZdmdqRs0AZ7S8F+FqHP/pRinnnpVNqZd3sf7/3VNIoGME/G8YW9Xfz
J9luTropCFAC7lW3gWOUS6oXr4q4C3QGGNDG0+kiEHtkSbsvdMdlJSK6BCkkbPjQ
Lm8saXn1POJKlkwywRgaoWqTsT2DcMreHAf4gmuPSzve0xDhZvmSRqW3y58y0SPW
LaElc7dTaIhyPPSdtjLYWJOcQ9jMBUy5bif9wPekugQ7UXMSSf/6YZYKsy43EIN1
pqr6rts/dwwFeaIvgOI6D0SoYnrlL/H4g8algMMmcQtWXGNgj88K1N80geXYfzFs
Xfo1Ar3YsjMb4IR3DigdKc7z7Xo6It4BFv+pbuSWk4KPzXKyypZKSlf9ngbS1r+R
fqTLggCtDn3SQTmZ7RS6MEjDeLmWXrvbpAiVELceRVmjk59bhuiIYFydwylPzf9r
2K15tMdeOoyCHZhVLLix3n+kNGn8U0lGKW66E0XRgCMegqg5PNhhWtmbZ3Z8s9eO
3VpQhGJEFLw42TuVd7o/YR+1sSy4MRP2EczuAzrfg+S8rXQxbHPTSEtU1qzU5XgF
/LjavNuAVE8SLW2XGUb7Y1vA+Xymy0y8qV/JnRJ4C7siNdWm3fyVLZFCrrFOl1uW
fDVZIrTohotdRiODjNU4KyOGiXZg1c/0xRjf8MfsaMbSTs4yprMMAuhuA4Olp9kD
N4mmI4RIBl49mEQ/yM98jrVAe+VTPyWugCHRPBaukUg26zG5o1AO70MHR+cKImHY
5zx6dk5PW/Pt/vbskzNp61gEyDnyF68nrf6b7L/cf9nWPQArvV3FeDtnA0CE64Eb
GwRIVVq9xhUnXDlyq42Slw0qLSPRpKOETbRIqvzW85M+cb7a9r1K2fGUYOngjHtT
/Isl3wiwVYDYhW408FrEoEp7EiTwza3DCxuyaC3Tj+ERAw6Pxw+85Nrs7zT/oTh/
u+mtaUghS/RRxP5DW/N0HLRasXJN/9ciWAhdUs+dQHgWbjRWMlsrJu4A0GJRl2K8
6CoaWXhRWsfvDhMUdV9qDgaLtb4A+lsUcjOTbEN1XQWTzqsvNFP7OlrYinacPr49
q9Ee7+aP2YBinypND0valnjzzrGG52plebv1sk34JXb+xd5mmCj9VWnuUM3j4qrN
gknn8ng9obcxHZEyAYKJv+6rutUZ3XkxHowfzY0EMNOWEs+iJdIo2cq7O8yzCu+m
RAdpx2Ckn0ZINfFliz9vpWpUHY+jABzRoPlXNm6PUwqxrXi2rKSr381zGi0vrBlI
cS2T2kdPm3RhTs7ghN1gLrrOGjOXdAW2clysClac8ew0z/4Vj0ua368YGDnBRVnp
klGYNLm/d3MQMY1q1YKv6k2mp7ClsT/TIOme8c31bj4NHn/8ygo3hkOYDVgovQgo
Pq/zXtXrnqgCkjcRboDZ4RDUWlS5v4/CgX+sA8oyLLJ/SjaRszHJLq4jHjE/dVYi
5OJVjmw1OY2bbHMd4fRdzglLZvI1IFHbxJAFGuQHtZA3mXSaK417xO/PMaPbSYu8
axENfgsnrC1UEARch43FQDQOuAigEFr1b3dTfoN+lR9h4L1KOCWxIcFV/yiUxiMK
iURlRougQ/3ZySdPIqGmlMYia3PFELa1+ZtGJwws15AOncto6Bssfe/F6oZfLqWi
jRKNo7JsZpdR0i3ORzkm9C8KocbA+9bWNzXy66P4mhJAYwuKQ68DmwCJBfR4W/Vl
nXfmNfgDQrkKW2+Knz5G2VGp/rYBjKq+XF9vkwpNSX938HBLBk6/VodniD1LdpFT
J8TFwzLulsOS3mI0ljNywh7t9Q6wgRgUaiPq9f02g4V7AEKGmL9lYkBvREPpgRrH
P3yY6b2YOU9a5iG79ZCGkhGLQyQ+lG+WxUNzrtu12bcCZUhK4iNGGcdlKurZ5sdj
PWoDM2G7RWLXfZkN35TELT/e9d+cG8YB5of9eI4Z1B3bY3N0gDsw2fDvTWklUS6W
0E7IMn3e09/PWzgK/c6Tv+f6eIpA/bC1zyj3+emHNP4eZiiO5OB8seS9Dl21kjOj
YpGv1c+tdip3p7oZDNmTKmuFV5VfgBdtbX2RW6MsDCftiCvYTMeuGW+wpTYlphlH
iNHPcQK2CjJ4Qz/BGtCAQDWv35TktbCuY4jV3cepjGIap5hlXYId4dsnoaHHm+TO
qSU9Lz3bBM4oXw1RGBTvE4qa+JATSDS12ZRjHBXOpR4d5CdWrZpYOJGbLpT+zaKI
89/iq5Oe2ilLFViSR3jTH998OyoYnPaZ3a1lJ+KJzNzx1/7agTMJZ85GSm3RhLvK
3LHw6+pNYSWEpI9vSOkkuhX4fvwnbiM8/YkYAcW8qOl8CiDfbzbY26BKmHAPxOXF
2QF2gcs9N/YWAY5jv9isNaEuXDCIobBtGkEUPEq8moSX3sMp0PQmdufRJEx187cY
YmFJnmXPkfn4p1HcT5iRraq553pTer5iwTNjDjwYECqcwr+Bl+cmN6oKrZZOanFZ
QRhzl2mwWLkPy6S5lBrqQ4B67RCCOyX4uGLPgevvjGs0yVDKK5urWIfWf93YYk8N
xYlPlkJkNrFyyIueNDujoEMnnLlP7xjXzbBm2bOVmXi6jcaF8arnx0/Qqyk5I8eA
boEbdoPLa3jqtJ6us+ku6Hy0is7g7+48iGLLdPAITolRTl3KxgPFXJQTAptIyNkx
Xf9jP76meZOOJJE7YZLckuvh6mRQZLwighm7PtnxhjEi4dfkuedtSuegleMd27a4
BlK/SrgaqrhAFsco1E1xh48CD0yflfOUfCDMxvzENoKV/cVK3+Ztr7WtBEaiSXMP
3ctjaMp0Mt5smm8Z0MXllWdxqvaFtQ3IWWdMqgn0NBdaVTpthMsNe02Yy+RbbMe2
fDvmt3vIdDfB6hVKQmqeRtNo71CC4GIi3t/5HGsWA+HVBOaE7D5xYe0/H3VCPC/q
crZgwRh26sAp7FWWyorAC+8ln+K/wsENlhPSfAUEewR0lnfI+g9kNj8lCyvtImLu
Zq7n/lO1iqwqzi8YWBUgIffdHJC8AAZxBBlfMygL5m2nbXb87Znt+tzVQ7W9rMpu
EwQVGdyu3vJJ3KE76DlhgKEXzKWuiUha1Utgre+elXdsHxr309RUBa27nW6S8Vm2
UjURqQTeVZB7SwNCzg5A+/XG3GW1Nf6NVSZdjbsb/4Wm6FMyMcpeno58ySNpKmJ6
W4mxCD6vxqH5c6zx2VX3+OxfT+pHDLOmc4h9uSVjHbufA5JAwUy92Ngs91LhURXx
z43s6WffaiN+FcZVHoSzn80MDnf4WcIWzf7T1cfKMQeOyIFjEnjTgbvYIIM5g/OC
jw5Lfdp0gs+HPOOWNcEuZuKXwJqMPeIBSW7FYw0TwocO1QCpaYn0Y8gUM+45cK+T
yVVcY/86xOSrI1iQP4AWngYOZ92k8ltdEaAFlkqCJGUyhwkrv9kZhiKlBU2OAuqk
Skc9ecdif8CEU6S+LmHYVpKCiIQN51mIqiz6bqBLy0vI/jPKW0Xg0vjK44l0sjRF
XvTpW1mZfR5mwtAE41+M8jdmVAqH7+B77krkGmI2CfvfDju4+Icb6fJqvoQX3Fe8
QPb4SSS7UQqsEiroVOxUIy161IRBGiB32iib28gdZY57JJABWEmJptTyb0zBRKiZ
nJQV3rZyb0ubcpsmKMzp8PpvIEp2evGeITEGGitCIxfO2hGrXPFXuMuZfada3G1Z
Hv1zrfPeNCCaznE1oF2JGoh1ZV4MCehUIKbmT6SZ1HMancFNGAHlVQo/W8cmi9x2
6xtUxHpKX4mRnMvsTell+lcqJXaqd8/jvLS/AHIczL/7t1o7nSqXG7z3rmd3UuRp
tLnYrPuUQvLULuUZGkbkRA1QZuEmlHd9lfvQW+q5NwJHMXoDwkEtHqb0Kkr9VVSe
iuh+LWbsKI15ltFq3H3H773aYcrSP0JC+6QN/t+RHtjiR0CNWGWHPHqUovKwbBdd
30HuFoZk3k/mBehZWOVX9K2rYJ7vhBijLtr0eUbuhHQ/KZTiS0IqA8JSR5e/YmRa
4ZHojmCeHiNJXwV/2DgfaN9WyZoCbZhvbv1p04OBx3GlcCZNeWYed67MP4E/RlEt
gUXu7HVXZEvBYkYfKVbyoVslkOQyz98JLaLAumgfVPLs6qFFHxJcjcXhCoW1l6Ot
oXKqAmtNQYcYy0yzdKfXROys9rC+eaAaYYHXufeoIgvjeR0KZuI28gjrHeHJ9lAx
XdbN2PCKj5OHJzISDScAyj1uYaVXn0aOYFZqg5XdmbYa8/4hMbORUwGsUct9jKsZ
VV/42FfbmPzQfj+MnU5bCOMogOBBb5A+50BbBc1tTaES8NqR/uOLwv0sPJBsL16j
MLPNufAbfkBpHENOWh3lAo9tx6ZOR0Yl+iWcEVplyHosZubwFHw3ic2FoRRgQ/G5
LUhqZQHVMEAcaaTOlFs1NLVndWDFnj8lf0wEesGFSsmna+66M1iQxpMzFCftZ3YF
U2NEARv5ySHvkpy7xevP8h/oJhgE9WNyHr2ymt7CFK7T88CHBG94p21qNJ1wZX02
gnm8xvj/ldsQvENVZBBx80oqXnpDq7upyIHPppNOnkAsYtDqeKZ13UJQY7tJKNXh
ALyitinr6LcDI1PHbif3lJSkGd/0Uat1gWyx64wvNyL1k4c+rXOw+/fHR8e7pL9l
Eq9+Tuia0xw2EIjWKtE1TKqnqW2dYwgNG6HDXEs+alzmcHdkORKGgi7KMl2s8D89
vpiesiH5sIZzEdF1eXiAzX6vIrV1a04RCArcPQcGt1JB/Lo0Fexryny3jMY59L2S
6SFvUugcR23HYklJipcVZNm5csbOCPlxcXV8Enqk1/PV0uU8U09w98GRZSKJ2qKp
dcoKFslSCZro601em6EkinIcle34hI3CKBrtkFUlfHQV0/A0e2imWVdeYogJTw+7
M6iyluC1S/mAMXKnTbhdGnggYsA9DGZKobPUH5uRbb7Ccuo2UZR82yG+pkR3zL5U
VkC22AenbA5w9xw1vN8DWqWqmQ+S84DJCoQumzF0kwDGQEyVTWN8btKvE94YLFQ9
PN3ru4etYRcJSTh0Hv9pPrMkX9NYsSSDxjG71iF6OuSxlr9vUabIq88uKp50GEQv
J4Mlino2i0cLR9t6pYS5zuNudFZCmYKxccc+o5+LJJpC6WNYOTPtMnCaaGM/IOif
k9To2G1Q01yOJGXrFxqPAuKt3YFI9HaxSggq1jpbUYETjtdaf5Gm+VenHlDx9Hvu
+kQu1CGtsL+IFnfeRr1KnQQUhn/lInTXYzOKYENgw7QS3ceRWfnitADjwsuJ9paC
SPIASidGbmOhrkGRhXJgD7YkJVQoBLKOh2VfZwJZrc7Bg2/9eb3PYcqShteOI7NB
2QAx4sHM4sOPrQH7YVtnUfZ8Zu3Z2rD5vzf5K2uuseNywsgc+fhoMfZIM63YEix1
UI9EfIoRi+6VgUzaX78ONLaaEf1mpodByyYYkAShfMP28rvqVWKyIwYmPaMTshIG
K1AoBsIYOFgUN348btqK81Co7KJ7McNvVHL2hdt1dVf2VAaWvQzmot1LeTwLokMZ
RDnNd4yM4CPjf5iTfh8ybFPhHUoZi6NJJQ6EvGKfgkqDkut9iYGjVa9uA5KbR0Yy
rxwh0Ltt6qw9jnjL7+dMnqhbCWO7GFXK2KiUYd40EXBqlPG+mRmgaayGeHrfzLpP
NHeUC8wRWxNk80OdybPKQAJHtqgwuBABpw/4IivdXwng08Qqasz3e5D5h7pbYjnv
d7dPRmYwaH4q+3RX6DGZrfkVXelIWotb3KFTLPLch/fHO4MSzZF3Fbv5sNmGxCyT
NtzH+aIAg0/ukj48JZ3gQ/7d8fULeD6GTt+C01dNIeSGC29WgCVIpRfY0lg4VE5E
zPfJlaF+6YYWoc2nHugiPAcQJnNW0bGzUCbmDQCNlRtuhu9jXu9c080DFBhoj42t
PGEM6p80CBunZ5CkneDs9yI8V9g8unQKUHafO+x0XqOIfFiNdP9Rk43k/PD4iXSZ
yQzAJbRkNG81Z1EoDyxbUimimkFGHIZ90TB1aCgfxso3KIFoOChK0JVAVijK9Utm
dDfyMU3ssW6cYwR9pNGZijhaSrRPVQu1XAQaDbJfVhQIj6EMUeiKKqJNdEADtC/B
WUX8MH+Qp9t9XVZ+Vkb0QA/vhIwj3F6TjzNAYhcC+wsrFDYhbfx6m8wpchR0kd1A
yACfCi/pxpj8KCXTaRDDr6Rg+FFHytURQGLOcYCPZFENsr/DxhXHFIFvblC6rmRK
0fgOkO7hAyTGuPOeqE7RKf/V686Gb2GyXyn7uQk5ShTu+fAEJBicHAeV+wSGdiSq
5SjFElp/B+aBJ1GOnbDp0JHeA7P71dUTpjzrrodFYic+Y2QL9GpmxjKGoAW0Z5Cc
Vr6ik6J8aAnKRgjnNdrLCLUJi7RvMwzUVtuVfTDih3XhYpKIR2SP4U7vXs4Up4Q0
mF3FppaI8V0gQ2Zzl//WMNldNLLyXI46CyeNyfsCM7LtsztmsNvc5Pf84wnnRSsT
HBaJ47RJfjyTs41Tw6/yQSo/f+GAAQ48lLkc9LTfIhquqpOnN/hcXIxTAEVe6bdy
x56HLRDl1PfqyXsH1naakk3BP0za4GsfxAE/sP+c6bW29jEqa1qrK4MiDI27U/0Z
zIGxGhgi5XcyO1uPkTBTaMtHVTpKsSCecjxMC4VXliY96yDqasJndqf/S66Bdg3E
5pwPSTYIgIVwpW9oHaM4TagRGuhFqeVkAF6YS5P721SQa31Q8Vw3JlSMifs60eLw
x6hjfEFXigsL/ra8bRr92VfqCTKhIvqStCXQ1fVVDmAP3vZ6ynNfyjlp39UTr4c3
SvOOyx+KP5UEBDVDwaU1q3WgjzqVWShvZxqEOHvtySW5aty9LbmKDFfwt+rD3M/t
tJ59u56YM2xSP/+rlHbNh1m8TQvSoux9kCmO/I0nCuY/1wGmvGoYkZ5/obvheuRc
U277o8wV7srzj10R4qvs28vl1iVr1ZXczpt5AQ9j+zY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkeQQsjs02+HModN+3bYj8fFhx8GethCStRSPt39bP2uuEoFjzMLdDIKF8d9Rlhq
+idZ58hSMwg+wnz/e+ZLejJppgXwsC2MN6IuzXb5KF1zSTIIxhdJkIBb/zxV8EcV
DQzF9nCeJ9Hzhgak6AlY8nVyaMfWlh/Yy9ZBH2NrI2nZH22CD+7IqA/5VcUNiheS
aPTNul8is8dyot7vpXgBm5OXac2UPmt+D9WTsI2OWl1Dp+53JkPbCmMUbtE5qVCD
3BsEm/ToBHLY45DIIplKAJad7IlL3UiWVE7L9Snt6/TM33prKMEMlgEWK7K7bDiK
fPgNYcICw6DWlJlXosktiDdLtnqU6gNrggSYayPJ8okcIeIY4tz0d3ErPIUbOm+N
PDEe6LKiskoFlUCRtZwnxT/Zf5sno7WiwDwCEjB9tNp5+M4ftqz7o5V6pjWHscOb
+vCJS1eovsqRra3ukA+9hF+l19sp0BSWSYgIuBFmB1GGMTrh1hMNyDfsqtAOkSSr
Sh7Sa07WgSO/WvmRxRG5TgwjkQTW2yod7IAOWkG+SjXeoLwk4+RJ8tME7cAeywHc
bLzupTuqeJkRzTirz4tbnZuawIt67LM0pI1Ei+Kexy+Gd4OQipnmJMZfi+4/OudK
SJSwekj06G0IyNsKa8f5Og==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QS/iNa2ebnW52qMhFETdxmFkgZMTNR40Q6vNsuprkqIhgdWVcdlDBCrNYAKcrsA
2T9eCH0Kkf0C1OglFntBbIJGPebGLy8O0LRkoGnYJf7/rtAm0kd5U5sLaxxLdYn1
QaPMwcRWiqVSmzDa5DEpPPo5hWYt6vg+FWCRT2v7TDcQXrQhvjQBWSiPysvzWMfc
iudOqLCsGA6tMSJQQdOwvcRxcz0iccmbgBValap9g37qkaQa3cKMd4QAPBukI17W
9t+txy96TU3WXuWJ03hHwoI085HBJVDHcna4ue0CshEdUQKk9atwL6/0mUCRxXLR
xf3kzEIR9F8eDslAQ8zca/cqdShK9CMS4RPTi8AFgUQrFIhfCUXW0zwvTyn+U1Pd
+6DktSki5cdzX2FbIbEzlLgtBLiePSETT+1rShObp3Q41XpfCNTKPYT2K9RtKfaP
ZXsE2hbm6rKdra/DxPJTIoNUjqjrsNMDNlqrmP9y5c8IA9myu7+sECVZT18iY09y
qorBaTF9/jLug3hs6gutD5LSBzod7LfiD8S4Tk/h9YZTSG4MUABixg7O8hM+zTc0
XAPF4KtaB0pXkk6/80/YE3PdEDtUZxtsTOWw63SVyUIFjvJOJuyIP1Svj1lCRCPC
tFMnl/KCBcR/XSgvunRird03tE/FHdRlaPr1Pgw2fExBwLcNOiUhZK2hYxTqzKTx
h1F+cshosLYsBUjybQolFTNXamK2Arkbi0paaSN1D/UR8dHBlJ+kAhTmysV+KAyg
FSq+9a2K830QiuQSoCv2aw==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNNU2fHa8SDahOutCaNrkVLg4Nm0EuDoisl+5dK52QHLDmxwyiuR9YZIrdgEqY/y
El4GhI7G3+iuU1hrHAjg/NGFtPXWPbQCHbO5fyRdDWQIvWby8QpNa87I2dYFkND6
ihxJoL5y9px1QofqmSvvejzNq2+90sw4f7JuO9oVH+3C2n6eMclnXImY651VXTO9
zQhRHM8jJfmG+OOsGHFM2hTq75t6xf2horqWk1KMaSGwqK1Svp2kxJlW2nA2qMmU
T1/sbIp/E0omkAnc06r0o5QprgPjWfx6AEBOR/1EYOi9EDu6H2a6OgUh3iizU7Im
T5Ya44dUt/+gZcka1EKRk85qSvlvJt6hkTLMiXowDWFb2jkz9l+ityiYa5YOGrXy
+IKu6nzLiFcg2gls9nzyCgwD0G1eWwMZYf+bPBxYD9moWE30wLrCslUhbDE1g1x+
chQm9dlzEqxlZlyzW893hwR5q6dHjzLXwbEwAxj05/ZCEEDNgD7dqcMGWQUrnbuq
MYgBXXvVKxB/tjHaPnWFfT6rOf3w6kBRAYrvSR823gjuhLxSQQGcRjmeWYRgEX9F
lm/dZiDZtNcu7P0YgtsePNli/5UztXlNE36d5bBG/vI1sCK37aeQBhqcZIWZvl5S
t3ALAgMf86JMSNDjX4L1G9giJLkbKhkU9YtLI/b9ZXklw1M9VTnid0ABUX6SxQby
Tw93h/4iyBuG1+vE3Im4f5r1SweTgyKmqSen/wpBI3Jxg1eITOltH0IT/IPMCY8F
Z7SXkljPyIVZDXEk8sEWIDjPyU6l8P9X0Wa1x9ExH5q0aWPV8bFiLeVlAPgj7D7p
2b2e5Cf2OB5nmO7iAYHljw==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GNt0RN8CV2E0Xz2iaTxRFO8wxQJf/X0YOj0zJDFfkIPr2Ggwmo6YILAYIQ6kDEt
qV9mjVoQ6iQKdfIMsQjq472eF92Eate+Z5VYiii7mAq1HbH6MSewL68/0LzRe0zj
njXigcxSaFF/ysVSYH2xOdB98UCvIL2QaiZ6w4B9yvkoDspctduYCfc++CKOsuvn
LcaJDlHv7/6wnzvfMM2+fhG+1JQ5KmUrjXJP/SEda/cpddh+winTTddFjMVWXeUM
yhqWWv3e20pRtAK0qNs+OA6GWtILXXNbLm3xvX61PgS4UknrJoP+6B/VOzjBLH8T
fGxHneTG8IttkxTR9+EtU0H2GFg7HlbbJzzTMWd95IJsMpqZtvF29/QNP6bwfF7T
0NFb7skcI3acTfbG0Z1YamhCKfyLkqjmEEWB3E8DlhnYRYNWyl+t8p6+5pH0zBs0
C+Fv7+Al0CMlw97jdeZAEPW9I/tFbapBV3/n8Mew3meNmfrkUWtBmfLoCVtP+LBc
ZQGAaX//ALrJ0wMU49fA1xvOHINNh1YtRKyfijX+jxw8ZGIABrfXxOBj7XnASGyc
HXKfkyrCm25xEzvXyZdOe5StckFxwsRiEjx0Bwn7xHE1qKoFA/JIUh9RzSOHIn7M
fVBio/X1brvyhbwqFWHMDSbdadHROj04rh3MnK+zfNvaDQ65Gn3K/7uRavE8E3vg
1KVatErPXnUq7qW3Kwe1iqfQUtqqe6wKzRucXFDcczNZBvNxdqkpOdN5rs1WTP2i
H/CNEmtI6WrOQtR6HZc0zXnhodjifh80chGcXqLpXuY1bTjpQjtMNO/RLqkG587l
mq41uXgLqBhcp8xwfTXQVfV2pRdGUnmXPNK7OKklP6k6bMkPw9bXau1EOO+RCro/
wmu3PqacveEEZbrJOiTRa0EPckMF6Egy9+Uiw2LpLOd9zTHMto2bWF4ZS1WYykbN
9ulROjQTIhV2OyyQCXxb7fn+vwZUMzen6/M7mIjr3oCubP3u7xRPKcG6v4JECuT9
bIn7GiwOxDoG5bvH9yCGMijs6mkvhe4B9shS5ExZJ+P/0dhA+MCspyAVkJM8bVjE
Lpe24E79FE3XIeSrN8vbVTGsH7S0dRGQipdOhLc7L4yvtqa7ZVM3QnSp0wSQgUAb
4NQE6QcNLr6MiX/Cph2EoIils6ka3N6wrxpmkgKYhyGDoaQsihAuL8ywUVmU8bgl
+dsYnDnJvcG+IVb4nXc1n/1AGIe38fH9ELXLYMAcK9ZGmKkXcD99i6PkDpG6sNak
yh3g+fA+Ni29k6ZdSDg2smugGOjkN+wBa/HpnFVi7VqyYhMInG5Glo99BGWopuWQ
Ynmm/DdM8uVQUrkMg1PVU34SJ2LfkRYvb4RigyIhJPgXKkBOitcW/rWss1r8ytKS
kwbWAmnglSltHZJaY57SPzjWs8AwVx2yKsqp7cafa0id0KUYbGmbuYeft/OLReYN
0zpiLWpAxPtUck4F2J0HVOQKIgaLlL8DR3BK+ZksQ2wI9PbyO1eFJyw6ktcNLczm
9Hs8CGfQsjALEtjgEmRlGsNjxLToT4LOFCv7m4VVkiI6kQL/ZwyjYtluEe0OKtRY
4c20J/ez6+0SZpt74+Jyr8bIVEt2H++FeBbHsnohJkGaBis1j0n2NvJfwaYPchx0
hNqFNonMhtcjdU7XWn0H4KqV1615BE8uhaC/2qmKwCdotLebxhvyXSjZ0plEmpRP
S7lWmTzngDMg5lb2xoYJ/U6XV/j7Sp10Ddd4OltndcORBzRaQrVebk0w23Lvr5tF
5uaa1DlSTzNdd0O4CuOg9B8a4s1pYZs8SxNX8dd1xRFrZMOk0EGgqwIihhqLit1/
8+G7c2Ii2ZzVZntt0Hn+pNMQ/kzuhdk837RuhZnA0vLMHcz/Xx5g95RFC6kRthtY
nm+vfEcUwLBjyun4KZPVrqXpRmTheT8Bm6bwIzV2wBmUAQnPRhDkJJXNhZ8Q00Gb
sVMf9GhK93JpMmVshK/jtebCBxT89/tTEvZbiifmOpN+ZN0tjFSXmwzsxtKU2fUU
vKKkI6dA34KSUgW+Kdkyk5znT3998IPXvzG9P+bvjbrkwpWBBXdFaUPofrbhUzFz
7N7HFplJPqF287uz6GOtev6cTNW9LjvYx16MaywKnyJdZVujpwnNwzQjpxi3Ci7e
MD+an5spJh7GA4gNUAyh1KnZr+R1O9AewlHalyhznhf51xzASM6UaANAFmXIVzlb
E7Ws/vWtEYUQMrq6ZAdbBA8UUPJ/VbUODGaC7Z1MNwUBjONPFLsWqkPPlP/CU3Mg
UnmCuvTU9cwP5YsQ4SHTJh4yRfgoNGIafmBf4Qj3mVWbrF40PBd/oYk1dYVB4n8a
XfxkAEBbTMLANncIat6tVxUs43B4OtKbkIQZmLNc6Na5FCr8PFpRK5XBIZRHhspJ
4/TjDr8TWuNgunCAhF0NToOfqS+KHCwQ+E+bCJ4rAxihkgKefeK0vqHTFhvUHJmH
dTDMowaUoq8Q5eW2Q10tJ09TxsTE6D1TjeN8x9Ruvy3/GUawLABhn1kGtihSFfTi
A3vE9V705lFl7ImrsMsiNW7SI0txP8YvGmEK25zJKyMdkSfKj4ivuhxI1B101NXs
OYWp/uQuvdwWoFZ+Z8it/n58KIFkR78RY6X23e4op7jvulB65NmQJn1FAnJN7I1w
IJcuK9qfcBxc5HFIEbad0K45vg2udlZFOHayWhGEYmPv3bcHVGoFRMyXU8J82WTz
xp+5YfFHNN5orsZ9TMmn4xbjuTqRZhpu8g88FOw/d65qIV2Dan9NUFsXxHr+IeR+
Ourtq0E4j0igo9yeW31YJnqleuhI5S/pL+Cf1+ip0PO2IjGyn+etaCAp3BZDFIHM
STUHNe7L2PXXPIOO+2eMA7gj+EGHzvBb6jZ1jIRYd46ouklbh8SfToHKvtEDQJ+0
bN9y72WN3bD2WawE3ntsTHOqub20fO5qiSRYl+80wJDd4f9CBT1O3s44BCjx0cAE
yRjIDcBh0ibnDVfEwonVl1jEPp+rzTYud9mTUkIyPQqJhFKb9CWK+iQGUQyWpLKv
7xdygryFNewes3QT9hV336NEzwF4v2GzINq6bPOMtEtV0ozbmB0WMs2mcMCg+cdL
ifL2yadPt+MY0VFgmb90lLr9h9jxIy34SMkFyURXwopqmVXUPC0FLzKa19WNDavV
07ljpYfSXPkgQ1ViX98ewttJXsGGo8wfmrwkHKewb+apUc0WhR96RsmimImghQNg
EddlmIPuNIDq7TdTJ8m2bvEKm8MXIhxlvobYjerOmgsyZQZkAWPl8kvCoL8NwB7s
//jruQQwCwMNKLcENTWZan+uisleXKPdtRUzWQWkWf3suMqCGZAPnQPUry+PejGq
vWRffWcFdd4WNLhMq0prU64WlidYl+H+3jo/k5u8dOJcXcbXzAI1t64n2N1BiReA
DnVuvYIfml84RFFSnesRFfsTY/cATtRBSYZwtZKKoJBpuipTIG5OMjD0dxwAHhXn
BHmDaiEKZwUcgvCwuZZ44FpIXGywdpnJLGavdu96mDYrXWnlLKWhHiBCs58tid12
1eQKRWrafozL4dIITuSZhSIQqz6o9M6V3Plg3R4xklbr8y2Iu8gNFVeHs4XKM2T7
aDQIdNCBIBxYfHlrDssOZ4//iKRfBcMm6+Khs10QP1Nc+kOarlNG5zxVZv/e4/Qm
95Tk24QnYcRQol6cr3JGjfF/Gpcl0xCsOOqfblQ3RNXPmfx1DGYeEdDM9Jv7wdqf
mnCpTLLwaSM+JxGIBUhm+anm8AbA3WfiQ+2euS6TTfUK8pHxgomPuO4+Tj2/hIJ7
PhXu0GBXzz5Puz3KQwUWAaPfCpp4iYQ9azJyDo51mRSGbIq4tfgsYYQSihs8rx29
bO1MfPrQ3TK9X14RUz4myrty8BIhC1loFGF2JFa+SUGcWErnivfRZHPlX/UUVoDk
BQgLqyYAaPB11Tl4JO4bhl8YOdGQq1x2/HipBTFYaW0DG9fdpwRTHWIWlevnYtvT
zbwSg4s603vGBQluEt+tmGP8YvgdRBFCdqszzBK0O9fTR+lyyQlugw5vj8eBke0z
3xMfpK7CxvGri+qnjJ0iyqhAl/jnzdBylK1ypeGTRhWa+mo74y3zCKvD2Qx628we
ZTp0RjWgFcoh5RswCxmLxIiXvfb/9b/zhwKGuMbNvC9Mh8UoszmmjW333G83wpjZ
0MxaP9yt0Vt75W1Tpr2pcyjRAVpBPIfSQf611Z0S6APD3k2geLOT8KN2K84n6YnY
n6DvN0JZjMKG4/oBeTfipGhCQibNjquP+fS2NDXEoO5Mj9PnChVlb8Hw35qgIdBt
3poTtZkIFPd8bgLenk1GO4Olz605fwxxfkeljhFIMDgJhMyTmKAnRo4Gl1nA5Tcp
Duf9x4bmhmzlJKCiXpDu07owIxsxd8aIxNZxnHBpECnxyJjnCdCkD6d6zjFtMUC/
tWVA5SFqL51ebQPQU3pOoNEvV//jkn9BQ7AYgdw7HZx2j4EioedVI6GiSdkkSQH3
fGZFXtvtGUBsrt/lxKDIIkNLzl2nx46GobPZRscYheKoxqmf2mIxbUZhYM6Tfu2B
TStZZt/h8SfYfFbhtnieREcMU0dXe1dguBTYgyyijQTGASSPza1Y55qKW3VnnAyf
pQx7lSDx7N1G2ij8SPEbxwAbLR+fLLRABK/YNVREnSmVUBkBvrMao7oTglqbR2k7
jv6ZHbqV4hFQMvFG442EdvhXmpRidtGS0/8efO+EGbpFFIMTatQh0oiLjlvsS39y
fS4QYmc662rnETQ3oHw05H+p7ZeKZw/LqMVSNafz4rd61anfINbgDlF87Bzqx2zi
YQBBWgLNiyNLJ8KD6oYTgOIvrYlmCsUHXUjDOFrD9Nb4IXQYM7ICsT+rR1+2tjXJ
NnEJsep8okcIEuG6XymFN0MXbmru3v/sMJUQhYD8p/TaoTgs+UlFvs8BrkVTM00t
425Euu7u4JwfGbr+Q4jD4UFicCZc1cRJTM9v3bC/ZMbeGXEbfjyBDTSIk4LKQqkD
5n8fM7ce2bhuU58bC52HWDR6P7VZEgo+rtJuArHCJasQFgNQKGtRRdwIOpC6uhbN
o+Lz9HBLQjZbMQUiu38wpGhiklpdMWR01IftsWBry0P4GHmjI9bfN8jF5JvXG6lw
JAghRCe1bMTYHG86FfIKCy+kqAdKiglmDbHYBDY7/fZF3Lrdb3CvUVgh4CwgM84/
cj6CSDBzsXGtcufYcH9vICoo1skQsm3EtE9OFtwfHfQ2i5WsNhltXrr9jKWP6JoX
yZRn1PxFqbSQD/TY9tTMwlzeynF6vaqT3N3OHhf9J/KbY7mXwc5xe3eNUE2+lNlK
PEOi6DQ/sdwZ/mofKq40saIzqzj/Dsx8rEPZt/08i6iJMyTLetrtcFm77xAX63Oo
YnIhcFzNNfs/gHtxSm/DFHd9o66mVGnMoDZLdUm87J0visKIq3huewM76eZeTa0x
/vK6vw2ZtAml/K1VMirLryyfSMS3ERF2EDjM5t1GJgoGf2BQyxAtKn+gZJa9puZZ
pzWhvw6Aj1b+dTNodXxAcL8ycfBWkWB2SxvWTcfHVeCfFNNf9uxi2OaEbruulPvL
3ahk2HWT7Y5oOYK9dtTqcBIJXaegFDzeC9HG0QmUR1MVjobWdKXWFfFHJlRn3XFj
MfJkpuchK++/qbHoyfBiQ46mmI+OCMYzSJmMCEpDYUqd4mQhqIYYOItZ5S2Gxfkw
11Gl3QmotsreiZDv+8IPQ7jA1dIOT4FX+V1nvfRJpqL7tw+g1lA663KeRHQcb6u7
31whqjY8nCGJ7cTXNwhiFA7cXxO5nT396AMAKcmW3KyduC/r840u1GXyAMPOMz3m
fNNebVtK0lxivMYLW/6P9xyrqWld0RoSvxTs9EfWrsFI1Mmh2DAd/tTkWgoSdrlh
0zH1IKJGzBxFT4a/0OS4dCr4No88Ywev/MPx2ZxhQNnnwoZJ423eqK5NgQ7rp1vI
iCzYoFTqtXEKfmyfoB1kQZu6CG0Q+sLpMrBCxOxSJHePiNx49Vd5BVRuzGs7Rzru
St8a45nl6mk2I9ot6yP2nbYBxkgyAsM7et9U5FX38OtAPo7kKCwedfdoT7hdbMiD
OvJIRHrMwjyGJA5clMRkQ4UFMsrzuCqgy/Hceexs0wVzwqL0k+xTuSpwPaywVLRB
68roTTXUE6TQP2U3p0lwO9KGLuPFwoYUIxAJPWd0XksQF98ww//5Ep+5BMsF16z2
gcd5QcLHBiIMhqoXgvG3QMluZS+VELT5NkYc7YYkJfUQFn9iX8ilOK/IqWjabgvG
3LRUlzBHHI5TMBz9EEldeRim4ay9cB2jzPbDQzlO/qHD1KdNriJiUrtQMpbmFAjm
X6FoLMDieTYci3ktTdq+grW3+j8Q8GfR8/WjxLXCDRm7P7CB8PKEexDRPyalfyyh
evlbKdG4qhPys/My0XXUVKgyhLE21yGIYJIHVnpOqHfPDkFk7RQJaVvGTas9NDxI
EGWAFGjjmXRqgvJdBJ/g5rKSUn376kRIArz4GL2RZubbjpm8r3fCbF9OFD2jVkER
nHuqkRpGsvMAuwsLl2stJAeVO9sFlLQGrnOy26LPbDiMO9fZTRHhUZOASHvnKXO6
zgWd44AUoHCNhhR6Lci5MEzdU1ZbHYSaC2y2JLZTVJTUjG7+6zPul+5pVeqCogbB
JWpFsOxV0NtYSIeu5Nx6vX6K+uHSxqk9dcnNJolciFrCupmBt1wtrtDC2wyfY4xj
tRvIXT8pO2ve3rpTJMVWSXZRwOshtKy9i4c+cNfOUh4JQzOvdVJKSQnUtgTkxeT6
Blr5Vh4qvneRqzAJNnxbOBCoXHM2jILruwETrP1UxR8KTdrTxewUEWwnRdpru31M
2YjMdbTHppwrB3Oviq/FVFxCv6s1qwy9ePN3qYEh3mp98JXwQI6LTw+n9fqa+L2L
8F73oVwaM5K1zd97JL2fIJUXmSlKTK8X1+UXVZ1q9BMFmShp5I+Kqym4qFi1qNv+
quducJkROHxwj+6pqZ5Jo9kFp55GTP6zqFFdkXYLN6BCfc+9GQjdUSvUbAa+q2OG
M8fACOK5ma324OchO2zoHfexVBTaPtvl0f0ah7ydlzr5P4XYGy4QoSUiJo/nnrL4
oy5+c9Tjjst/p3OSFoSx7XhuAqB6+sjXTth8Vv1V55jQSsvm7Co25enWII9YN4je
1w3ix40HY5QeSk/F3PSZkpE5t+NYbPvTfOMJP5W9VdsMGQjziqyfz1k8YaJA+n4h
+CuODZX4+kizBFperkgwM0pjvIUlTl1vuQwSsBwY7QdD+CbJnNig7MOjMiPxWcVA
MXz1ssHKgzpoVi1i8gUIYAoPGgyr0nvO6degr69vdpPBkFZnzs2XVesOUHtyKnJ+
TFb3tdGgVDpm9TJMrDiPf0m/L9ggMunx/D6osiNxjIPBem7iYpoLthVo5Cs0bTRr
gTJzZ8RVQT5tyV//bd6Naqb0ELVVZywq2gDvC4qdd8Pio5H1O/Q02THHLU6k9Rhx
xDwYohoPPrv6YPwf5Qxjl8qrXBBXdu4xR/0m+egklCxMXf6n2NYlqQJPevQ/eGeM
02d9+u61gcCpQhjONEcYWrFcaqG7jtbh44FTHnOLQst1h9RtdAPJuurCv2WaRh3c
2OsbAqJy2rAiQfuSqnGTBHrYiRZckY8ah1u9s7vw94tO/VD2C/cOe30WlxbxCi2K
qE12rBLxRHnHDXXKfeNfppmiof5kzlLuH71nV/u1H/IednqJMZoBUaNN0ED1MFg3
i5TTdvh+8yFnl89fWrRJs6YNcZ7dnQ0fxkew1k0Ummc+nka1+N3U0X8a0V+nQCNO
H6lcPKVY5sSnukVRG/8ftsCuS/W3Qi7vz+YqhtsVgBUtvAawA0+lqSXbQ1z9v+vg
kGtwN58fstrH4jF+Y5dfJJ5setjN0GJpNuChZyP8xi8vgHWRSTJ4/e6V2HTZ6gOg
pcOdE6lSSws9vD9Ddiscv8TyoYIH6QOeH68Bzm6rMRZrtNAiNVLn1pJz1nJIJDCY
1IygJJAo5ddbnW9MuIqosx3xDpogVKqBOmhzhTghx3a9sN0F7SPgKjI6dZQCRtUi
Cb8nJxS0lc2R1675Lz5dKZNWflyRa9N5DuLkEiqzJ+8/ymXddJ0OUcH4ANX6g32v
GiIm26cgrJiY9jvuJzfdJgBNUdG93MfiBw5ucf5Qoe2/g1KPJzWW9waj2qej8zzP
7C9u9UX0TVlZK0/iGtJH1HcNahhnRkoHDalWTxEpP8GiPMvVCKL2ZW76r6BuSCpt
xcZU6mHfuUxlkDV77QG+8Y4cJCLH2NqbVx2nQOFjRAalenGmKUPfSfAG47o2g8/3
nyP5+CJDMibOCLswgvXtvcouxAg/GGgmIvyD1HnXT9HtU2I/S+QtQVhYoRZHsqK5
OgXH1mpYrjW11k/LgEJGDWsGOp4HRasIBCWDp2uPv4KvpfQYizRboR6C4jhu0Vcm
bvUg7HPZV15o/1eSKM6TaBnRLHt/uKaOTxymGs7wQ80geCRqugiXxzNJ522LIk/h
Cnpd4yMaE4YzpcAbG9yP4c9PQe/zivgrFyGzQedB5OwhTK7w3NrpA5sLlpOE+3oX
9e1++vyYrsBPILdhUuZxtWjrg1Le4mTMZ7wmgUgcpDhEw65X4L4Zghb83xFCS6Zt
xiYcFqKfbyQGLbqGeHd0XXWm0qATCUB6C45+px6dWLKOYCu8mzXdEu/tolaW71vJ
8TbgSO62sgWzisT2ln/8gd7GlueGcp2VUDsFxwd7IERLi0tdl3MBhrN6dwDQXA5g
Bg0ak8DzRYVbsuWwxU1wIIlYITELQlA5kYGTzqc1H2zzUSNUOoMYtNRo6giBvuJo
FMlhlKyOdYbpCMaKWxz5TM4BXhkUFu3kHediiI5/p7nzPXIcHkElgWQ+tfJLyzVV
MV3XJ3MfH60WEjs/+j62DXZYKz7bAobmd6iTcs+5cigIHWnq/2pBKgR2zDAlND0B
7p5hp1z8AtCcP0qn0QBZ45E/RAMOz3yjSol/E0mxmtjRMcrMhUapvF3AqVhxUhB4
SSlesQAE/UVYcwDWjODfyeGEo391gSuo+UVQ6XDn8K4+N5dNrBYUTeHJvZkt2zti
TOLbfP2TIgJQ5pNw/2ERGImx4Lg5jZNMLuyRSJUEnLx4FqZ2Xg5FzfpgUpFMQfKU
8taK/Y4+j1Zy2TyngXLLoqo09pZcuhIqmFYZBqTa9rYxpfy95867MpZIRcJNwNyf
X65OSjivjz4/lVgQ5aWa9yVZuc2LWABjJWBQ8mDwDzp6Yd6ERpvByMA8aEI3/VZL
6hqIwY59gD73/+pjuSFM/R1lVeB1g5H/BU1KV7EMpQCiVcpuj86IiWEkyjorhYC2
a3T48NBbSL2qkRTffd/qBldMsEzsNBuwUXIv0FBjGOMfiZFMc38dwWJFs0cpDNXL
DByl/qRNUw1eBHF3jOJRvwykkBpu7nL7EZa6VAeBs6nj5TXqXL/poYyez/jFOwgi
9HNkHGhVmp2On+VtKutINkbkCiiiX86/Dg0Nlqi2/nKUxRrrYL5mqrjk4eT42LXg
Iqbo7XrGb8td40lGPiQwYRCNbz6qxLyJJbNAdaGgJwEejseIsOgF44S3aHwc2oid
uDbcdNKovxVo2gvlLdbEBLHtkz0vLRs481xXypj731MMmK+UtliknQnXMlb+z8ee
NCKvlELvoxD9KIfltVYc4P0FvdoXMJahWSOvsYaHRQttWH9Tv6OQJ8wPeRClhArR
BHD4CgkVbzmrEJmaoQobOmsC2gnC7a67ffjIGQENV0oyySm5J9I/jqqjjFsFhjn0
OvRfDlYIZOW0+kkqi/MZx5xxio4Ot2audBERWs/MmSfWjgSbtZaEAkCWxxTDahYv
ChSBy9syJg+Gpbt8JDe5rxNN+SDAV52DgYyuA+2Sgy8Jz1Bo550CDjT8eX3FR4Yt
QEswzVeX9wbGWuBWs2PBPMURW9vqu3sCAQbUpzRlKhMvb3rOPbjFumpIk/BV2D83
bW1lHwNc5xP4fIrQUzatV63Et+6jT6srZcjelCtBdJhja7Jb1Yl/WoemkNbNlQ+9
SZYVdhr/iy6OU0DR4RoiuRuhmAu4aLGF7DhhANcnbhEsP5XAFkDrHyLT/ivVi6+8
ubZMpTfWfvfZoxYYUIq9eS7JrMkpBJ9gGH+EsakodsNwgbI6O/n+W23GxWbQvJM8
eNNhrWqWKdLM3FtbiWGKcw/Q1xMEFQwAEJsSrabhyu7qjxnHA41VzXyapy3bwVwQ
LRJgDiL3P+25uU7CCYYlQGV00F+JLpd8+W3UoHbJKp0NumevOBTNECJez7GVm1H8
NEsdyF0Yx0UPEbpjRjnIQh8hjff7M/jnoljyJPj9DNf7Lvd9Lz4c9Dskt5UGfpVa
J7ZNBPvdHccEhWnTWOaeLkXHMPVYfdLghuQDTTEDoKu96WXDN3ihM3gw0ANVPHkv
Z2lmJLwyANdJYQtj3KfwJZivCK7vrpHFJIP3hkmqOa8OK/j53Mvc13BLPxenk5xO
ZMuE5f7L/6++rF4txF3mErML2Zn56a6wnwpCiot/jmh6+Xv6YmdmwfoGCI0mKyQS
xAVbDFLsLxGiNuqGGR9XhvczzlBjGg3dmx7ksVBeBjsgHbyyPq4fVSDRR97wPE4v
fEdyX63ZtE4ZlhGAN3YGBGJnQdIAbnfcGZU5xX7RFoM6nif4AB4+EjYVt1DDfBn8
vbRlAyXyNbJL9xSQrmDJW1KgkGH/OX4DfAPRQ3Ynt9W4UEW8ujMay7SH2JYR2LPm
5InpuX6iPMvL+ce6tvx+SKfL0W7aojZf2a0IW2SMuuEfQWqV9q59QJ5WyA8cznqE
+9EbiMzMdBLSTOUnAHOrYM8ZRpwAY7SkTitLA4xh+gnDsSjY5NmoMCqbYByzHkga
Yi+D2ffWaQDv6IZ3IPHpUbLJt2CMJG/Tc3mMul3KI+2eYtz6+ggJBSBu0pTgMCX9
zOmkWvRhQZ2BmpE2Kt8wvjKQAWEpCdF0vqvTOTMkaTBfbBLTt7yzp1xeqApT3pXE
4ssdkkkCJlmkMsBWewuvhtzYtDRV6BktRGF2liV2k0Q+72nI+avKORNoQenQBUav
vvJII4liMtje0lnV5g8AKMm2HosnvOlS4ATtgcPfZDSObH9MJ55ODZtV9Q42ANtU
sqcnHKmLVFN7ebyWZEw7U5ahlZGfRqJKFBVQQXHu4kUxyEwvBoSKdUwkwk0X7n4s
v7qx4S5iVSSJyps4OrW071VpXzA46BUV/YX/jh3fkFNIimQgjXWDVZitSeDISKtN
nr8oRfu3XkEIrzUmKIJcbjBFMyTBCc1vaabDDRTeURmnRerFUdfWf4RHVld683Vz
AH+oUQWAlDgRxusNZKKGF8gOOlIMVsHIGVPKWt1vHVZoI2k9AdgWdtJg8MOcCwvn
jOjbmDnuI6wQN9N1TDIykV0nFPVe3Z6N1sPz8PDA2u/ILY3rwTYxvRr/3juhE+GW
s8W6qxNfxRwvtyDaGQFWO1mao/RcImWeB3+J6Qm+CiRGTs7MzUCDLjLSTnkdma94
CySaOroGArDKyg1GzxBYj3a7hXtgqRwv6NKR3qZIrCJWfCkyZsL4AKyXY2IQTBoL
1Zj/IayE7TfRXZN3jqyjZMgWTXfvWCgUjMLUStNrxTwOnTHe7J3k/q3jFNAJyEJn
Uz9AWWLOkreEFSOCQzRr+CALSwsFCEHyjSr5BFBPo7fexImQHb6n5WvFdUkCxH2L
0oogfqAY1gE26aswIwJBc+soEQ0B6E1vI/Us5vLRDjZBS9CPnA11hNiHgoVNW7/E
hGHmDJzYbwPq8tyn0Rcz5NQtXYZf3KRj8EarQ8n/0jBfAk/Dk67vJYb5/phXTf7n
JmtJDa74803l2gfMc7EEH3DPqI6D01YyOKLfxaQtPlekk3LtjagQkrvP8MhDKRbW
ILQTYfJeAs1uig8DO/yoV5Eud340z1YLTFA7oPIXJ0uPNcWczc0787VqGxY/lZNT
+8AI1qpPX1Wk2eNC9v6bW9z3Pw9/BJW5RB4PjPZugr5qHiAeqxpVp39qnsAdZFP7
h0UQP24wO7y6gdG7R35Wpref+r0rcNR/CDAEKbzGR2Q+DTDDMLMfLssUxe8Dghb0
o0dxnVinLpz+ijmAgMpwI1A9h6PPaqM3k3TK8y5eUwC0KC/PUeTnNRF5LL7pTZ8D
pdVDb6rKV17p8hLHtHuSxwXxlBr7JOALuvlEtL59DNrKzRjQtPF8pRCKLp/FHwLr
+x8ats6RuK0LPHv1j/bohGQXSeT+padPLTfkeRBjsln7E27xtfiMep3G8fkxKvV+
d6wZ/GB0ppKTGIgK3ZcVL30FRs4PX6Yq+LdZ7GG4B39LHccAttw6tT/vQbqxp3+v
krV9+NmlDg13Ih8szgQ5uJyiojlYo06iJINgnUWMA+ctCwPxnoutifZHCrOo43Tr
fd26j3hGOc/OexPTZq4m8R3aF0yL4rIbuuJAt+wojdbR6SJMU+r7Rej6NT0/BOH0
xib07LRYcGcU8nA+wIfItCTxSsnYWApGtM2KPvPJWuyCqMrNV/krUbh1Hmf/iaa6
RE/IoduYtDHy0RA0f97P3X1AiRRTFHbrSmvc0ZG1viUELzAhHa/EudEUaYEVfne1
3IVo+ig7dEUpWNRUta+eYZu7IOTjVASQkzrmR2a+dshWnnEdRYgyRqdb7+9fazE9
qAOmuScpITE7glBk7taao5YqoVKU7TdZ9mTk1+1XmYpCdGv7mldLEdP0EzwdAiQp
d5EmQDkslhkk9gRxlaqwJpDzukBkLwPMjoFRWLxnSS376x6H48Hv8WiOzQjEFwVn
gkOEvwxjY4MHEcjUQoHosTWenFYE5iv8VY1Fu0GQwJVn11BhHhPqzf7+ct9myK2g
Z3Sup+eSzJyKSXGMgIL/0DVwnPmNeQBeaxp5Iq2TP6SzdiS4VhK5ROacnk2Umd4u
kQsHj3jqVpErbQrhsfALLy4kRTzRxUyDqPmS7CN19+ashbtB2aYZcUImLLCJ9eWA
aWNJuimANIEKn1svRuTQKGbDjiVVk9/NAGRaPv2qy3eNDgNm9mRRmze5uhGw0yAX
Rm8E++DYM5ISaVFbcqXdLyB6NIudvXEMcLugbcFO/gzpTxzDXtaNIn9bpu05WNER
NNXoHXBeswHscI5pL1z1Q+L2dXFxHGBqHu/VQmMs22gAY+WmD+D5InKPUkJrOhFa
z909BlIHlXJEN+oCSCS6sbs/PfsYDub2tPByif7veawJzIDbhD6Aowkq8ntzCqhz
tZq8I9Wodq82t8af3KcpqDt27z2nGPXTq7PVP6OMjaQnFQ1ZO4KB4YhMTzI5T4bW
BElGqhi0d7KfF7lE0hP3bycNtrD+XEsJK9AIXepO3gocCCFz4U7D9+DGH8CjPZvr
zhqsd1UmlluxUdqV79rFCIoy8APZo0z2cNKYHooaMAsY99vQIl7YzkYqkykTQu65
c9pW9DjinKFBw1yHaBTbuuWOYN0apjTZdhq//Vl5jBQCGndpmRGFEQZdBMynkNsN
CzlD4+VoP4NhnDGMFkYjq+lOJi+fe8jaCWQxLtqsJf7d9UWMw9Na2ye0QLHgXhB2
VzhGl7IrWjobcVN1s5l3CMryLUD5ukj59l0jBFBnH9OWhxSMF1S8U4CEgXTLZb0d
gkx7u1fOak2KO9X49WUtjPJpNAAUy0Gq10MrwZ3lveY+b0/LfoJq/ciVdjSnOCby
CChbk1OkfqlFJYTKIlxEk4qCulCfjAH297mZT2rWHInR11vEyXb0vZpkB+nhGtz2
H5KXk6CJOlxvDaN7ZCTjSNxp6mdE3CnNqlZLc9UfAWXwn/2Aj4EEPoZ6qn9aa+Ky
5qFPfFodqVT5i9pvaXukOZ5s4VBZ/uVo9Fz3Eec1vdqCgwPFqwrhROAp57uMX8qo
Skz23yw+vNNexTq81zRu2M08pEonN6iLJJE112uKOCd1rfqIsuFgssKoCVdPKypU
vXJzTJgIzKeqXFY4j7wj6d49eyGqOXUkOy7w0py6X9RJnEqzGgOJmFGcYelLpQjW
UVqBs568Nn8Bx2iore984iv5R08JzAAVSTd8da2ugtQmOq5o1j68zYzhRGKqIGF2
wDq1LPloAWVRTMCIAjxL0+H9H0XLGOmVBQ9smCz2TImQ1wH9WRUEmCP2ABnlY+c3
7CfbCYye6F2ELg46LCY7ispCJgXAom9viTaKHKLHPryI96JbJI+Ana7VIfklMRsX
3QacUfx3HzN5KfCRLVCoGWC5wyMgStCtu1T/mWt3h7jqQhJIlyvX8DxW5vdXQpSc
af3ECg941nZdkoJRGKIORoZYG9HCas+rB+4yrZNr4h4MBfbn2KYLvzSwclvRnmAm
WXJyArcU+tmuReyasQSzLW1DOVwS3Ma7vLDpHInmtNRzfJHxaLZeNYkI+Ojt0GIE
xuF08PP9BtxcwomBi+IwmsQ4EY1gY80lClN6e/wr+3qE5AYa8pG+Yp/0Va+zuv37
eOILapVcOD9UwxWevOypSnOlhS1U50Bxf/YxeXtNpOzC9LNuPhUzDnL9O5RS8ZBS
32quZmGOe3J+aP4mXgmYc6K8jqECM11nm112V/Mgsvl28IK3++UtxqElmZI+1xrC
6KjuwaEo87OtGyWJjgZb/IWHHpV8+IX29uzcbog45deQrwvqZ8c9pSfafE3joTsb
utY9Z0PSHEzRICk0YZTJfxbYD33boVxKEwTz7xW5OynCD8CfIPLC3Od1oufUkYbn
HjZSQKC7M09PDEcUjMVmUzUmZyXxPyNrWC9McmrLz84Oks0ff4JAhHtHiux4cHGI
pdqotOpiKmdT1mDj9ElU+txSiKTqktkaKl+25CdtThbjOnQbBCLGe9lPKnfDQ7fN
nCuOarBu1Y47HXc77VtsDXb3cJAuGw7odsNTJXy3U4Y5YGMkKEtlBDhmtxp9SQfq
IHO6STZgzENlGu42EYdJKFkF7NBHzSbz2hAZ4vBLNjZT81trsr49UJn1CmKfvWE4
dHIa/aO/tmWEiWIu05r9c2skX3WNwZFhLLXhhXHSrwgH/H/ecRXY8dWFu7xkEN8y
eH65XWbYWhpzD+MzrzCO90YGwkiHBbTqTZFVEKE6u/6AB4NC8I8hb5MPf54FbygN
CMT7nVXLpgKod52UIGFG30ndn9RgA92Ret7IOIXFWYtWB3qBJuBhZrsbGcRyJzPc
Kdwrd40bHHqpLBjgVF7p+HSj2DFDulQGd8lhVbzmKZ76cT5D1HOyTd9sKeLa+Vqo
nLA2B1o6QgkzAqyAlUu4NzbCVygkTRogNlYqe1ocgglyqAaRkIxTu7Gg1ZGfxNgR
+ZMGnmCylk4+nH67Ja2ONKwzIkcYdBcFKqUCohQQRMfMEsl9caKJnuhfR68Gr15s
vHSQTTuKGidRvzbTp8K+NPSl+uXyAYYWjXBACBx8u33qhpwIrvFYnx2QQy1p9OQV
DDTKeocHr27X52feFqRsyKLNxEi5b08IWHky5Qf99Wqq046lsAVetUBVeMm7ikpr
y9BjJWJX7hWtQSyCf2qJy6Sjw300bOJh3+S4+7JCazkPUSCqrcBrokTEk99/1muc
2/vdM5gjEPOp8VT2wEB3qwawDc0ZeC6s1Qk7nHRMrQDxuu4+oFo98zvKbNR5sR2n
iZf49akUF5RpFKwd5K+jDo0O+r4FjJGrqE92y9OzqZdYVEJXxTe1BIg3N9i4I2PH
bKjGeeBNlG7htl983m1d6Y8hE1ad3a3Fl4kMXt5ncpxIFcSLb/ze2dQ64uo2Xs7u
Xbu3VCo42J1/nI4ujfPATRRt98wXukpszaOvkvbPhzxAD7nNmQQjOHW1vejdeaUq
GfDJFtdn+EeLgJuuZFyUxIlkyDdw23uOboxDaYNIFCnLY/Gf6k9BPJjRilTJR6/V
0SttSIPs3O9t5MQcHIgb7WWfFijKPXYm3QXcuJshIm91G7QIzn1WgNnWzB6aWa8/
Q2wnulZCECuItJYuLI/Ll6NRTDBLrFVI41Dm7h/4/2whL96ofvIzlCmwI1GcVpFT
CRXwlHR5I8RM3xanEAlHei2dkELUEbzlrr1/4/EARUKzxpDlo8bgpIpaYAGw+am9
e70TpuJyn2sapEO4IZne3jWKQ5+mr2rNGqujm4zerEy68cASLoTWSaJEBdq8z7uq
ktnJz3+EXNffF/usavXpT2gdRDGJLtNGHBI7EHIoSESFQNVjh+EymjGXjH7MAQII
MQ36ZQtpqBFG7VJkuMUuHgBM35/L47liD4Yuk5REK2DTFiRyTrXIVYi6WsNDvG5U
GdX/bYlFZdZ8nqXe93EYB4fSICydpRiCyCrPP8PXEtzrljUo6IhfKjUu4XeQvITv
0P/8KVPZNC2koLcnsN7RZhgstmW4nOFPdlAnjfKH87aqk+Wf6IE0In1/qgrbpwBg
HeYrvz+uYIneYRot0D10TAefK1K4mKpZpERnkoc4bipflI+fBd4hzgUIw6D5R6RQ
uiuCYnuJGb198RXsUxyMcttEUidV+QH6QpxUMcu/e4c2w2iVIOaFw+Rxs0hiPiaz
hsSbvVP6ZsNdEbW+ocrxKaTpNWo1a2Sd1SCiwtdLy82OSeaTMR9B8ZEHh7DpjUrt
8V47l3YxtKa16TNKKTzXRw+JfIA1/VKa4+ZeBofW3p9bXBCn8KEuDxSgIl66wALv
ylKBS7AX8W8FZOnFaJI1YEJKKBdA+WQdsnRbKy5rX//Ct1lNx4u/vTfbcw+OqZU9
laWJW/iNmNszNyISCRlwVZCH5NMx3td5unbAyZCw6FbAI72UjMlSEBgdtcUC6KFI
uKtpWVu7ineeAxn8vnKbMacALPXlzOu+x2ljOwgvhKzXujYaBsZaFShjMDMqMJ20
l6XnaWpe6sB8LDYKHmBMeRfaFK0IF6kGy6aqap/w6vtgfF6Ylcl7u8Q8wt68n0x6
Lwuw4DXPW4l1TesocmazM4z4sAH6bgJRVMvoZewHpxEWAZ5t0ANCLxsf5I5UTbY+
TNhIZnvUhYanyhgCdzcTyIqQz64Isa4v4KHL+ddyVUXRkwaRLRPnFrZXtAtB9oNN
5RVj4+eRs4IV2C+mikMhCKh39P4ZrjnkctWvFR4K++q6WQ0OW9Pw9N/1BoG3dmSL
zLyejVMlE9mInKckYCCZauvAoMBdI28dixcjjoATkVxr5qcnZ1LkSJjH0Mqcv4aJ
IB5+hoKj50JA6wmuB9HOqml+BCMGvfN+8Eccvnl2D6/hr+Qjnx0cjVuhJ74OIO8g
+XIWiX30Fldn6Y3rnRKx73rPLUKy2sXTNjcqxb86CGNKBHaYA1iUAM5lnRGXs1Ol
gATmPG9e7cbwMQJiQyV5YlF13sVRjL0YEhLau3mSXJoGKtdiIFi6ed+qHuKUr3iM
quD0rCvZlzUibKogGdyEKebi0RufIWiXLIA7DixhlLmdsBLxayqCnCA7cWD6gcLR
wCiRZ/tdsaemxJ/JAmpDZlxD9xf7u8u4xghol8J86DTr6beC6w6/9lx29TIcfr+Y
fiGGri1jIEIqn2m0xP4aw9aU1tGvzqw2W0+rMQG6f1t/VVNvsEURrnc6q15wvLk0
dzB3pdbAi903gJDFumeCKMl36UMfgL15gnafF9Vizt8gN++TWD514MAmeJPkfH0N
m6fLZD70t7ZTaSrYeg5m4gF757LnR0usJ3TXrcf37zwmGAcvjDpK9cb9/6fdWLY2
HUWH2guddMNeiPXTjJRSJ6pSkwtLN/8sSt3gaYVC+trrrsW5a/v9DYJWns0l8vdX
2AzYC2j700LpkX2L58kuZprkjHVInzUMaopFjGOyNn0YoC89+wcjcouqXCUva+sP
ohfnbamTPNLKmt6hKVcvzloikyBjrSuZ9JbOs9vbfv+erh4B1AXeb9GiiUYSk3Mz
jyCKsnQZbC8ZICWy7VJpRpyYT2nU9eS4dyOhidqwm5yeVf8BxEbTgLyMDEkR9oWp
/ffmRpn2wVqbN6dBAmpbljnBestaA9EUDtvSDOgCF52PU8YuZroa9gxdsLDt4lOL
j+EEkf1BucKEFLHmYuiKyph9kAmSzs/fsl5YDMrDdF/nRLA8AcyC0n17dv37yKSj
v8+5Wpe9kalAQGuc0Mfa88Nt2ldiZA+u5yYe+Gm/x3JWDYC6HIU/+aS8QDmrJztX
ZQ+tGwJG9m7nqmm1/eRGCaI4J14d73o8sMUIC2IQZSzsAMf14xM3To9Ml46Wp5iG
Z2zNZR2KRcR4X8GvGZzY8l9BSezVlcNqG6TzAlNVaYl1j4bm+dcPilNbsJVS7GeL
wG65cbvFC/w5U/A2N51B58KfsrjKT8l03QYqUIEbUiKGKHeF5NaWPrAjT37cl0/g
zMqPAT3IGEq5+sfncnsRb4E8ok8ZAuoqEkrQLWeQ2b2kkJLDIeUCSpZ0UAXeLolJ
ypfjUg6K+DVNaEMdRk5/Oa5/Cvf0QixtFawW/gxwUURjWRWkXetI2p4h83BfNONz
G0HWsbWqPLFvBZ4jbrqeIokr7cNofhyKBks7PNX5gDa+Dc9DXNaE7eeHLlfyE5lj
K1BiYFW/QeCnFnLIu8ME81N7g3tH79qmGuCubG7AE95BcnhmbvQ0oaTq9jZ2ayA9
p50/H+mbFsemgrZaTS3THo108y6/iwgG6CcBWyL1g463BhMhk5jaBYVuAnhXhbmC
qc5bVJ54vcDObk2S9bdM8KMtNNR4A5e6hIpNM8wzlY5zEwWYFQ2F+nI4svccy760
liSeX7PqluxT+aWs3AD19r2DCEgcD40xfg/JqK4imOZbQQUZKLqZtqOx50gL9j/d
jGs/PtQ80e1eADgaXNZeMSmtj/BcENNk7JjSRjTqaYNhvjvYok/fTASjNyiWJY3l
TtMXOTCmfwJqju92Yqjx5SEL//gVB9RTNboJfDgx6Sut0+mlu3IABhxs9LBw5Grg
r1b0y3QkbQW5n0zLlQrodAnsScl2V64AEL8UYRcdMD62L1jtJcssCYhQXsk6ObSp
7Qq1mOPH0N/GubGb4rsMOZDKgU4srph8E3l2ieR6U3wIFKDCMPm5CrbrShRZnXX/
Q4jICNAPxUorOo7Oq91eolSO8AU0iyGSF5ZIAaFto1BljFwjLYw0WFnpCftxl5p6
1y37+FXgkEt8IYorbOVu3Tb7HRaaMH1/63TMEl20qCUmpZS7UqO5DHwHu/rSzXrz
dGbYDbQx3PpwqUstNnAZkNPTVCvIgcRFD/xivlPvRK14vN33vr+pCZjJKNC1CWHP
t/49DUDQ+M7t4sJSoHwQUDYQF18cDT/4KI0grV954hrZzDDr7ZTSoox9x0AXKvwb
N1LfVA5KLmBa9dZfRHUXd7WE7PjX2wHA/+2Kw+NOyGJ+BFocd7MUrrYo1h6NyGm6
8CNLleeAxDICv1uejOrT3/3R9/Zk0LZRrkqv6+GYcOcEg73PTCXeH5pPFI7CoSkq
LOQIOOfrEBvEm194n9nkiJ4cgQjTnHj7O08O+/65DffiakiGF8XsvLckGnYLwGRD
nYtVzyaE54SdkepAxM+JG0sO1Fk/QGK5BXFUPdWww2CBG1u296Sg9s6bAWE6YtzO
Nh4kbk69y1+DULiag3stjrrlMLUzg4i8XWBDkI2YKmQz43s6Hiyyu9o5y1HFIbW6
NAfgTU9xlYB2wqQ+yf9HWNhjpoWF5arJHUoFw6LO6BqfZ4Wgysdb3q1kaqnkSdvn
w4mVAnyopEPp6CIugUJSwd0evxum5oJ37b7b6U1XtJuT/UPFN373zHhR7Mdvh7Ac
aZwFQlX70AYqnGfTLzQN3nC7AodnKjNVOnzy1CwPYqvjv8Cd6yi3Lq+feT5NcTU0
lzNOR6QPjDyJpTgx5rnBJtJIyQUUK9MWma9C4/2aBTUjXrpxdjYoYnp4H+1KR+Kz
O9O2OngHoZqA3d+NSjPq/XuNhD8ScwiXGWzXyxjffgCeow9DKCE7z7Pag/U8w7Bm
M57FG/CCRGLf1TXcKoLj8NCGYWvkD2hnvtIazFzlE379Bgf27unPejOIfBGN4X04
z7Ou4VLINUec3wEexP7XFQGoXg57HHE+vTV8dWKHMkNqcAp/wvJwcqC0rf49jvtc
l/0F0wNusdRsR/2gNChw5PwMyga0WcdAzkxyXuL+J2cNkWQQ2Fknd7JuvE7fE/XB
8p1H/54sio9zExCfTOxN5pCKidXbiS5unYmTeiYQHSS1fqx8TxsBAtepxVCMZMGb
a9iYu2S213MBO+aBUrfLTk5v2f6aJAPbvpx8wLQkREFcpRWo7Zi60nP9FBcrxKHT
m44R2dToYvufWaKLnmZnUQltdC9/xRFX1CvWI8799AMeEdlgLnlHqHrIAHvBYSIh
kkTXt1Meuz1Tm5sE8ezwa5hvoF5QQtbLbCJeb9FVMjZF7VCeo52blCQ4uciJvz+9
+TETMvCbwI364pl0q1xrMy87xS/bTaCvSBIgNYynn9Gds1t028yudEvZaHr2nebT
V6GgO0he1TnVdJhdFgUu82sHsn7Rk8QKq/QJ8JEcyZCbvF/uh7FmnirUrtYiwuq4
vy04Gjzfb5BxGSsF+ApAu+jaba3tgNchwwBShh1gmJ/9dAIZ0EEHj0eQRp6bNI2C
GJc5JZj05OAYfpgMzy3nNtqZfx2bosaGHJQVUu9s9ypcvc1loe1ZRMfHmqD7PQSt
v/PS/NWF/SyQaMEkkVXIkgor1mzLXBz3nSfkSSy2Ahp+IM75BkYkow5Jh/Poh7Wz
IaouWuKygDbjhEjON8VSTIyP7cvWDZMu22yOKcLr04KCklNSYvr+mSyr9Czk1EBz
58+5maMJEV77jG/zmhfkfcWLtGqwgacw0eo1TEw8j6UR8akOpXiQQRYzlknp9MmR
FyypGWfCdyl2UE80wfg5Ow6qpqOM6XFuT0RGtetCjGddr8O1ERyJGwPYfq7Bz72x
+lxQMgS0WNivaDp5dZPifuIBD2RCrUEtMvKL9LoljniKacU+6v33LZAB593V6Mh8
u8XUYPFmqz8EfINQTsWYKE96w5IJBgFDAuZQM1k9Dny8ECy5f1CQ1+4w4WgLMvEp
lslzDIy16YVmZd/caZl9OTVLtv2lf4sCLi/uQ9rFksMm3QbUvUxz1i12gfQKeRZg
J6f/GvDAGZOTq0WbeIxUoZTbndhV79tO54idLnys4FadIKgjlDNypWQ+eYZpm/X2
Gcsg8ppAhmDbglr8/UaA0VpG5J4l4rwi8yZPl/9vjOYusCTOZq5HWJFJqiE8q1gz
RgG6T/aDSalqHR3Vt0J2pca+mHU9U29+lwZeSg92hO//EIN8ArN9quGr9h077QTd
KukFi5XQWFhFAN3xaLdHaHNOY+ueH+d4SlpiuMeQsu8wDkOo0GiLAcFk+A7UsCSq
4atjXXfDlXyVXTwL0Bh+vElJRepcfSk9+SAyBr4tz+ld5sfsDGvRDXoAtobDKZcn
eM5+VP6vIeDBWxjcbtwYfpnd0aJUnkI1HBjifbwoN3CY7UD3cAtyT6Pv3ZGvcYbb
WigKYfjJa4rQH/cQ6gI6rE6g7MYyPO6ihYkyueyVhDO+kxOY47fHVJFZkp1Qje8o
OLHI2566+iiA/CTrx0l4jHz/jAp4A8Am2TXLHI5ut7qPhtPk921uIjTI6OmybReI
fEh1exSkwALDN8Q9XCcSaWq2tzzci8w4HvlOr4lLH3ny0IULGwUwZPFdx5r5DlkX
2zDJe4YwOLGrjRwE58E/6r+dHjF7hlapJNSGXKiMYMvvYl1txtL9LyiKD/Dd7Y2F
hz3mtolm3AoGVhz5otoVZaBZxYjucZbubKUKl5ZIGseV0VfN9hjAwjExLPRc94Ec
vMsZEsdTN+9FbSjiXWhc3BMS1R/1xe/Mkg+guhtiAiz5hXL/wLTOSil+9IEnnO6/
7nSsu0SF+uO/6Ldn9D2jCFfB71FrGqKjFQhPOgu/tC+n/FKGxHH6t7dDVDa1z0Dh
KH2kmdZxtjKmOrRRugIeuTfWjicZswYDJMpffGtrBzo1Wl0io/D2A+QiJC878G9R
byiAiaHsHgS+sSxt6ZVIY3Gr6ZcXC4RosqL/8j43KoTachV63RIIXPWz6t4KESKU
Zcfet3M2oKEyPySa3DI+1PtlsqQQo5IdchsXxtozX8Q58/+3VakHtVttHJTh7YA1
seWd6vgS14aeNnykkhwZK/cNOLVWOO5kxe/BkiXmoCLa1CQPVwvxRvHYFMzlDKOh
Wuq6nQiAc32JoU/d0PYEiHHsb6jyXMECrofy0zK+JZv3cCGLxbTJ/qCuoiMRUkQp
rXB81CDhCeSqqb3m6go8Nzv6iReeU3EJcuzYrCsFjc/gIkgowvUw9jdUj/wqD6on
63HtwlwvD48leJmxCpq+4PvNfcN24zy/y+al8Dx3Z1q/iIRwcI+juLDp846VN/sO
khRsFaYpK67J2B7/BBRpOQ7XRZAub0L4i6Z6YMasXd91sxb0GouO68nyvE8LTW0H
rMwVbeI16L5Cems1EjOJ6CDYXM/CUavEIxpWMmOsv8gOjK9V1VXWjqJ71yJ4Xgvq
f6UOJIdH8oMDB0ouVnQL1zVBUr2PZ0Oz7opgWCzuebc3uIc9E8SjdeKzBNd3hs4C
MQpx5+8CH/kGgF40rPs9Vg+mrlxOujS+nu91OTXp4z9dA+ieh29NrXxQzUFbOs6j
WsG9r0HR0eXt9hc7e8NgeOpB8Yhb5U6NDk/l/53YtSuWn81vKc8FKVyHQ0SgmVRR
4D/0YDKsnKZUoOQ0A1ZMhqdY9YGGZrBkXeW9pX0Tx8uOPszqmS118Rxo13yec4yv
eEhrxGfEpidQtEBC1UuQvIqL2/O9qjYxiEPw9FC1cHj5VaunT7be0S4gNkb3NkfY
rDz4h0ZBLPo2lxSOfF3+6qxdSiWyzpaRYCOaU1Q/oi88/NZguMvvFvoU+GrrVm3H
C69qNk28LTeMzyjZZXNIATKfOGSq231Jc/55Z9oxW3ThFlBwZZEwe9zAFclYXDgq
dA7HLLigkZDSVjnR2SogAa/xpTkSV2afat74oINjLhBiBoAtk9sALs30RODHmTmS
5qH6Pdiq8ukJaPwXfVMt0vgCz96YP8ARmC21opYpxpBwzunt/9/ZFKzJS9zHA6vT
FJslRntlxqf2s2KKMUHAL5xuhj/s46uJTESv8P4Y00jbeYE+hLQJtvgUL0uEdRt4
/oj9UKR/weWrGKtbIY3aewKbVR7bmPiQmzAyhBSDG9M8HkV8/DPO17EUOT7ar/R+
OGzD5mYlirffFYBRzF0usmgynOdFo8/Y66TLy08FN/anw00H5VwYKIePdeSCldw+
BQXewKvlixbftmPoiBDB2QH3uYbVm4PYZ0Nyqw2jvuBbaxv6m0ELdEmW/tAf1C5g
Rf7d79CBzjOyMbWX14S6Um//jW5cInOoYssLSqyQcj/s3KWLfNrUlAIaF4CTDmdZ
ef2hGLOh8Jr/TbGumds7Ppfb982Q8iC3EIa9gj7xJT6wHycsLa72t78dO4czyrPs
CbShbM2Hkjjt8pBuKMqomkXMABY1lUrwcw+FDXYer3mRhD1PvhnhgEQBGzkTPIEx
LuXwmzVwv0bQelbC1mBeo/APLggM9IzVK26vSkuljo32jwVR8GRAalt8W0pOSSar
+22me4uoeP2aTNXinN+qRZtusgq4G4bOiNjRR6bXF3LReGHshRpdnz4W9/+9f+/Q
iK/ZEieLP759wdL0udZi1mtVsxr5C4uT4mUwlBiNVaf9VQ681se7EwZehf8RyoVt
M/ddboK5Bj7IxHJcaVrFVsaVNPtWPB3NWMXnHpxk+wQ4llwRSEYeFymx3BF/VZwF
gcjoZceUSZyhNkEhSDgtQp8w16I2+SZs6UQ5hsBpK7wUWxby1M1JRulATUgH9MQL
S7uKcfw5hEkTEziDtzQ4WKuWjZSSYT1TO57aXQBxE5JSB6R9dV5V9poUGPNvBSq1
MmwoDNfrqqtTUPe3AksJ2a0nFHdvDy4rUWphWiqCQ8KXUVgJ4Z9L84hLmchZXpNu
PpeqnlnDdTmfNt36icgIEELOixjde7ecUtlkRuQyxgeF4d6v01A9/EwwpCC6UghX
VbugHUkgW69FeDycGjFOuzCzPgTbJPROvbLimmEV2NaxJpMp6w/1NpxhaG/tqWH/
ykBwRO4U5DjY0iKJh/Gf9g53OxJ+21oKLP/LiBSPSG0zse7LK1EG2M/TSsdASbVv
b19CAmSqkfJoSh0foJgI4K9JVvPzj/f41bA32/tCNbmCY8iuWQYo85+JmcgImoNo
/iAAqL7TpNSS6To/TTBd7Bxw3nwly6y882WLxKwvYMkCSTkTYawcndSSxlew950P
sdZSJM6eYPkyHwvrFPTIXlhL9pZHKePN/04pZjHl1EJGSOyPlag3cqMTRlr9B9Ic
8Gyb6LVcJdMNuWi5LMDSKju7CXsiGMKDkXIFCZBviDzxirQDm14FcHi9n0vhG0Bu
rmLh/DQQJs9xt6EAMWWo0ZkP0tM4WDs+hnq2hKmHW3YA5tJGn7IvFoYoDVEvOu22
VvGL53MaWQ4BSNetvi/bxZYxwn21+WGr/UmEXL9SOfmt0sUfOGz8Cao2uKoYqAAH
msZ2P9V7X1BQTB47YftEm+IY18C9bHc2Pg8zJ4yIJtJKiqwL9Ks0T29BM2fIpUGv
pxfQyDo5gPCNb6b2PflkGj119sK4x/B83yFistEpkEdG22bai9NVRyh0yDhuVOUG
BbBGoj6T3z0tv6i0xa5o5NcHvwiNhEna8XFgLY70dlGN2jPisgC1exs65qgZV3Wd
VhkswbrXc0akKTa9vXJW8CyBe5J3hJWSl68xVCUWObmS56V+zhgMcj3lGcSW4RHM
R/KnHi8OhhPNk6aj1g9RcXnLiPEH50XIsuqxCjbxoFF9S6rqGrMWyeC3Vw3no0rp
6gqSgnZinvOct1how/3qmaicZD/kp7Skkti9/P+rdB4qTdp0kWR2lOOJGIPap6Qt
VfzggDXt9U8ZXtSucREeEcKp62+egGVKuUZ8Z1qEXseaGO9/jJUXTsG4bVzSFUQu
R0i5J+OHElMPwTf1etf6z3iRKXlUip1a65nK504FCTNGf2j0UEUAJZWZogf0RfwF
xZWiUHjPje0xjB+s+7liy3BkahLdAuCKxQueQiIDOOASZnK4otFDmzFhGiT3vJDG
dr//yU7YbvGeNk5JciSkYQY0IjOdL3SJesFkSmoDE5t52ZSbKz8/u6/EvMhU2eCa
Cm645XVd9vgP4NQ2iURLPNFf7nMhCK7Jq1mkClFy3xuHNVa1tE3gEl1IBXQu8ZyS
Jk6d3FM0tNVwDh+oJQQ3IR9pvAmQSDuZr3b+/Dm+4kYL22kAbyUN9D8o4gsCjzH6
Cly614gN9kCb9CZ5u6sRvhqFOPrxfsbJ/5YEVIXDCsBpqOH0SfDeZ/pS6DoT16hG
oCuK8T5dBRdyplOBRpIgYq66l4nozl80NBdOgFwFPqOlMXWc1DgqoeWIJtBI1KV2
Ds977dbqWOlqAY8+vlMh1hBa7Bmq8bwaD8tEjxFaSLGMw35i3Ai1DavfnoliFjPR
W/TvCa3yvnhwa6Y6reoRkj+bbAm1+VxtukTKsActT4nHgVFp7xa7mrklw8cBW3Lz
liCI286LjD6R3UZIG/SE42OXrGHTfubKXCP0xw5KUAHjJn0CJNicjBdR2p05gqGv
u/7fOVP60dcYuketuALHID5qmnxVZmbo8RszHOm2rKEnPKimqiLkNMvZQ8OmRcGz
tqaw5EKHVo5raB6hWCbUwLSsxIVEQXlP6aOT2eK6HAej07TRWc9tw4U81Osl+2ZI
HIfU8lEMq/RJ13OOZlQ2aUIJcneMxoOnkBdKadP07Z4lO/DoAUUH8G7k6s/KZ2Mf
8O3PaAGQA57rqxmZes1qQhyw0YJSRmAFBmw6mZ3n5TI1w8FokCr6dE6hQyRnqrpg
BAfu6ELr6AnpynaP9tTuzeH/3D7JIheHj/jIspil/KhLNY5lk99sgZ3aBmU0ytx7
FejfXdLpF55F2YFIACyqadr0Gt66dhyOs2PD+cDzMk5CrWup5GoClMvm1wYRyF4Q
+zux1OYhlv+XZV77v7hKN8B+kOkD8JBrL93T/5+bUSu3lDjsSqPu+Z7Kd9F0vGJB
fFhrQkDhSnEC4s+fTrXXqIe8WXrbaPO+HdZvVUUP4iko8dEZrbBQlmarrSZlvp+q
4cPXIk+bqcXyiIauZbsWBr1J+geIer2fKwjwALhY/KXNsLFxq23NeweOoa3vJi29
ngc4RxDVGkQnAOkR0+tMG9aKGtklI8AhJSRfgPzLq5dIMWCuepLrPHrnmxHZPQre
vWFaktuf1n+33XJmzc+oFppE3LfdqM1pm2wBfK4rjfFB2yOKObG35DbIKqsuzw2a
3p0u1DSSKG5iR9TRRaQnabsLBjoAvTNeSDOzK+Vh6+Nb9engK2coyItfeWHZ8L/U
Zh8N9ouWzkyYfgP7YimVTCOlCTWt9U6rFrV/Y+OC3sFcEpxhI9dKVqygvHsADqtn
MMNnOYd4JWTlLywj+GTe4nHNWoPO0Z57GwHCIwbXtXdVckEjk0wFyNeqRutR9Ky0
Ej/r/dYk1i2GFRbPYAjza2TblMk8fZapO4w92wmeLZnLaxSZFVFcnp+4NQURZy2L
IUGiUejw0N962Ryx2OOo6SWpOgQepgRZIFyV7bkbe77PGdCkdKH4ZdJs5JC2h7Oz
En9GihhGdy87OzFDtDvgqtQlcv2CwQ+50utjFL3VDlr1mTyHszrv+kZ5SrEDkolo
VFHwoMxApWvM8YiKQvDqIqKVoI0xtYd+PIxEQbif++PtV9EhXRLsBNfZUCHYbqn3
9ws1DxnOr4azeZzMAAe3OsHgR6N2wcBT367cKi6LQuxuA0trBeOM90exYQOLFqYt
7IQajWE5Yj/YHgZf+bI3ezkBKcqED247cA72aM38uICFOPWxpAo6oRXYhxehPM2U
l5/niVVXRRXtpNg+ag14Rwedh91oOyPwK9mP8OGdBXYL8vRBlcC/wX4muzZgiEBm
qHdfp1blTAf9uF2keqdVuHBS5ykUx7R1IWJoJ5wD3/4d1ZqxHNDGN8ngbIgmAw0t
N8743cmVqkBZc90gajwV32tEnP6ACxcfwE1N38yhEMvYyU9bGeY2u5KIJesH69pB
wW+wTh7ZZofsky/p1xW6MLY2Tv8eNUS2iaQbbgEluqNrSY1ib8pAYfbUuNngz8/k
nJErx0jcVyK0LRlYVWLQkcuHQUo/HcJq4HSif/OUm1j6duzgz5sbv6d+ghuC4d2F
tTnKOR2r0NVtzv7M/pAxxdymEGhRsMw0ViDnP56ZAi/lfV25jFoKif4ifDuusHpu
y2FDRv3Cp+3FI4VVLWlevIIRAUgp26BlUc1etIxW2ffRUHIYuD1qxSxlXtcEpBES
ukZcAj9nA3VierQnZcOhuXRwZEDaHqEcL99N8aIMoTMvH4P1t6ZI24/+4ftRn4Xv
Aa7EF2Yov5H1cdilYO3a9YEfe1m+PmgGGxAfuhJMayJEPCIMJTBMx6LZpdjlRQP8
QLnE219ftPbnJbZYF7J980dAkMdvTP0+a86ikunnmcpQjyLrWy8ThLRTCu/vJIPU
Rv9IjsBNtexxBGfWOY74Xew+GtVLEiUSbKuBgrTgIZSedojlhF+zuKqQuFpBYGOV
lwifq92Czcioj7wQzPVjhjvJzfnj1ckIXKlRoWc6VX4gLP4exhOIloPhFy2BbXti
3+ShMN4VjyPSEzU79zdNnj2ype7B8q6ejPOarSgeDntdTR4rn7UQoibw32uWkAQF
IM3RWlYoh6K+i1ZpoU32K8E2DL54lwvM5m+2r+h+4WqPqEAZ2sJ9Ml6D4RAo2pxF
GfE5TwypBUxJuNumb4R1dQZgi6mTEMr3wT7yAt7v8Qwobi0P9atB1Yz5C0kje8mH
9vhg6PBpiSqdiCefGh29exweV8mzn/GVbZLYmSYg7Z4mozeiK4btDkZgWB6Ec5RW
kd60g8eqBIszSAm4nxIOS9qTK8oGGZ1gThyfKngzCX0cO7hdQY7sqZhpsCfzHsos
Xs4uAQB+S/KTF8ZFIBVZWaRQcC+cW+VlPdQfKlcAXE8qN9LaCVqQZQWerMFmpp1U
uKoppQFvF+n9Da+tAb/9ozmLWxY2p6+b+gfKQRaKETxm7Mo0KxZVYFOYjK2nyWQD
Zn1Cy/n/KGxRFGby17Tc0jFyNstxP+rhH1BQFyNdgIELi2y3KbjMcJWxdmyJ8w5t
QYqKUT1ng5X134mJhsqvSD6/eTIBw+eMKKdtJUbyUrl/9NtLOuWT+3+XcI5ZDM5F
q6OZy1B5YuXFfU27aLgjYsuyTIFdjgwWRNr85cDoEG0TCYE98dhzROfxZTUZlFkT
zMl5QhdP4wM9uqr5biyojj1gh1lPHia6jeG9FeJkNYJmUQNwJBkmCAFijPLc+Pk9
I8RFjsGdizNAG+RIiyToZfixIvN9h+dMgSA0OOA9xJH13EqEPcHu1RZz9tpWI1QD
uHbsYCP5QZo0/dE0zKYUzNkzKuboa93L9VboXBnfiA0UkK36MKGPdlUA1DsgFXYc
9/DIaVauSi3aU+4kBpbjwAB89djp/nzrrTQZFn+Wwcy+NUKHmNEIHXL60fLhEKNl
hB+QoYayDqgioDAs2NGgRrQWpedhFEHxnYl1fo0FDs5TPEv1Wad400tM8CJIZBlI
/9HdZSbxdYMXRx2AD3V8GguKADg9SZvrKKOiL7Xl2cPyOlbGByCSEz9vJEUw81GU
LQwCgJdxYmIycp4n/RtKMIkDJ22vVU3vxroFqxNuXQS5LowOb8tDqoaAD+8smJEZ
SRVA0oAv7j2gndGX59rZEEDqjl7MQOqUbfoHPpvM6qEEo38elzTmIDvK7fT3yNOX
eyqDLz8rXsoW2YQcWcfqkb+PblKjco0k3+9/fnOiyMz2TFeaTpHuGsuYeEhFE/EK
DYByRTxYwXSP+uO5pAb9YsMYz/PoFdGkw1rBTDC58fw4g5tLEM0Z84MZrqge7ytC
MjmHuFJrjzlmqf25YXYizlH/u71Tv1CAR3WXbeN4LI3yQ75+1h3Dz9LpJaEcHrR3
wF08ckpObu7EDm1GWtw4kH49h7CFVwEArhK0JW/cT8o4aB4Bi6OEf0n14oaPwLrJ
yYCJZezY9QbQIwQ0leTuWVCmXtpDCrA87Dha+XmS1sdDQgDCkxNfhmLwOdaNfwnA
6hnr5+DE5Z2khOkAfdVtNKZXvso5Hslc5uHUMIYwsmBJXKD9gCiWnl2AAm9v0ycX
D5vMSXnfhLgFG3IQ2HmbxapjEpxa87+pf6CSLGG9byVNuHTttRM9fjJrTLVC4hUO
3gHF5mDeBSVb4J8K5/5/aV1BcILQgYzfkUQjyBX2sYxS7vC8/tleQPqqR3HbGLQ5
0SKkZKF/zGPhkaro+BEizh0o29xIaJ/fnzbdugfK25s0GDyVcBGxUs4rLDLSlJoG
+RsNVIMH4k4cNCou0+HW+LSn8FQS3gXIfDybUgRpBJYGnVB5PUtC/dbHcZs/526I
S0EmrP9qeH1TmW/ivuaCKNyYRh7PWFPIJccsZeE+P1dGmRYjTMspwT6rbOryAPSz
KNTsDkE4qxtsEkjvF32qdk6J9UTJrqdiBHI1dpC2Xe4KqDUNLHp8Ze+iUwGjLSWB
nsmH3hOtSb7atORlSF0H+AHs5y1rOqx0H3n6V0Hk9QdHELhuJBDbEAVDHhCe1zG7
xcnpIFOexPIJY/N/L2ujNxIdzNtvWLyCZ1Uxg1ksfC7C5RqyGLIv6I0CNg8SMlsx
b+hsOb/mAAuO13co21I6zKkAUI33GDo+MF5JPKWIcWeM2wl++zNJr0/nX1RfYAa4
0eizUosJbgvB3m28KkhNuo2q+d4A0XLr4Wq5tXOia2EYhM6469oz9t+syUYtQKJ6
MIKX/2hmt+XFuK2NwraidkQ0Qu9oRRHvLdblHGo5c+GopHpn+frZ2KNGhFXg8Rma
2kqzwzXaot4eZQtzZs230N6YQLWmdowBkp02cI3GKCd44RliUaDXVd6joH3S3mbP
RgXzE9v4yRxAjeoYvpqWATfmxuGZWD/NSGrISiciGWLhfTpAbagIH6tpdgHgoBFJ
8tC5Y3rTLo6EAhzSJYNkxnWINhe60bfe9RVnekskZa22q7gDJ7AqW3nedHhN8ldW
HAEkqCrYNDFxJGJC2/IJk0cJJTc49GMrbqO5i2WhP+yTeel1vz8nJIJnA32LrdJw
Cb6albGqbf9vhqxsQcq8zTRHHhWxAnYZcBQcNpYqhGMPcK+MPhQ/wxknyZpGbS7v
FmRHDpVEFf12TGPFn7YpzzzbfZty//64rmfDnQ+YNXu2iSptgak7qjs9esnyZCTd
keOF2+49WhbrMDcIhJtpCMCdzS8+sH2ZuUBT4GGQ4MyriaWyzBza9JdvrWgWFcRm
sJsMH2CDYNKgfF784FtlRNmxYevxqONeL9FFIT7p/URJCy8Dq1eS1mDDO2409fYp
HZqXm5LQKac7en46OVFy5GilikjcXxyg+/7ANdgBCBF1GXteRsGLdGJ3wfYF1yau
JWHoRRoxWhLMAQ0ndNrPYny6UAeKxaukzOSvCKcOuBtEQSKyVwJKb7lA9ycH9Fo4
ZxOGdPxMp7RNiCrxJTAcZRmjmxg/GXdeMYfR9kPbDCu572DIJq+A+uqz/BQElaxw
xoWlfi4hz/pvzO9ufwnrbJvSZ7cMf8H660vE+699AlAQTaEXzDCU4FyiOCYCBXFo
dFUaJLWujMg60pSGWCTB4m+6UEoCUkud9D4SdP1U6cuBN/unK9nvlnTWl/DuTmSP
9wTSYTZyaetS513U7UmG2dlXgxqhDsnnVRucZyxfhlv4M0lvHGjG6zny6ogeo1oq
uUTOiuv3lMxVzHjGtGkGg5EG6Ybw2h/quqPf3/GOwYdQHhruoQv1+H5wH17HJW8e
jsy3Tkmt4CODgs0d1GspE3+j/PNrl0iaufQ6AwuJ9C2WQuWCQrdbhSTSCEH7wnBM
eLIyZWB7Tb2+MgINIVsyJRorwQZI86SFVUxfGNkAhl3Qje8qhXcF/f9a6nZ0Es42
hyC7KKFWfUnRSezvJ4hvAerd8CuZ3ORsdR9r0UFLoLRXMAWabr4CNpDA5LDQ5jzB
MvpRK7DTY7ksb0npiBj74qDAIRTqQ/wNRYtKjYcAGHOpxNNBib932IIObnGzbRS4
oLuchhkZYvx/D25rCgrX9rC64hDxiWHlcElt+QjHqMVgT2W4izvDt1O0WYSKCP0K
BrQgjlMG5i3pMvab5Acqx/dnNOScogBRVce3C9zRLRmToUTHwHOurzqbcgnjj3v1
dxiMeJvxB0RSGNfHPunRk49R2Jpd4aLRzVEtVcrvCU5+1y+QTIdDB68F/VfjdIBW
Mbn078ZCPAYaUvhxpgtlByhf/ds3aHOFv3c2QO0kAl+q7TOltfDshXxXYdUQODB5
v4ar7ioqQFNueKKJ02WQJi7KD/GYp/FJJ5nb2G5KZb5atkZPwzG1I4mYzUbzKz18
4hRx39XQWIDCIUt8cKlQ9p+uWydPFMqWhGvUT/oCpb7WKzndWN7R9XMZ/vhDG7Ex
VoFrDHScvvUkMrpo3vigSvUAkmZuNCrR5LuN+oDZWzFSA85fnlaUey0GDp8exqSt
mOCSyy3VuS5yXFw1U8uQR2VZcPuaemastIRoIPU1SlZu0kzc0JmoKLae8C4o6tvH
fSOnJZQIH/NzE+s3g1LULsDsVxc1a5h9pkgZTBT9cuQGz8Gt/HRiKd6ots8FrSDv
D9/k1nFNeoGq7NMaXKsFk635VP68gloXkfDaFVu0PTwLUqaidgQVAvq0KklrHguC
NJ3cSoBl2QGuKebPWUEEr4nxMe82tpltDeXcOf/0glzTG9p2s/Z5iu1vMhbyWGTP
JxPUqkq+x7t0QlPCxjyVHTuTLVW1W3osABMakGSvH7qykQCYlN1GPq0IAvGI8u2X
vghe2DABLPnRpHaJ96brom0CcSNiGvsupV9IpC1inT5kVckiN38W4idOsRsOU99D
nm9Q9si9UjSJOmOXHxOhdd4LVmc6ngy+jsQ+31KCvOESYHT1s/9x28z9xs9uFcnY
9h5ZHeduN9h4/0Lp8A8cSbrzaVjchrp62zKLLqhh9/qlskPpOWINglFzQCpNi6kk
PBRmi8jtoSNa6Ox/Qn8jnIf80MqdUZ0RsyHO4Q3AgUwgoPSJQa/cWpzCern9Y4kc
PG9jgF92hcLi7CkN+bEjnmfThdKbjRwgOClbyMRBDGjtaI4Wl9PDi+h7St0MXmnh
vC/2v6UQSQZhpXozdDlHMdvY7WbYz26dj7NfTwFc42up/jJHfpA62hvVCgzcTXP2
qncTMJhweVVEKq0YsN2vGmwiRfxTsNWoSCbyp9TPecdwCOWD/P0WSrvugPEZjB0p
lMsqwQNQbb4kbxvpehPDJ2/shpejmjCZD0h974yrTOTiFdNJFyhbMyvfRKbrkAyU
2H8qmzC8ZpD7TKMTX1ocDYLIEMFGPfwE6T+gIfzMOYsoayK11Plk2w9J0j/IQa3b
75EI5SWodlN1vSthRGrDMU+RAqg2z1nyH0tvsME3ZtZ7YWY/cVo2saRh9rztwGRB
4oi3BQunFUJ+OaQSqMeX0VZoxTnYzUs/uXacF7w4dOhLDOR3yHN4Tz6UACa4uNEJ
4EjwhlIRdK3WMXozUqEdw+AUA+pg5gawUfi6pMETehWMCvCY22K+8VqkhWPVGXs9
F3KmDxHnA0U1Il49FVoRErCiTmaGq8rXD1bmZ5Xp36O9TBJ8IopFiUZ9EDHTrCUS
u/r7rWchyUS9rY0GI1C+2kO4NkD0MV+t8DXykEgvUXNthBf378106hLXvhjHiK3o
GaCl3FzDZbdgu+M17BqJWbTO6LNnQ7mqlSlW2USgkyYlFqHs/imIgQgPw2sZHfiE
JzaQitYGOyHZvV+OwYxfVAr/a8cwbfzyBI+r9m0V83BqkKqD/u2Y2LRMr7tETubT
JsIowqkHz2G2OVSkt898EuHG39iXjME9MbLg8yQaLdvVUE1i9cuYOowyqUJY+bof
zaSB6QnbeRzAnsz0ShWGiUlGGkdWyISwsf4pRkkRdh/TTE/be+tmco3Ls4flwoJX
vNHOnBqV+TfSYq0KMywd+/7MUcCepT5oiMuq29TFFV6FcYgKZIIlAmhuhmXD/Hau
Hg11ogfjo1QKruWNL7jpnmfZ6DRcJzSaqHE07UmadgtdL5RO2VTbloA4n6yn51+i
7wQfNVpasToC7l0JKImRwDNPP8YYLAyxT2EpN3PeP1sv0wzgaIeO+ITwkua70zZd
D35DZtUIkMlAhimi+fKwH9vvCKbbKkOFHuQStLqv2nnxBbOc7/jP2HDlV+IWKL9F
0giuhQozg05oOEZDsBnpxu/EalZg2jcygrZ7r2KF8z6m/R3A8lUE1CM+AWKia4QW
qnE5Z4mTS8NIkj4Ef+hxlXCrWl1Hyh3fW3oJ3xF6JO2D7oWdm50GdWi5k9ARkxa5
icjfhA8r+MsDA+/Z5FczYRGRsGdZqZUUmVyuy2z/Rf/TT5NErdqUlc2A1/mbIw9M
ggDkiK3/qoUBp4fFLR/tg/HZI/p6+6cw8g31osGPjKH4XqFRaCfQVmRTYByOI5sm
nkGWV4Hzts+nT/Po3hDTC9DiSoOtuGri0kQ6333zkVpDWH+pGlXJhSMwEFdEpv0K
7AuB4ZMOzEVfJo1lm1Fxg27foaXM2lXKbuhn6y2DgR4cUYU8F9JyAkshD0U8wRPV
xJKM6MGLGiYmPGEzWONWO0mcTqsk/c4SfZUwm0evPeZxkLtmwcUJXzrriIPN8qv7
VW1hW6Pq9BHeNfLq4nDZu9rCaNwpWNK/Bl3Ydzn9Asm6wQx0o7/m9i2Wg6DaMibW
bB/lFJFvaXTUW23xzhoM4syrKoIkLiEl2WY6vSi/QITol8IbCjAHQ5WGwz6Gj/xD
3zpXrwA2SfnpqtQpx6S0Fes4Re2zoGeqgi4+UWomch78WUTsjBFZesGc6XhFxJio
oPhTFzDkg2wygQoKfyGM62uvEZUP78DxMtBl6e9iHZVr+msXMnR8H1b1ZaoxGd/M
9W8IOPKds44sHW7n8nIQi73GaxX63snmCTakMAO4ADHBb/L8qw5gfnpC4QseCFst
Qd+WrpA77I8Jb6sDuR3/HfvxJ8gPpOWrwJ1SKeD5VpcB6BFk0npu3QjCqvdbSAfU
nuaOq5IsexcE+wQ2cXoJIZ1nbbtl5VhnqJVtevcYxSf9ngNnAFkkNg++TTtoBQkk
zlz1NV6VVlbhzJEf9IfBhz7DiwpJUH9KTlZWxghOWavNPWlJzkLnu+CdzO5GQanf
An2cpsJxvGXg17bU62TBlY9EYwE1SbiwH+g48mn4h6JnVGWc0UzPPXV2ZElsWK5V
O3EA33p4KTqbUMqiYgjI5LApF4z8tCFRp7G99A7Ldt1QSikjfer/RyjdE7Yd5qou
6Rh0IMooTBChvmoTBYaAh/2p3wW9GTKbZeMjOho6PD41ziI9QTVxXN8CXuGeVm02
KK+G1gKdToxLI9FSqKcFemsIeU6yfvN9VuedKK66iSoozs317dlC5NW+6FekrG1d
MQ6TRaQKEwrTTFWCd0XmxnpEohm8/7vvebwfwP/G24JMS8/a4Tykmn41XDVf7g6N
v/v00riP2lR22QDg5Gr9GC6YuVzMyVcLyeCYO2dGhywwmCEXx7ITlmJlx67VFhgG
QHnVm2Phcls9Bpue4VettsvLxiZ1qBMG9eGS9weRkAIVgxw8Wr/jN1JAf82rxOUY
en1S/nue97TmYXZn4EMXDyo7AtabjshaMMJKRYrF8wdegraKLar8xIfm0pQ6MgZ4
3oDuWJaUE6mB8MqbB0JAYPeb5MsEwBc6cP4kx4x+MIzqTUR8/7figATJEuFnYIJc
HFxKh1jN3i9Eo/dhTD+zA09NH73MKGgrVgOxAed9RLejNTx7bukRtpDj0feEX/1/
GQMblFeRKm43iw/P/ECIG6p2IiuUsYo8sH78erE9AFxj36Mg1fgdoZ0B9g/G9+U3
96T62MsV1FUP5Q4xwIpWvSfMpPouE0lxqKrlaAoChkTSff+whhiRVG9Hu4IzAbas
710pRQ0roJOgsJyHOOYQhHXDlUbZQjr6lHrUmGMfzyHhDuQdlO5gvdp/j3Gspsgr
D9/Zul2HU45b5oIuRnUGHdUf/Ko/A17Ash9hkTucURb3KqXA1JIn9oZRyjPifjQ+
lNwDMRPaV4ZXNjV0SBb/wRYOKrE474nVbrqa03Ij+1Qtsk0UWtb3ZUwBtKThjaoe
UhhhQoB7zrNtJjoCjaeINz8QoB+bmuTxQtlNDdCwZLXfSpVxsgFC52tS/OLyfcu9
Li+79HXCcuAj3ND5P+/1rL9ouJXBCKMHXMNhv1fg4ZsLU0ilW7RTKNNhmQZbNpfl
h4dBQ8060JJDsEpPlIH9EArlFuPTtXLD3OrxS5ufZlOrS9O0aNLord7eFuLSjxGK
Bf/4Vtl3zGJrNfj9ekcUL3BNwFxvDSe0qYb7V+6Iuc7zte3K2n8z0QA4/G+Iu1Gw
yrDc2ERk9NsDXSd0E3T5XSBPABCVhM3AO1Az5u9Jw5q+FHxOT4Z9LibvPEmBULkl
kbSZJMARjclstRPJ0/VMnlyjgiJ26S7R5JQn9wJuAC3aLMBs6RXxNS52LThCqOSV
9bnHwBvUs7qwXtpUY/RFHD0p9UCwc8hA6EFghdvY/+OlJWHteZPPcKottuVxZYaK
wUAbYF5JbiJsAl/V2sddeZrSMqKYlmdky6x0eAVnCZjzuWHkVtZztDOUbdz/w4Zl
VSn8vdWOqsm/RF+AzXv1VVaPMQWxSbLTlOJuywoHjY3z8FZTAygFX93vk9yDrmnO
a+wzXzXblLElvs8Ukmxq763oecgoVt5onAS0WWdn3r/0hDaOz1e4FuNJlZZvtW1T
loqG4zJvqpCM0ue6H+KoGYM1uYojdSq31GXFUcaklds7sszEcs0Fr5Nj3rKMUv0l
Jp2AMSuxmBl+CU9l6Skmn8sFvJoKQYvDXq0eOHATVXlo8nqZvvY29QNaCbseF9FH
CoMrZZgiUwkreGOFl1BLAF4Kf02rg6njXYQ4G1y0nww/c2hOoN/lmQhjI96WmajF
vlzMg54a5h50Ka32uIHjFK5KPVndefkyNnezQ8nS9wNgGBflXfqv7b0yfyLNizaE
x5L2PRVX85Y+dg2R0GDnFUxmUQXomhpuA3pBvkz2481m689FahrMG+HRYfOCzSuD
A7iJwZq9BREyrzJBktEOcN00hkjIhR0rUCI769rcBlXb6/8cxWoKOOtokhOIwD0d
/WoMw9cNTClPu4bgSp4/IaoTiPhiuXZqVvv4xhEPYsBNoGiAQvbWbem5/ag24iYO
AvaTQDeQkQXaqZvhIh9Uy4DsGee8g/yvWtnt0NhpzfBvE3WE0HNpCHNQacL90uXY
EDn7A1V/w32kxe3vLjg0PVdSOIA2rbZy3hR4ittYeV1gfdNmInLS4hPx2DxsRZg/
FXllOsevwUEHncDM0IHHyjrOQjlSnspeyn3isOAJdjY3cs42J9ZDcphhCx/Jlgcs
S7Cvj6+IWN4IPGUvPZFWRD5mdM88V1p2GoYcfHyYF1/5l76YwtAhro0KhExwLxY+
Hov8W/yNauqv5ypx/pY0sIfGBdvhJ63sZCCrfYBrOr5wFVsToq7Ldq2kvhlLRvkn
ZS3gpCSGVdhR+FhZ/zYiBUxemaYvaoAr7jLYPqrH/xh9qm+1CRrL76L+UsaISabV
g7slkyDskjgk/TBkXFcMBNM2Yt1oOqzCjRn6/i7HcJe+V7WvRbMYej4dLWNmCpDh
m91puiQerzf2SyzLDs0bOa3bRKagFIzEIEEsvItofYw+zXl/xDMsHGLD6qmG17xM
YrPJpUT7/yz44dpgZMQsMCkqy47E7hbpSbBPDMZ23LbRoSBS2fxj32DJRNFlfl0a
LI4T/qpPHrGZE67sUzAGPLtlm7SP03iHsltVDXjHoR/joIw6k4DWIihMpRQBV8jH
BWAG2rW+7CUg+6hm3aoyjihJehblmPMAciOUTMew1SJaLO8glUxkIXPVSTyLfJf8
0JGUUYqei6o5iMXl/mDvSRj0+N9NY8hH1Vr5SUdAnJHXY/HwnBebXygjfmxA4Rei
WoF+rSFW4r+J/vOMv7zbVLJ6w2lnQTNG3+BSB5d7BwAO1GsQgLDndRJIGZKuyvQI
uvvAKrgwoY3xZGZWPf7CdlbbzLKcwXAiMLS0DlCxZQjubviuh8hTOuCjGv1LUjbB
z4rqvew4o5mBYvtxaJsHjevVzeVr/bDxYfpl/Ro+YPyC+LllsSLHLoyczlNmkB7f
IRCRTawNqQhKpNxTBX3cF4ejwJX6raY0ayK5JhuHL/Z8hv1tXlpx/T2ejCI0s/Uj
Jlzlx+aFtMKXhFluic+Dkywel2JTMQ7RFSMxaFflZNV97G/Ozy1JNGw89oPH5iU6
YlmgqsJ73JY5IjvgGd+ewOo7GvFF5dwcHWyGKs0/tNCXVFryAFFHX0h2il+Tj3y+
/6d0GfDE8uHG37KtwH2t6vhSES/zhuwgnwppC32FaKp+V0vlJlgOXDowDDREZjIR
UA9qhdG3Up963tkjRF6Hqza9TZbkfhoS0ODguIeHCEs3ruomghv6uvi746ib+3Dk
xXMWF9gnq7J1IIe53az+rYEgBXd+PLSssHMUxyfoDxOSJdUMWX4VPTpVFzc187Xu
umF5jmT/VdH5m37/rqt9lAXNS+iA006bJffccGkiZBJ6WkO+6tla1xrasyWpAnN0
x7bfNNNXiYeiKDywaaltfvdEHFdb+BO1NM20HZYomS+lnDhi/S92syFuQhTn2P29
WuXAD93AUR8fMkt6P9CWWtmgGJ8bxo4oHnNIAMNac+I7vwjSlx99vT5OW5rZ53Ah
JhnN1OojA+65BfBjUvop0kVWNBVMWgeoOSi06t/sog8H5untaSNMSARyJChBQT6W
jBgqy7g/3aFqtqhqyCehRR7HJ+DxyKFI5nR94gjthiLpepXBBeNHEwzlI3RwXrPD
BAszM8EeG81uLdenRODYHweULs/bqkQ3onOCawbmXrEXSSK+bKdJkBCjtkMk2LLO
VfW8B4pgxAS7vHOaOTfQSON0xRFwG270nVX2a1JgsoJlT6CZcf94uRBayzWK6IBy
LSry8sfcLWLYzyljjONZhNUDu0mwOXjxWE34CPryLDkQUMA8sD+nGoSt6LMXAuDr
fjjWf/dfj/BlltKIlAhCieDAvMj9FLUqzh7txNFqsfF3CdJMTZcA7f2xGNbyFi8B
TmMsGWkrA0ef6M1/AlUrUvlIusgOD5MOTLfiDn9N+gRNJqgw7kWnrEwrvCpwwdyd
D40Q6sk5TEpkkYU8VXOTvD3KQeeq4GjuBkuIvKjNl4olMGJ61zuR5roQ7Sv/Q0Pc
9lOLa5wHXkohRAgXnZSTVa8ky+cHaTaAyPI9EwlaWT/LzIphd/YaGYJxQCcKZmzk
EfzTvClbEnWYW0vAaT/kviy7THOsFQ8Utp4mcnLuCf/2dxbNlI3VK2vnq9XD1vDP
eCMRthL6u0EuwAmLRq43ky8O82yBMl7qcjACJx0z3s4eIaaxpPx3InlgU15GbRZe
GjCnnzKMB15ZeeSVXOtx5VGEGSDPceaMnFYV/x6vJy8l6rltvehtusZUZI26Shwe
wX6JQUVYR4cgiBH4rEZfJZuDRK0vRvJzr7q9qI+caLdjzKPzys4OF8RaYbFO1oQ1
eKOUXjhOS8MR1bcgkaYKkNEJRX/tTSsvDPR7o9cz6ng+Q4uXlogkfxA0n/NmiN+0
xyKflbbWI/Aik552Pp9OqrHxRTVqtKkEV7GUoV95n6Uqqw1EO/qrJY46ZCjsQjxq
rlTEnTxobnP5YuXZ4uATcz6whysHemqc34YZ2wYNFL7opCXF1yjuR2ZESpZ9WuAa
ue9iAET6rfkehqtmOhO8wUSggH5CPCBrgI8tZ//rNkZmmRIO9ZM9NHgwhTu6vjae
wQJOlA7SCotbv1zDglxRQwTav2oVTyLyX0qpXBdlXkTez7HG71qFEdN6e29IbuaT
i18Ku7mE5MnlAWyunur2vjffgVc5cWLGHGukFq7lAzGx/F2juBfI9UX0mKWJUJvN
T+HR9yAP+zqyH39j0GTf+mvm3CeglQBllLza5+fGFxAwuw4qLPLO54wnmY43xlMg
CintDl/wjWYt+OgS7QnUlkkFHvUJ4hXATRd405Hbq8+MLRyAMui9vRJFNxjtmZxN
1akUw1Jfk+CFKm164+aM1C/vNISnYsgcGRXNpt/KCoHRU+rq6YbX6wc9xPiDK9zj
pxIYJoeNmGNKwhUtI/xd2meFlSyj9NiUALIFNTjd9i11e0bdsMPeKLpNOr3l4X6w
WfWlDdS/MHvpcnH4Q7ilsc+2/PIVW6nv3P/tSfy4gD941txJkcuLcIyuoMLu8WFm
pv7DUkmG+hn5N4s67FGM6RfWwUabBhT1P+CXiwfzaWUvFPDKF8GT4w9I+i7ksIkI
BQXFK+mCLSkblAVtUXjP4fbawO/VwFIxPD/txayhBNzyytpCopCXX8WhfcHjcRH5
wJAZCZJ0OTdogro+rXJofzlD8Wr+gdb+qh1ceHKP7W9oR2N+qeWvXd0+WIAACpkw
HXzq3+xqDFIRy/5ujmiaRtu5B5DFgbouqAUP1VsUzBbYB+JFvC8Q81hgl2G7+9kf
vbzdgx7Ss6bDXbo35HnjZXxwYdcmYIfG7uSTi/JIIbb6FIzhHofGMKt0Z3E9pXNQ
o1mpDJ54XvL1WYiH6rfaio5XuYIdY5h5rGiqfgWXV9b6DXpJrcfPQ3gvycI1TBPJ
uo8+6B3+9pcQpP/7JuGrkJzElluo76qSqJjpB7aJnFv4ToL+Mhf7x2VsdkDUr1ho
CVV8mI59ULN7XiSxazIJr1CAe7iADKD0s8CHobwy+/BnNpRawYLkAbjlzaWADRtM
CRpJIOR5qVTdrQRfsO5sU6gNLTSmlPNC/krGTCFxg8nQjtFUYFr865mV0Uu1QvjW
maNhEkq8EtZ4zumRuLh2/twsezK2UE4Lhf6HtqOcBL8cF11rrqqOS65tv4FGIyZM
fSlK9XUZvSsAYvBql1QaTGJ58ojOjrqc1Yoqc5qYO7pFw7GFUKYTNPi1zsYVYD6Y
tLyRTX2pdD7m912K8Ik9sn4jaRstsXsS9Edquhxc73rATWb/C9JQWIF273PjJvg8
fc2cewp3w785WpZFLOwBAN39Q1azsd8gGDMKLDOR9QbsyatdKc/D9aaNjewv6FRB
MboWgvcIzJTvkp0qfEOc+nu6EuuJFcRkeZS5YY+KGU5fn8+lSQ8gK03Z02c2Ts0I
eIolVcrwfXttHdk3sbKaCNvzQdfBkvYfjmROFvvsw3sanFD4Lt2dgd0RbbIy+AQv
o6xWq+s5tciOWf244Ly23Umh2dtRcH83VW94vzygXMPTlsZCkUz4vMW2cR5v97xW
WFkKc4IcVNGpwTcJdvKa4XNZk5AbaEUiF2rckPDLMSpMzxeTdfo4W6GS9DluIJXg
AXZy/RF6CPNHPbu84QodmQ3rkhvKCNrWSRVRZCL+lg3jY3081fhG4HI3Q+d3oIBY
aOYQqmBXRixQAcjLPv64idF+qM7FrdQGp9EqSXXBNAO0An2ZYPxKbDXWOspCmpSK
ye7ENnFX8aLaWbtdHnpYvcVJ05VE9LVnNsHV2HwTEXbozE4x0DWZGkusDJEvIhbv
/649H1r9ZND4yMNAMmA93zMUt34Gcaev0y4FNoxqY+cRyWRaP9lrWv25bp1Vvg+p
51DhSG2J7mlOhGd0e/o6VtzHwUfx097o0ebcWovTDRoWeYbeh3iXGscmuL8e9Twj
rz1Mv97q5wn0Cp71vbZr5F9DvEqHf2r4JOk9/4AEP8iDf6nb2CZA6wfEOdJOtkcJ
db+3W0fED3luNhdZKhdR6RZetMsSfv6wYpcUzFP4taDAsKRNTvJtOlPiQUSKSdzP
UvkL/EiIO4EE+chWBJKk65zdn6JlViTo0AQpfGerV91kLkrrinygKFyv2/6iOs9t
GO+lFT7RKlCa4qLJ2CMw0TkH+mxfV9P3XAdQVRRx6mp9kc0K9GhhQ1SXsrMiRWS1
SzX7s2i+kDi2HZKpnQtLxPHa8x0XqvOxU9b0e8YrFgFgNGKXwDMcZ3D3qbjdcrEQ
q90+e+FF0at/25P1KmdXxdVEMsQOgCZjCdovWEsEOmLOElvc0tmR+L+R9XmfNKzv
NF7l9/7HIPEGjRc2tfFulCZCYjgiiEmZ1YcKD3Uakh4b8BVNDwrzwI8ZajtWq5p4
Id9hBCG326u5gKsYs0vNZcwp/EeYkqz+7ecRZbfo0xK9kHaMPwxuDi/XHvZHUQrv
jeM+EwK+DeqI9r6ymlku+JSVqLxO9cbiWr0SWRB46HA+tsay/1CJYybeFvETZ7s1
i279j/6QtGzJlcmlPJrPiNYeOAyLgFazmKZdIMOckOUWiceAlnd5dkTFnBRn31De
C1PaysNDaEy6O3g0kHGBvTIfM0lNU8wABVbL4rBMi9sFEewlD246iPJ3qzTJmiH6
awyeeLltnsG4YRFQrG8ZORpGErwIcUCLw+6la2OaGx1nMMfjwBWZMf1lW2QKC08O
4wmX6ht9JtFMvwP3rBnxp4oEYmkkLkeu+2Sl8J/8lZVqq1NiY0Ai+Sj69q/33UEV
d0zygs17yf92VlhSahlhmnjSKQ3bhkwJcNs0KXs0VoiR8RbBSN7qAGjZCW+eZAQl
kXE/Y2jXc+YLSvPgKUhw7puzRiJnrZ6TChkr3MMdLJP78MJHTNAqn31nkbPR69LP
DmWuzLqtkP3Cwibmb6fhaLRg8V1tdacdgfJWn8uym+z/AiVVYtwmgq7/wSi8e/GD
t7UXvw3zpXAPd9Eq+eMEn+DvDVEBzeITm1MMz//X0BiWJhsi4j5yU4yZUo23KwbN
lXgNo2LU23EBsk0uHqe6c8SKsteJuv8S9nj8fY/SMWKunvUOn4S1cVeiNXLlvzC/
mObxIiZx5kGKXdIC3jQuQ8gcWf/QnWCjRv4eyaJzW/p7nFqqQjzi5vE9CHmVjBru
PVXrcPsYGNsybJ3AfM48Y60I8WZF/pVutOgaEj4aegcB0ffhKr2TzqkZrI91CPn8
KZKjDsbCt245Zp/OYVXFlXhsxRkWRleOnzSBUpIa5eRKAKiVxiTWmeQ4H9tttAvS
yj1kJ4z3Y4xXw8Nljsfs+lNkvPaR/Vus7BTXu85ByW6871gEPooaXPVMDiibfD2x
QkMZoSBpKXSzGpgwsw3g16j8m3X56q6QfgD5CxZYKkio5prFwSRUrCaOe8Bnn92Q
DYwfhvJ+NzDIF8xcddhNiQ77X3QwJMUN8i5GZGCaOrfkly2lwCOm2C66F5/TtYSr
ge3gLvdTGZUfLRgOa1OOe5Hcm2i8efQG9uTWDLQq83ZDR+Wx96wkWLAw4eSkQkOB
6j+SNz1TUTjgtOn2iW3idlU3bHyUjsGdYF8Zh7eRrynnywVeZI9ffXD98nqaTXGV
0XvjO3NWAZiwMReb5bS38H3SNdynceqnPRDFIzm3eClwRrMuRQLCsglMW9xq1RUL
jUOlRNKbW9bTqT+JejMg57TXu6iFQCNGsSuoMe3D+RGHRdJl4VUHi6DfYL2hssFH
7+gnHpF442mGtcBYD0Csi1xHt31wcrlwtrhF1CcblA25rYOQEclF5tQJvbDgG87R
VygQWDnQ+kNmD0rBbHDzLCH7Ceb5soX4VKcdHjNtLhcI1uvC9nTkDlhxFLOlLGDh
TyMsl3zDoWST1a+j5XHOY2qPEjLsesMr7pM0fYtklaPguea/W+VEQg4xbwbvgjCV
Y9C8WruSOYOz0j87AQuONm5qZpzscYQnVhFgXfcUctHvdIfsrp/ijoh5RtymYqqS
iqOELmUYMXsq1P1WybuT08dCyBoLo7lNtwGqOTDtT0rdZYb3AOIh/QEmNq9/LEHQ
T10XyAaDaar4NK0ekKkXx2gaky6x9oES8+ljBzig/Sbzqy4zYNrOzu8Yy7jMmQzL
t3updAznJhl6ujs+icB/PW2P98Weu8njfLVcs1xoFYthfqZvCyBTRs3/PDowe32A
cbNjZAoPjKhhnS1MckOTuEUER3vZ7cI9wxnANyaxSTNlb798CRAeYR9BGyd7Hvrl
44/aXYLjeYLgFgRT0yMnOVRPZ3stj/UQizJHTSzKtwVJmiN5r/f9R0E6AO2J5o/E
q7VdkCBtYvRuljocX6Xwv06C/AQ2dK8jhGCsLRQv8mIAGlFbQUtM0UzZ2C+jG8Wo
fRq3DV4Hy+1OrlQiryfxbHI3jSWdbq0m3pY8S4NYclgyRHVzN5BUY61Bw3tBbspF
U+75UlKW8acbW3E7FZy1L7NmF7zWDHCcVRvvHYdKqc+RymnwmZTqvpQAh3THKNr3
mmTBOFbyK9PreubwelmCwUccHU8llsGTgG/S8uGhCiSyG43DxA2Mpfg8NOVyhE4n
Fw1MqbdhlssMerq96LnW5x5eW+jo427ZFbYM56X1HHj13G/ZeSjwpPB8IL64aT//
/d15CpMd2aNVZUFCQA1NSNJJ8bMPzQx+t4Rmpuj17t46wvSdgJfWAw+utWFcAm0n
HNA0P5kArd2xvfmKZkJzbjHLTM7qeoeprAtCjUgNTatsty7N7NGSL2GKdjbJ/CLA
leEZfyb+vedbn0UMYW6H3qAN4hKjomrdsgw9UAkbIqraTSnpM/lbW+CZ1vm5iDkd
nDhhUluAxM+2epUPOmuP2ZVCOfygDJsAPgPUkF44UCRgGfqvpzl+Ob/XRIOTPYlj
dgYsvDb6RrWZ0Ld0fwhBq4C6E8nhQSYLs24X/aRimccPxiMW5HJZUQ4EspmXbAWC
05ZXH6JFtCIxhPy4WWDNLW8C/Ri44s6HMgEVrjpSt80mweRo+lyjAmxNtnJVknj2
/QX12gY+5QgFtaTBK1TL1uyAfQCQeUxDCwrUU/CpRt1BKhJaPIut6EOhRiD/rv99
gv+lkJ7JtwelZLxTtxb3BIDg7EBnUEKDctWGeb5R8K62+/TYia2CMBHTO0+5LBDp
gZiKbT8DikwAKrQfUKDuppJkk8gr+iUvg8R6bXcQ2pPLNBuuzauSbeDDWxzHjDVW
fz2JS3/5tRG86FOq30a/QNlkOUEsPo1RcB5szLukqLDLTELC1QLqiO2uGeEaTPFw
/NUGfd1Ye0qMMKEjld6QACk4lBifnwY169uU/elX8wwIy/2eGz2UA7BHb07hTeBR
wqv+Y3iyusvCVT0Mt90dMMeW8zziS2oFcQsjf1CN85Ck1Md1zJRzyjvQwZsnzm2l
5/mlm3XmsYQ5fpKjQ3iArJTIQnqhjAEqEkiplIzkubbcBBJByQ43VCPOZqjjQENH
vvvRSnO5YyVB5aJ5uLiT4QPbu/30AEw4TmSpaofEK+njwIL9dS6kkl+OCPsgDjcc
vv4Mb4k/eVRo7mQujUY5cI63/gYNEaYTm2ocYIAjEMIVxtfX8mLWEXtZrUpDQlSs
K4tRzCKIEMuNIvbORtQKQ9E/iRVD61SJHgN1Xc9pmpvynXyqJaeDXgOmKVtBlBM1
C3s4A4M2WlzMJo4Ar6++pv3SCaUvsT6D/iT70MpNd8v8UZF+ai4XwSeQV++lZRyt
QxydUFUTeCdKpkSWBt/UFrR/Vf5DNTzYlXmb771yCjG7uXqhVlJrkeW1X/YIxiTf
3+dfs8G6xeRTbmt5YR580g2cUFDFQxR+UfqONlg0AjZLWYwX5JlrVvbJjyjynO7+
FCD4Re1lR9jg2h7IQFoOuIbBLhHQhAAT6DbO1GSr+bTXHIwGAXcqV7bh23aqGvYe
HKUdbLjs3uR5/pJDeFgf74t5YBNalcs6NhTVp/sKN0aeelcER6sztolCqz0RPQmJ
P9Ww8eMT1/eLsmQ2Xs2Q8CQtGgOfQAJNiKAC5px42IiOcEBsw9Vty9uDqZZoiN9V
tBmHG5heWYLg4faHWjkhegJ6sOApXUbnFOsxYnQwxQCi9GeS3SxWk2I6tN2Wz8FA
Ak53+4pd28yQ/kS79HoNlldIo7b81XplmqqD60HC+T/5uO/MVQQkJbq4lJUVuTHy
WnpQkIua5RAxJ1XTJFZbtFflqRaCfMKt/yrE5P2vJWMQfi9r/u5V8sWKmMpdNHIX
YCt4WSzZDO3QkQkbXc4N+FF5BT/6lzGQK9sadHYdIOLlcZTpgfCV04bQSln5PTqK
yM2qT7IMk5oPO1HG47jBb49IRwwoYVjwPPEZGOfkXr08HDhVsOUjE6VW69APWkyJ
4f/u78s3FO44AabrGyPBY2FuoVuyC5DgMkihpjITyN1eAJqN7pwLXM5okgtxzBfX
deYo6Kcaz5a2QoWDBskhpSfqdzfPNmkIhF50UrWhbKXGsTiIgorFmO4dFWwmUsWa
EOV1XU/tr21ecLoHQZhzm2N8K5hTid8ivSkeWNDiiLlHMEj3Cvugs2EeRfe2DSGq
SGKpx4g+rGJ+Tz/ywOzVE/mp7IWzgkVlnlQWNyWWFs71f9gg6u5Cjg56C+Hst5uK
ABhl6SZDGyV8nd/pvyD41whuQtUDxIFmgZnoOcQ2WT5FQp5o1PJw7l0xWp4N4tom
C9n38/2JHySKYio3JvjMb043ybWN94vSnzqLoYPMwsExb/zR60DuoqCbZijPvjqM
AKHxe8iu3wnBDGbsC0KjQr+2o2d6ixh8IiYGglHN+SgB7vzN77Y+YZc6oedb/kDs
zBOu6AA2/tFX2ctdkTl+RPCnpimBOc7eWJccu/RIqtfEIIPwSLxJUjpAhThwUiIT
Z3XN1uJ4QiNm3cBj8ZVeIgW325mm3BXm1WVc/z36lx2gwMrjsjMXdsg/xFJbRBaR
Smp5wZYknSosSrH4UZKVMc9oe8B2lbzVwSv2yMKrC+8AI6be+a15bnFEW9Fh4iNY
dWRoW0sAuRN+STleQZgFpKM6GAe1frsVyx2xxKrtTGMjYx2XUjRoY0WFBuZgROf0
aJE+Xe465ASHa18sW8RoUMbFUg47lG4/ltWIzVJ60MFuvTb/ypYaEFA8ZP8SrAwN
rNyNUWXF2zMqo3X+voCGktHeQMTPeLYNgJuyCsfFnei8mNq8ykRDjsllaCpGzlpC
yOnQoLMjdI22Yezi9ERK59YZm3VhkGuQQ/xLtHmZRNzkVWkArifiosbkQqevdm39
NI+VCIm3wiiN1pMLVv+R9Z3qCD5YQwyBWNpqe4VMmXAyde7kbywpKCkTR4iOt3ig
C+hcj5rzhRx1+bNL5T/BvHWkMUuG5AE36nEOm5r93/k2UT5WdWVo+Dhu2n0lxDsd
ZlC2xEZiyop3tY4LM44opAyV53oeH1P2i6g9+sr9QWUzct4lwNbgA8JtvrDnHXRU
DN7C8798NzPaXZLEuQt9cHR5IA2TSUooJemgnXHpvJcxkRQPwn+Fp5HFaYJhPZIW
6cpQ2YzBP3JpStf3fGaUlQ6wTzOnW2jupbdiDHfMu/59JA0aPU9x3tMYVM7vMEFq
QTnu8ntD+ps9FZNmloezCd6XmhezXF4zeyAiHlsNpT6RnpFINEIXg4YRBVkY1nTl
3w9X1we8J0NXvFrk+ZGGDFdn5S5DjPbsxGMebwN56Ho9itzGq/irDfOS4lc/GaU0
2CjBydiWnCjj/HI1Od5J3Ta5bYXSQBmW0AdPnTjSjk7RBiTQQ+SmtZDWGNVdth1v
rhT1US2Yr8xWl6GVlnzjrIbJdEibQNWvr2ePVSWJRhXQ0/tvSXc06j2/XD9uEMjg
A6UF0BAOqUHUNYjtknxWRDa1mscq3QgUGArMX5dB5jbsB+8BHy8z0vc/isT3IVyR
zApHOtCRuE3bTDXc2nsi/GPG9Aum3/jQGKcmhCYAdybee/Ag4f8ysflOsgm00P+Q
WdROx9H+JE4QM4BuP1f312irbMg2nym0mUO/9o0NJ6OhzSEDjc9yBkm5gK35F8zM
v1zumwUqQq6HWoJWbDKEy1Nd5W3lcXo6QtFf+RwUyoBTp0k01S5fX3aSsKIgYqlZ
I0CGHFyGa3XtwLb3+3K7rAs7WEsQEkwmJvMIX5cuuvy1ohD9LR/kfAfUEN+oREZo
qULZzPCI7VQt3y32G+gIh2/AohrdXXuFqwytOs0NXijJN49ubDwCa+gxdr8fEa4H
NII2cVGkiHWvnEZh+VHxh2dX5wutL+cHUOSaivMRG7CX0vuPhukITb/EzcuKHxe4
h24nuAJ+tJcijjyDyGfQE+zlhqFBalid9ZGtMXsXtiUNSTWtrpgIoLplK6u1Q9Pu
M4L9mYkBXcH49+56L8N7fGE7QnH7sDgk/k/+iS1VsVEX2QMZa2c1+R8qUrNJvFCi
n5QPFlhLHUM03dxkBCX2o98unnCEEysATW2hgWiVGp94oiFowGnXUhqWFu2IFdRs
/3TrUtC+gyWMa1H2qafnm5yjyDRiXGDe1vKIyB5pYmgagLpn8sX4T9QsZsoU9Qi8
y6ht8pim/83eUl0bQajdS6DhlTciDDwFxKns6DQMfVt6y6tYlK8wxbpDVCLhTRQc
26Ugz5BK4mtLD9NutTNptxVH7Z15o7eVlqJZBvWWI9J1DRpE9qbzU8wErnBo+sqU
jWuGdsPoMjxzLbSlBvBCnLJJcOUTVhorZyvfUwkUBq7O3U48HcXlFODf+n3iYUai
uvziVvA7iypbqwbEP+e7BINuXs7l5VUOQNizHPmvlkhoyWa8BAhuOdEH2jX/N6AS
MvXn+BdpCrB3nxrQBVLMFE+n/B/s1KjYDa5YO4WlL1Jl83VIo81ejyf8Gl3sjfKx
qZYaYBNAZkMUeLpIQegeQACuorY6qWgXtgHMupO56lSAspkj3x9gfYIrQJ+2fJnM
0nyRCOY8PlaI+lE8tW4rg2SfX5NQSIKKymnojuBRVa2q/ObDyK17GwUh7gGzKcQ+
q1I2YMyVMKUCVY0rRr1sEhDGo3HVkSkldncs5AKZ65Nvn7YoIcvbNyHGX9HaIblh
rXl2awlyGpqWg6G/6Fj0HNIe0+Z5+7t7TbBJLSN57OY3j/VK+mIdyojuYzrFpXWz
Ov0hRcAq3pLI+lva+dzcbBI8bkncf1j/xxA2gzaeRhJXI5paJkLaBR+gG9POvBwc
7Ka7BxdrRdn1Bwi3Rxe8195VbcsQJ1CjIPc+dVE2dBQDXW7k2sK2UmKM4wZzZvAF
qH+yAYsePcOxsrqWAPXhJcYRz05jakfdUVHQ22yQ0TrBN5K27jh+E3ZFISEfXULR
aAIYBFiPuwI1i54Cu0/0COMorJV6qCZf2XFeJPUhL2wBp1OEMHVheMqsSM7FYwIi
LHPEPi7aH+n/VnzEfDScBzynOoooIIxrsDMbkLoU1kfT3NGKqoI5NDKmhtj6jlnN
3A2JoMhPxcZGWlip8sIjKt+DuNwX3VZLYKMVtk2WSkJazDOIfJK6GeYK/P0Hlieq
ryME1cRKstLkbUpxWBTRLieTXjRoYxJZ4unX17xl2KBFAql40oSf5dQRFIV1IQ/6
4GCz+VnDBQWSQdd4IA8b7y85OrSG1os3a5czPfcREpzUwk9WKpMmEag/1h0r6EEo
pODzkrV0KJ057gt85l4VpnXybAswcKJL2g2QzDtgIfkMiJNpHTXfCXY8GdZp0iFl
fsvXVql1zc6XghEZLJldGVBvi6LHFS8OT0rlt7IWjxBeA1/JQsXLeOgW5ysoaZRw
zL3bt/2cS2ZMIi4iIJzOPxF1oz3tpeUB4vkGw3ddw5PwruS+W6U/btLYguVx0EJI
okYTRKbNB9HsDeuVrUUirnTm39VvnuJ7JGyVYFxXJEYbSqsMLYyaFpyCKO4LTdox
l/DOu9zQOw3NuEW9qvJyyB4n5V37uRLkxuWFYCz8iDWeftjqWE0qSRSTvf/SvN/X
63ynQm1ai9sIAQIX51+Pz4yjsmCq6CI9NM5/dp0hXN1v2OhXMimgzTAfN5ZnSg2N
NKD0RDxjB7sLmzqBvKIMgavoAwgkPuMllhQEcEgTKDrFd/RHUN4vh1FJUCrc+eyI
pgawnZdfiKqoroYzFDOzrWFXYaFYaCADVQWeu9FynHUUZB0DY4yv15Ld59FYWIk1
ggt8q3RXp2fh7AirQ6NoHPgWEZB10KR2y5+tBEooOm/fHiX1lEDjy9hmKyXHEOlo
m+FNAg/12t0GwCLuWapr9AhuFQ8JS8CS4pPMmsJrtOAJ2nET0s9Ckp7dPVpnspab
DO8g5HXddIAGAEAeeSMygxnU8mJvMCn2DlAbQa/kS+a6GQxzZef9//36hua3kodN
0k9B/H1rSl3imgZSGTCopZCNNuJmuCNlOrM7J5EZZ/CclHEHri/GX62cR61dMREo
6czqY7XR5FnPNlYtGo+0hXDhwTxJM8xjxygkuFG0ZP1DfPHryPokvVzJDlIuQnYV
jey0W0i01i27v2Im4JYbx7quAbi+vftQ3WrDvFEBCEfJcgWzdZ5PTagAIKchetWi
9zaoujYb0BSOgiqtlHdHjQrBbTp7dwvBjrV2zgQ/6UmpHUw5tJfdf3hn38yJxWnN
zVjnCeZUzSqxbvgemrMTKNAbhWEV2bj6P63g66GSBWQNqmG+Sl29qWyu1HoOUNTs
ev+l62hYMr74z7LOusQnsdEw6+bpwMDt/YQYjFJrBSumqJZ/lQZE8R5SeZPd/nc3
Wi+xJMKby0zh25MFD9qlWIJu5cfgMudLgQDJbYu3DW72bFAAhpNb1WGoPVPVqUQ7
+DaueLIVFhaKvwV4zGJoQpvzNPZH0Pt2aLkNaQ4n2IYDQohbs6UIcZCfHFmp9y57
df8wkMPNe0C8ZsAOyHEl8JVrhRFIQ6gLrxdHwBOSFOQS88Zbu2FcWGi3PTk9hD4b
69/OTOMw77WqL+8tjZVomcj40Ru3yS4V9pytVsCpO9242hx4mUDpH929ZkFqJsez
pXVdIQzqjoOZQerLWqQfZ5twdq0K6BfHPPBSIFFsDtlyo0QTgAH1UQv65WORXHGF
Bzp1s23C44jLqMOTMxCuTijuPLeSk1MSElDz4ARnQsqMj3jmDjDRhwaSDAwTpx/h
Eg4tVvhdCeInMMxFVx6plABPct9Cgt/dq9QJZS+QALIQ26t++PCWsiFDSkiVk8Su
91PROFyqGb6OTYxwLVLJ6AFvn7hNIwfPl6SobuRbhk3k3gwlWI/HlNAmFW2ik/Ci
1gajNCcp7PPVLHpRR+bMt3Rd/i86bbR1yl4CkJZVy9rmeGVDvRftnTy4FZ+gIBHi
cThHtyeRV+oSZMKoBUmokh7EY1DHsv2utEHTbnex984lbq6WNGwQbl26iSiw8kFU
YrkF37WeFqPQaAxQEurNzo3P7XnAsffnda5ZHVBCXbcQdhP3M88NaFFDVEEUEoj2
1DPl7ru3ju+YE+naUOQfFVwFNGEOmXd70pFnYSdqUE6mRsdgVAX/Zn7HlKgQghlK
QYp0zTXSzQVqi/Hx3RujSKots48alJJC+tA9xo92Dkx8myBMj9bRCQr45pv7rVmf
/s3L+pXgYG2CDaZ8liDeAQRbFd8rT5WVAhnveuwaIeL9ptZChU9bSXWFL0YGR6JJ
PSl3xT1Q+wGe2H2OnZzUjrCR3uhcXMaUJAnQufxFnCm5Bqbis95hGuTLqWnANn+l
9jnDvrNyhLQDrnMW21oXZBCA9dxdDVaN/IHe7efSvuf/01uefNdPbxT9dnl2HpVQ
pGUpEhq6ivR6A43XSUlVnVIeUnrKBSHoGKdtRXGJsZ5uHU7IR1vb2lPQXAyB6Vyy
BuMxSIQlgdCTi05d22t0PnfOBIKjg8HnHJ6/iG8azsgBEdJ1CRWln3SjfE+ovRta
VfS+uH6chrn576ktYIoERAzORsvwI5H4KP8jRFUBh0iXNUNrjqorJCTXrXSEUcKK
eEFhVi2oxCoLUk7+A4cVMis0H0tUD3wHrXiuk6NO4fWtz60jRjbGMlP4Igs0r3Lu
I9+LfMwiEGRA2L9AokAK+dDETxFAAML3wIPhUgD3PaREcljcRE+ZH6wzewVnirob
JQpCxlI6exAichf1/usGTQWeZoFkUt+zgYToAbVaFd2TL+szGs4WBBeAsXwPh341
vkiyx3HajE5uxPjSSEWROEGHsyy1sms8Hl81ndVGSQhjZeANSfdKFEMO6qNhXSm4
enHGI36hbTym1cT6MXGrAH2u9BXx8Do1AH7Gy7oRfpVyIaWPsUcZOAzkBODU2+87
WxkFlPxJib++2hq7YAqflDhsc8Sg4FuWk7f17mCYisCsz06YXeB/9jCPNw2Y40tI
gSJcpjFw+YTg8dYAmETEpwZBPZE6LxuON6FebX95O58a4QMGEG2XeI9e3IR8U1l6
WCHflnaS63V4BMtv0QJAXqUz1t+PTYPMALx4gdHF9Vv41tHJ9NoGBUOF/T7nIIBB
3Ge9ygKb23XG7VDdruUEkbPPvXhjJtTXNbB+YWtAIcTYjpGOAl8B9xsSBEhbUvQj
aopt9hyJkqY9N/YNQ2q/rUJPs7IpswkmP/5GOzIGEqU8krwidwj8wA4+MO6FK03g
SVNGhfkoZ05yLIGDPByr8YoMbd0P2V+WurECm4OPll3BPLJqyEpcDihawz1ae/GZ
lARYYVHLm7It8E2M9nJtiTXLmFDKl1XJgKS/bRfxAVJGqA4e0Qi//maA1tE6/OU+
1QbAB7dTa2wWWm7ZKN8CdHw4OqsxHquUPHpIBU/9Vbhx6Tjt+yripYWbUGMq4p0N
FpuwPkMBHLTyzF6953i2KYRbYe/bZR/cYLgx3zqBplRUtjCQs2TgatBq84Pxr/77
0q+A5tr9V6zq0s+e5fcdd20ch8COoxImdJMJ55MT0P5XnTqQra+DduDDGuiBcSiH
u0o3L45sAMIC9MV8lvbyXa4qy1Ag9BeGjzuz02gr92sIivz5u3Hu7LLgjIh+aGvX
PBrD6IJoXWu751BOob3BOGEkvUXZjDbKX+12/XRCMfMmDnCTvSj4sVvy/vBKwiD+
gq+1b/zs84/24hCDf508vFQvgZYVTQdvb1C2s5KEXv9N7eGICBmX5SVZUDhJ3/EF
E8aL3NEFA0/Z5QI6wvqfRiDAe/I8jEILYK8IQvkAyIXkMNSLjRpOE5XM+sdm5ffq
FkwYZOcgcicTuhRpG4tantyQG7lSbAOG55wcwV8stqGyyj0B3fF2q+erJTfNRtiT
CdfGVO9CZjiPitc7fJBNOkBKQTpYnyUr051T/xDFzCCja9SicYezUOprQizbE6oP
zNG/Akham7hoPNm/jWOHOJ56FfAYDuT0FbYim1nd1Ya4HInfGLI7zTkNRscBjJ0K
pQ4sxlmunef1e6yHS5YJBxfIRtp7i2zZLKcx/hiPlK+Ww5bgDho910tr0F0qOJqn
U8PahHSDzX8FjGrrUWAx12GnbrJP98N+Ht04ppXpIKSdPtCNQd8yixbzDNf16cND
3wXdr0WJ99X28hktqKfuFx2Yv0B0ScDl1niqXFfrnFAiLCG3VsKkwBkJNi/GnpSl
93G2dqw8OmO+ydqgD3UN95HVnqc/OIZLNtyaCp4O57ABZLkC8IWtwsHG0Leh1LxP
fKEPrFRCoVuJTKZPjG4c/eF4Q5oq5xp/f7jsET16mOLVVFmfUEqNit5tHjINK+sU
i/9fGTiwtww6EldW1+Gtsk5ZgLQWg58+4DA+VMl0Nfl2z1+OBWnhPsaLdQRMurFX
odU6dbW+lMhUq4bCQhECH7KOlXGyVdpHfIOQKyDNInimAVSte5n8phvOfoAtUZ5q
1IwwLVuSrXnUkgdzA8mN/d8Xp9/9jaSqr6e5yTGuF+drrbK+xSXv9jk1iCWChNb7
7j++Yg2HaP/+ojt+AeKEsa7DeCScxzR/ZObLUru2t5YCCepMqLn70sUoVAMWQe9R
fPF3O+XRSDVtC5NSPXPkh4j+5VvMKKLs/us82RIC3Yv62vo/8LimqJAOHcyeh/kG
SRKN0NXrdXt6AUv6By/UM3103DDXfmMmOcLlv+euuwKIqmJa/Lhen6lwsu0IjVFp
RZ2cJibcPZrr80hNGAsCQvDGZITk7eJXU/AvvdJi/U5hNEXYZnsUnp0Y1AS0K/bn
IfHI/0TWIdoP+UuqqvyqFjZBDJ+eM+RKuVReF3igxqtKFLbqjugBN6UaR3ttX9pi
TmltovkFsvJKaNvpndyRREl6l7AqoVeTtft30de27M024hqFSMyJrBZo6zo65KEz
tXDi6xUCLKERxc7ZMNabeMVGXaYGAi27Sjd9ur48RxGlFZSQO/mWd1uNFileBD+F
LRylDPJotuho4VfbWQ/iqDwfZpclKYstrAihqWoAgCOfPgz0gPW661rQwY84p4AO
zNFwDeIuo5Uoy49BAo6ER7182qIJgD6u8lbJHIirRguf6crwGLzca5cEoH2NZ/iW
rYuWe/dZBfIpGzgLNuXDIY+b9+z0RSaetHYrnKUpEsd6v1em/wLdNbtMntf+TWzc
WUnxwI2A+XKK0neBpYZS541ZK6DUFQ6LpnOdo9rPXJWff+5p1LpFV7GU/8/ni4Lt
5D9PGFPWfYHO7eITvJnJeKJwNM3UpsUUKBat4AJvE5rBCAfkZNYRmQrVV26S7N8J
HPb2nU73aNLAfuMu9fB6UXHVVLCtCmRPIXKFQx9WSCdl8diRNv0hBZmQVHIdb9Z4
b6NqYNddcDqRuh0tNP82Wc/4VSYpNHeKu0Q82ddsv6m4aqLywuhLE9K5YxzEfXK7
Crdirz+3HN3cSXmUP6bHKL0OMO07Z1nTkXz8T/Bi5mnd6eyD9kedq6yFjLFuIKzs
Ri3WHS+BmN3Ue2pI74SL/pyEfR8qcP05X721XEvbNNopNYro0o5yvZY0mM2tMuD/
pL70SwPQHKCgxVJkQ5cWFuXxaHqNnL79x6Xk9s7/fiHsO+yZpGmOhhGY++Dfl2py
po5grZjA/sfHPOVhACIPYk4SVNv+ZAxJjqcPdAnq0x0HciPxTe9PliefPrCgNy6W
RO71ptIsXlYwJoKQR0F8iUAQswM/ak17H5EnAqFmLMBSovSUtKRdjRqNRl2JnmM6
qBLU/1w2Koj8O+4wGlqr7PryIsLVXALfFXBekMajcBi15UDeLr54aOxTpcrtMWjL
gAkZOpoHkSz4mNmyX4S8gFeAnGIclhyVpR4Ba5H0rTOzQc6mMAD1J5KHwlhF57Qi
zmOw/14Fc0QLNMgxvGtUPIz0YibQztdLolGCUK3Bczqt9RKnUnEARETZn9SQI+cB
X3uWudW8PovqbveqmF16v4ewkRf2mHib+VTwa18PuKj/TSGnYkxEUefG3NktbvDL
8ERGiwNadcQTLe2GHbJqEfRTALERwz/HINgP+2P4U7k6AIT3rqyfPCTS94Qx0BQg
9w5K3+mZzWwI4WmxOO6EQ6suuE/HMoU+rssYJ3PmrAWpfx8zfFEMSpYZA0RSmkUX
uqkJ9+dO/QjddN2c2MxScTQr0FhRfxgBXzIOTrkBovfSiNHh6+zwOrOadd352p8e
cm44O2thf97dsTGmDRm1HS/jpe/zHn+rtDKqMyd18YBKS3Z/JzZk1Ya69CJLEIWq
L7fTw/fdOzcX0vd1vECA4qAfr7JC3POb/TdnRzlLBw4+6C4RqJ4EWqFTI4j898Bu
LLZfozKEDfZGBwrnp31yOy66DtvTEudE1PrXhQTzwLOTsW8cRTrhGEBFSy//xQ/3
AhROYJDmFP+Oij7rFga6yeOjo2hPsf4RodjBJBGIwtdE0SlD/3aI7HgURAKEsq93
3hQmFFiycZtk9cP+14xRNryxLcnh68tolKRgym7oSK2SfIZkGaVxcHGguMkC7y21
aOzqanI7vghKp01k4Du1R+j2/xdmcnCV7mEMVCPnl1HTIA3RfgNekiPxGMe/TxXg
qz9GP6GfAcVbKjTu6ZrxT+gSvBOZXlHbQk0QUsxmPFXsk6B9KExlxkG2j3mhTVDM
Up6T7V7PydbgWC0G/gGTMsKqu6GwbVc0J7KIMD+o+8J4Hkcxy3+ifiWaEF4h2ELA
LgECEmEwOdWaKLiCUVo8nFKleLJJCR9ZreXPHZG8pgGKv97oe9uL7/qOSP3u1rr5
jlogOtlHSHH+rb7gi4fgY2K8w/j02e0JNrotfm8FHIKUSh+deEBpt8FEg+7jx8Dq
cUQgscHQg0BPWCWcZsP3U1k4cGaJc0B89Yov2vuXa/4wzdqIlmTGdQZokeUGtWJe
qb6kfHIhYWgHrh70ECeUzoRuf4C+myQUkByPto7xSD+ePJn8LBibEzEdmk7f8gS0
b6pK7OBhLcgn20Ncn9J3GJXurXYDxJUd9QX3cv3QH2XeP9JEb82CAXzT3hDsFLKe
9Hvy3+mbtRTd2t7rUSRcT8LCXXp0p80T1qfHMQlNzuMytpbAfmI1DZ8d1dJpIand
rtotqGyYn4fZHHuG2oLbQ9bNmDp0dGdcT1pKiLiXhsadjheUhVjbI5nNuYyiuJJ5
15msHIv1MNZVkaYpFPmyDdfPcfz6oWfrt1ZUJNVpJJEXPZeXNOXWVBY8qxFKBSBB
RYjLMnKEBs8s05QfnDocPpIG1AS1T8W1zbuesmshTOVYsdVVzqYUbGB+wYBTqhn0
5p2yJ7l361se4sXYfmoq/m0JO9wSXZKjTIhvMKdft4h+m4TuxlRCqg7rzxBiE2+z
aStSU2eCKGE858DY42gIY+CF5I57wLlWhJg1FcrX0j+5Ih8djMxDNQb0y+BTvtII
S+Twb9QqQki/v+djrJ5uTsK+7U//kwKdS4CYD7b8RxW0Sdb6JBdxN59jjyWt5oqN
MyCSCGbIpRcEXNTr4ArJBWdCYwAWeHudZavKaFfPgeoRCXq1WkZLheoO8lAqoBjJ
gahLlRCDRLFCSVWRUaT3BwByFxkEXIEqt74jbuTZ8fe2zhRZwkyYxwGiMYyEV3Hy
RLleQ/5wxDi9WWKoXXDAAFGkO6+S9WwC/Kuh+9vY4CL+095h3sTEXqybdAC1A6Hb
ESLSNpsqVLiwLdUKfx1xzyqe3gfLF3So/N7wvh4Z7TwFlkQXTxpHgQtXkYq2QqGE
SHHXQsrmN0hvu+0y9M5TiRQ2e5JUW9octyWEYLklNqt/aH/rppY251l3rz1H03Js
vMkaXaaMBpznYnskhaH7iun5RFbu13+j01IwwiGzxRtd/EF/Tqd5x+swVYNUieNG
lnETW+dyQgg3fOgz8XFyCQasY6XOFtoOVcef/392a7hD5GsQdfXhEkmX/jdTknOa
Yoj/75VSdM39KSqrX+WtiwWoxtHCXzjkz716GbX769S/1tBJnNxaddPccpom4JaZ
bqRDEnQnOtqaV3lIR45gylVDLKYdWkV4Yo8mItlhCA0myVpN5G1TRHurj1A7hVf3
fV1s8RvM5dZRHb/B7ytq1zsddLf6oHgebEuS0iWZJGVExuIogkBt2JS21F4MpHQe
+apLLhJuM2ADzLGoz/Iq6uI895LxKh1scLsgmXa2jIudbcbWWofhVM0ag5CKd0t8
X02hSVIzRfTtE+dhQhrRdi4uW9lY92LgjhlwfAxpaWNuJU/TTKEpzT4FKCudaQWg
+z0FC8dnSFZFeAbGTCI1+c761DvKiXDUgVLuxJihnaIqRDr0FG9HPbanDQXxwZj2
MwbSwLTh7gDN8PF5ccPdM0Z0FX9YTLJgn1ALmAqajKWNdI/EePlOgigMWtMMg4hG
WxK9QKP9SM2BonjfK9IU+LKHjr6iKXET4j2SNVK5e5ZVKyOzEaBp2SVdb9rjLOdn
oWqgJDUxJOiMe+riIQo7a6eGDqW3kiSTOT8CSoyQx7FkBHznzjLdVK0dsdj1bmZg
HyKr76tGRtBBnS7WX/Nx3urNcKxW3c6H90deJYC220YHkUam7jqMfjtG+vgeaMkM
CRsDWHs6UEyyEr/DOXQG46eUQsoQKwYTBA852ZSDtf8ypkq5DcwrQTpAiXI+xAca
bZqqoaG34EU0kM/ocuTrpg4BuY+/ivYL2bmjiXysYIrHURCaSU8I+bpyDKeae7XN
HzeAxPvKyavb0cW0jG5S4EXOvhPcOVqFdOE2FOSih8ZjE0aI+0ep7bO9uOnuBlVC
9jViKqmT3jRKzP23ZoGpWX2bdK2QPAWJg1K+vjR0hFXglQH9/SPpU0KhVR3ljJaZ
pa1aEjOrVdPXCDlcHt/IpaMH57bD9GnJ1pSUewk+sD9zWVBTY/t2dKmfqLCAzkV5
Q0XTHFDkjlNZBEREqvGnvxPXmMfJcEe5tXw7OCIUVDPEIr+8iMRDDdMWgCzHdlea
n3i/9FflXDRMDIlv6xJ8rS9LGnP8ti1KuxxswNF/3zLhZYTy4OGMbQyq9TY+fKs4
UNp1Brcro8rh10g7firqZ+MpXUzscQ/Mer4ha5iZjhTbH70v+lagOVBUDdeJbDYh
b/vtITq5brRjpXfxCZEKQbn9B5SOyLSCLvNq1JwJil44YjTXboRP45uSKtsNTb78
hIIPAKVEpfOXdUcQkgXQ6xlOQaiMJQXMIlh91OOSc2w+HEd3/Ce4Fr3GzqctPTbe
wZ+Sc4NhVeTVpbuP3GiNNnBiM4lAVawViamXC0eQTMfWiXkVp8xMu2DjDD55KH8l
nCFzAsdwZtU/gnSePi5RCwsvYns2PQbae0nMS05sRdOyKJ0ueKC4xWvN7y4EaU3/
uoSLrTjvDq7cJsjM1LILtgXRq01XwoZgGDjfCegM+uTzuZHxbjwhyYmeoW50KK4k
yV4IZdqVuAWQs0TbsgIrr7W8LBFJcvfjiBkgns8kU7/wyOIUKIkDsNj6Bsim4jLO
w/PIf22WK0jIZtf4acp+HXWLsWdK8W8zvuPr2l/nFbYVf+zElwOZyt7AcXe5jVQA
B1VBu19MeMsFIIDsx0q06Ptn9UUQMlHwr869xSaihFQWqzJeaCSnO9gzdLBVLzMS
4QUyvdIX+dT/nLiAO56/fxvKD1GW2dnP+0Ke6Arxw1wDeb7O9v1KvS6MpOifI6oV
cT7g2yrd5HmVFjEcgAzUj6G26f3BjorwcYsFZqlTDAvQR8UAV5IqxXktYdQNM2c0
gs03oroKZ7+pXFc2Ry1eB0izzMO8thxe0Dk2PvU3DjcixJOS8PMUD36lpGO+QUKk
DPyaoBKahCmnBwTJ8ce4hfpToVN1ysPUo37d/vLWkh3eiM1kRFYsXmV10/0VkcjH
gbZXDRPsLjjvEwerzkgPDKqbQr3huiLTPbB6oiShR0o+/Ymypez0e9xM5tWcC8uT
InjbccvltxJI+b1VcIDFZyp3hlRVzJ3UIfVOkkZcQ96XNXuZBuNXn7ZPIS5m+kLS
ZFr7Kd5VNHRHS0DuB1mpT3dMHPGKwg6cfX7a/L14SRgufZoPrAT3CxrK2s9s6yGt
XdMgByDlGFa9aHN0/FyjY8YMliBPu45iFXO0kTUNFWY/Mh/HUoCUCSJ6EZbHHUvD
Vaiz3Rb0GMCzW3xnOJkFkersab74iwuUwEaIZ6nEy3T+ysIG6DUyawCIvIOy2442
33jfYDo4vJmcCPEtiSV4Utk98dbENazmNlDQ1K6wgn7Vmickmgi9YREiQ48CgFvN
ZkgjlWaRD4cOIgy0YbAy8HfrERkQmIpznhsPBJ6zDw5PurXRV2XlBjZrz2KRP7gR
d5UyYhvWgohK71na4VCUYa4pmWE7enEzviy4Qff55xjfuhTLGHRuBc6nJeJNEAqV
5AJ9HhQei12FEIpBe641ILuMn4gE2cETbWq4gtKw5lqP2y/BicnUfG2kBmur3Y/a
MR3202J/k8tXQLupS6FzIzOvyGYPVbA/YcH+RPMBcmMdz1B5Vj2aGkszi4UM7bfQ
F6Md3Mtkwa5o3G78QQ0gefUrjjJTQG2dwD8oH7OIRcbNtCeTFFr7Y5HM9BiikwAi
SQhulSXBfbQNF2XmlAvvdoRawfrRqPAXHjR3Z03C5g9JzjANXoptSYgqWGVSV89X
7J0ot3CPAozYKrrvK3pvtWpSZsVK4h+7joyTAgTgu8PdX8T1dfWjvY5EQ9ucvDHK
TCQiGizDcYh96726cRGv0S7nFi9q6jJsky2Mi3/j8ZLOy6cQ9eVyfZ6FBfvbwctI
bwTUwGgFX7V0x/tvQYYPsDzjXZdVVEp4KYxMugaXBqzd5GEqqzbNjY+oewEf+hOm
VdTFdoJyzftbdmpolG7tIB4f/jcy8JxitOOOzmaQH6ejkZaWzZB6ANqVy1uJH5Ds
ryR2cgSW5YxOKpfHWY5XCHPg4Y8TsdEMqdsT7xvsCpmWI2FKwhQBX2vIQ16onuGp
tH56TOIlLqssuXVq1gAvsjBhZ4orKVKOx6gWCWqNw1blMKz2JwSyXhEWqc8NIWDH
j2OhLn0ti8ylw10MQByWtV3OnUUnEd1DNvJXU6Bj/HfbnAvG4aDxTDPFxmwjm6bc
SE27SUHa3frFMoXJsLvu7jwSQ8p8TxfeKzMgOYP3yHL2SZBmhPRBGQVAX9beC325
tee/lrIx9vLMdX3z0y9FFIwKOezSUFtY1lT74jz0drIXJEZYfGO4a+UgCqnUYU8l
KcHkTOFK3wpaW2JvphIEJqFUxfXnjBGoqmIXYfoTF1O4sIkm4fEfnm8QMrpOR+7q
iAqTq5/mK1jLyJgW2QB/tLg4dYHkyQuEjgq9p/VUmR8ZiU4hBIgGKnT4KGSWgrd/
1gu7vB6Hgj9giaVcdP9AxxV/rZnOOMfp71Jd8w1DyRcSdqJmLJzb4LRPMIRPZsp0
r/zgoH7zXbpK0nXO2QDnDMQOQ2S6uRa7+UOOmtQ/gVot9RLDS3VxG1FNpWVB3cUg
vS1E4WnWUdswiWDRakACwDvvIemSIx1tlVcB/ptT8KK0s9QbUeSNF2NTRWr/63vD
+Sak4oGFljK0loOj+fSruFK038gHwJUbV0twHPfcdFY5ske2+Fzf11OrRCgYIyYM
C5VvjBEof4JO9Frt+7bivQue5cns6kGiPbma4seo0mNJSTuW4x2MTZoyzkXfk3mN
njNpzKxOqnON2p90DWP4JuskMrYuWHanDsrWpMexKviEJ/iFx3nJjNZlB7IxzJgv
Xt3zBvXzmIhay6NOVDi/HKRF/lTLkVCX3XIiKdFgX5oq5Mg7aKR6Zoct7w5VhRK0
MrPWG6XORXihmDq3KkHZbhLHPQNnt6CF0LvvBzIwiEyJDUxO8wIpwrYEOvMf9AWC
MUWypSnoOeu+EKkZVCOde+OPYy/YDOEo4w7kmn5M/nZFhAR1HRUw1GT5yUeD4Znn
QJrtVSj06UIImHXiTAdJYu+NnjzEqqYGbDYK9pc1c2cZqc7Mc4bxrtu6mF+nNdxs
53pTO2tzx5vZ6MVwk2l6OEPo677CYJdHtCXqaXdNk+yMBcg4LtWa0a3IztQAfWpr
+f7yWDWb+8AziptpxRRyC1+R14ajYta7LHfbndkkEPT0mG9cB1+OaFk/AlUjMN/R
GaQgQrlRWK/EbBcQdwiiOnee0bILQqt98wC/rfz1wLEIOcWOFCfhBb1QyU9jihuT
h91BhvUyaiCBJunA22kvCYdRiY27oFxbXh1lco4oh9wKdoc/eHt6/n1X0QIxzP1x
5w+G1la0ejg0OEYx52ieuoMoodsdwdz6zmv7neaUF01/CrgvXu0NBB5+KXiGfXEl
3zzRmjTrKKpidZV7QvdibvU3heIpOUdPBovWu7b5qvkSK+6dc/cvrbtnpwGhivne
9ej1UZcMEv7vzz4uvMSNI0eQCQgFn5llkUHRpFg81wgenvvSVX7oreY9kKdSO7oy
m2F32YlG9XQgcEycERnJ2mn3VwJ+lGXMR/RmwO+IMowsFXVvNmn8LHCE06TYJddY
LQpWcOwd/KeCrCnVj/a+sNRo8BtMHiLYkKOeiWxkbIyPINWr4qoh09f/+iUyj5Uj
4wMRR6eeLAdWEvEWCvJkacua16zOrwD42cSLP4kshPzK00UnhcH5rPjJerHrDB0m
Vi3tGlmOModniqHvwp2jt/2ddvrxThMiap+xHmJBc0nsL5DBq7vJ04MTi+wHxAgW
gNuEmyrNBTcLcjpl3KGbEcBzrIjwoVFnVBRecjv0/9DBNz96c/1hX+BVUYSURTWL
3T8fqWJXhtxHp5mwOZjBn2eWBggfO/zdAAjsy1pQwxkzkpxaJsGyBvPp+2i9U0wN
zwZx/LRod2lDKDkoJOdZ/1gblknXkymgKAYe6yxHGfXS7hq2QR6tEelHDBSR++Kp
vTJU6aNF2T+GgC2Y9SIi1RKIWs/ue28kPAs5Jw3EKvHTRc7X0q5l6MHkar5i938d
9p+J2qFh+lI4v6G3XG/1ng1UAHjiZTPJt7Y0p8Ed6UHRBbpiuDmJhAFeUF7QNGVl
Mb23+zxSMYCj3U3fdYN9W4CQwaU7rVYxgATH1V+r1JJXjOeieP+3f7DwkQPvh6nc
6DiamjouNeVg3FUWk7h+LNqos8arSp6slKIoRlvVCBqZp35jWr3tp6T8oRznmm/b
dM3mKm9NvgNEIu5MF3xhpeg7kJWJLLN8GKb3xh0b504LMv6acElIsHyCihNN6EnB
aRSuz0JpM+zpdbu6cw85aHp8OWoZ9EQUfirOA3rpQcuzBc03nYfEH57zcHDAK2+1
wuYTrI+Zo3iJMSG9+WJ3NiIiQf5W9L84P63J3w1hx+odg5Jno0WNgRye/FoXbB3c
Dk7s8vp8wUyFHIed5aTReUoc2kc5ha39yeVnXInqsZp1g1y7u7zjlaHN+jc+8b2L
VjIShToeAXcEJqt+oyhakw/8it6vCXHJmhYLbZfAqdWAYCfMCn9n+jbsn4UmlfnJ
jSJZxrG9GQRK6GoW0SW9PvFdVEVfs8Os5n6CZdfDF1eey4I+K+Bio6DJD5a/DudK
b+A9SUr/ovP2tLIwwK6WM0DuT142B1X/l08nFK+vr9Nn3rjwMMe0cidtUazOG6hl
6d3iIoTG5MH8clGZWvalQIgJNcTGrBpJQHBBnkkDLJt1tm8uSjgzd3J+HE7WGoJH
bgLAsvJV9dBHiXyRZAfx7wGnGDcy/TFyFxa5B+QD/lF3AIu6XQRRshdbc8Y020TN
fgIIfexjQT6UJRH0Y/fIiq/sWNegX+piyBE2w9dpqvTBnZwSArNRRtpGHuDj1wDJ
OhAlLNFU17eYzyqi6gnT6UZQJeuMUFhOpZXQdtNdgcULfLTRDq129mlO7vg2csD8
+uriXHtd/4Svj/7xxzWEW3Mu5EpVG/vdasJRTbVvcTDjx7ZAy+OlHfb/nMaC7HXE
7lO+Kojp5jB+OZwBoU1BaWlDWz8AHFSBJIzvy7OjO9VEcqiTNGme52MzGyLPMJOd
jEsNdJi8iHM0kWphdbziHmtylOJJqqQ5nVHMn3N86ZQ4BDrDeN6UHwb2vVIOj/Hc
bw/PrEDI8jYbbdRmwjNQTfrpvslBXUA8SR3YnaYtqoEWK/Js/vk7kzxJ2FTRJ938
U9c2Pqf/h/+zO6ahZ4CXfFbT7VTF+qf4HMZRD1GJMDMisyTCu3rGYXyqClv7+iwJ
o2yxGb4YMXvWNqYDlYgBrEWXqGw0YbWqf5f/YlQXnUrpbfECMEYdCFk+kawEvmJG
I7YdYC6QV3PVqpLLfwGG2RM6pGR8aZoGOyqmq3xZ7+qTeA1N7h7J1Ta8xIwdyLai
qi5nGNeJZ+RDWbGKSVY/EH3ADY5jgRSKhVmIkkE0ltBl/LeA4SWJndt1X2XtPyhg
lpuEjXt59ThGHSdhLcPZL853TEMzMlGltXgF0N95oSv039oeWGiFF46rPNMB3av0
MNbEGC9R2KoXQnOpGDBM9aE1LuljTDQ9VH4i/AZUmeAGYIhDImVr7y7vMMinIXwT
7IPOnyy/YMRgTb1XpsUyMm2UkkdT4ZweBQUyGs72sMKRb0Y75YPsKI6Xz3tnoQuv
XpHQnPEIJNycBLza3s9ckzJNV3oV7GAE2T5xzWFLOomBwGy/43VtPEtP/lhnBIXy
IQPQ5UzOjW8LUm+F5HAplC4mVLRQf8nONYMqHSD2o/tBt7vN8vWnYgQZE8eamB14
B0dJbo7672CvXtQbqVnSFSiId6xp2ez6FbU0RpAA3Wah5wFdzWJRoiZ9vnnO/fNV
wPDXRwxb3PceIGc9RcV1iDOZq3Q8KZjS5U6+bl4jNftMEIEtkPl0M4Jp+MI14/jw
w3hoMC7JhG8ZdaaKSbqfDz33EdWSPUTIkzAYLTc+ssZQimOOszH2Y2AEUDFAqwGG
U4Iph2S9VGyJZSLPQDfLHrJMkqRAqy8yKmB/QMv+EpUqpRuD0cgaHXGLw7iQuZ1U
QIX/rb3wrv3aFH3H1xXM+6jASBa5ln9bQVuxczJVXdm9KtoP4zDoalI2UBHYcDH5
ZjVE0GTQWBN0qtaLq+XVVEi5cDpnlOOIfR4VX3O/xU5FCKQLz58XKIIro7yTspC/
eiDpgjwiKmfmnaTBKPrjFG41LyflGzC3BKj0Dcj+GJZnD57o34fg0L2KqOsal4lI
JX6WOxS9E8B6JVQnqEPwytp8qLtNU8xGR6nitrUJsvGHhNNSqDN5dl9RbAUUvJSW
dLpNi00GKwwoW7pCIT93LOMbqkSqYI1vQS5x3UcD5fh2CimDBvJJxwAvv4UCwS6Y
9YbT8LU0gVK7KRxWUevIgyUDQ+NTRFrupFHIKNloBgFinPEY2swDkpKZq5h+53Nm
1j6XoTt7anC6PzpqbtnRJnVfqomZTuHpCk5+n2M30HRbP08S8bY3FJp1045Q9CSG
oic9IV/SV2BCKqoq70g0XTMfsPwzmCWBxB473v41yqZUc3XeM1vNRWly0OUSGeuT
ynSVBv6CHEiuEBjsuqv4lQum3fkC7tpkFlqiz8LmaNfRzGFB0yedF5YMJyiy9qqO
uKmBJfl04tW+N26+l+c4wWpOuAlx0pQ7c/FbCMvxm3RIgz7t2KSPFkykwGR4ZR33
4W9Mt7O5W54aKe2jvUMbQbYsqrc3BgWJp2YmpS5XfFV4aZtrgmwlEeRoLw0E8eqZ
VQPkqZNOYFYabpZIriHrIq5xlXTqbJ9d7qBZWnOSAONznM2n2lB3gXj3/qNfP2EQ
2dhyrviXXVr42Cwc5LCpxgffldEqOYdA/5yH1FP4k25s0hCfdR6U38JmjH7RBqdd
oPc91kJ2+RKJKlfutn5xGEPn3EvnvDC7NdAdnwIiNmSQT9NThRG5/FNVV77p4aSl
ToftFrnIg2dZnvDM0s6dEaLeE6s9q8aKTBQjUEJNM/x0S7jYqmH9nbi7k2FnKKgR
+87aHd1dqL3H0/1gxg9NJH3bPaQMHuf1zramkeLctwIZrdcc3ZSfpYU+Bbsptv5u
qzUfQ8/0MSykm15de4SdxPwdu7dOFlsZ6Qx522bFjfn1E1Xj8/N+S4eDzVDvppQT
Duv7hVOC5MPCR9N30qpFswOc8p6v/I/IJZEx1MwMagf15hNU26nBKG6YRnpF3wsK
LTHbAHTJgmXP33JCAxpwZP0KIjU0MEPlZyLzgPgidMzp27xfFkaqv3wz/zYN6zRs
04zE6ZrrcOG6xTP8ZbX09ujz4NntbwV14zMOz/eB5PAND1UBLpTYxgymhR9KqO1v
SG+Zj39Rxy0pjHzuRuZOdeYfE93A7sqd5wps+ba3d8U08VhIWY4c6MXw4GiQ6drn
OfGNoJGdQaC7QFnK+p9FnEcHr+iEzcxDtyA5U/BkPttn048PcTK2qe6WKXD9ILUv
OqFfQ9gDEJjieaM9WifuGdki6Nf7SsNdMipqrZ7/L0IxqhJApJ5rXiiMobJocj4F
DKGOHkRS6xrtRtUTSEiEMFZbLJstJKG5Ghs1fEq8ZMrvqW298XjgA8h84FROg/Q5
n2SnEKQoK8awDCyWN1xd9XdALOzaK1jnXtR6b3ONOE7Ltrl2cNA1dLT2/gFHPw1p
HKOAPfdrhRPJA7hFNPlA7XFsOcchJUnglyTOQj1CYhq7s9qDzlIMrScNQE0PHCAN
bGqOv/L0FaP5j5a9WWgnKSFVEqOyDZz9tywyyValSEnrnyDggRxIOp2eMXh5yZ7E
dMH+IgtKYJg+raeIt6FjOsrkdXJWXSgt++DKzNwbhctQ4Nef2KbtOi2qN+YrLSzY
kemX9ZdsRqRk8m54B7TR8gDQfQ8B+uJGEs96C0idpQ9FiQf++vWbl9EITClxLEV1
oQimnUN891Sc2xOtde1yrw3ilwhMKjFRtmzHNlVsO9iH10UCzxSgDXojaMk4Lb5+
vGhRM4H+rvlWH0MJr2XKlXTV3DJXwQoA/BM4dg0faEcuyYAUhtVKj2LHnXfQ28jW
L48pLvkow1pLc/ioquOgESD4MevK1s2WiCFyODfpktisD7KPdIrOGYPgXA9bBDsI
QM87UHeYROsmOO93tlqTd7CCEeOcxVsDsXM7fUEl+Vx7BiInejZIQyDgDxgwXEIS
wCiEx901XOdahXQ7EGXpxYhBTiuZg6I+lJKMRrTpMujjaWRqgxgnWxRMxgayRBhZ
TXvqGAsoUc8xpCdyTN76KrJLaUcDoz4nzg4Oc481CYR3LRAzjkLkyCceQ28aAhxE
fmRW5eTiz0J5MjQtlO2aFxgA1L2jKPqUpZrDgtXLC6ep0qQEXDHcoYSA8K8IDlHx
ZfagXzbuby7eDZKqXpU36bm3mqRpUNk/6nbw+mraJxV8urvnMg0kUMwcl9V8sEIa
QVKgbO3j1zbQBHIETgP6Q1DZ0FVrvcJ800lGwaC1WC6tzE0A7FM5NMQ/8F33jTCH
bhZiQdzSlHsahrHH77xGGYfwBbTknR7iM3P7cgEc/Q4Dp3gdfA+PPOQdln8ej6BR
CO1iNFmh9r1thSvNyeoX4UnuMlSfQiMUZPgR6wlfgXFQw3wUmHGCbmn7r2FusqUI
ZnUlFQj/OG+Az3u4mqzaAfS52wF9P4Br+W7owjG/CrNFPX2M6k+HwAGyICB5j8Zn
F6ANosp9gKNaabfCMsO2eEwS+1rVzGeDvIwKMReQVhyMLPUGhKVSiEiyvCMj40GI
xCQeDxnahY2VQ/FF69qoiUr04BkCGgA21Tw6yw+ljKt52AxhRy11qgOIXfh9wnn4
sQEEjRkHbsW9eZFpIHluq22o23BiGeGUS827W+6ZGpu3L63VZU9jPMqQlbPAINdJ
anN+QWeVcKE1Uunz5xvRvD3jBDvj8eZG/DTMJh/J/kblojSUCce0JeeP2u8GiH+b
8N/R6al4qp/N1zQT+T1hKZLnADCExJHe0AY3+Z8igTo1ia5yrq6+uJkvXIpLE+tB
MAwGCZQZwglN312Vha8/Uy1gyPCbm6uliqoKj/rbIYA1KA7plWSmcsbtLw8CXyoU
SCxi9oObP2szF1kxe0YbB8qO+oYd6M0pqtfyV41nGb9iZrR7QKNIC3VFmYr47TpL
lorPAlnsN5EFOkmt2kMEzfxI9GDrJtSs/kBxIZiG8sdrLzay8erAwYCtU9qFSypd
qzqzjpI5R/WpkHaxcvDBmT2lJrpTarWmoBi3Yle/wgAmTQLkPe1aCbBmNqxg/I/o
cvaLTQaLIeoSYYZfTQvlI6sCaZ7LmfEbnlnIazYHjHfYHSxSuKFSMwyo1JSzgxtB
sT5u6RUbsn6lmaaim3BFM5Rr8MCSbuYsb/v+rpzwRla7FPfPqmaLzrFzYpG75I84
Z7OuqNN4Fnqo5M1mmCAZrYOy1ZHfQEUarbdjw/J3/Z06ZBmPhD2Z1fCPegnTHoUX
d/66xwPLx7B1QEQ2LrkYLSkc2VTIch1yqFPSdViZJXuqMKCCL2SNhWs3ByrnXqpL
dsuijwDf3o+KOV9TtvM0pNOaC3W+L0Yqkaw+8OGC1ytT8e5b1kO82E8tjqtBa1dK
BAbiA5/TJEbvWItHFMtT6CL13p9vlL0nMXAF9og55biiVmxZT5GRNR+X6UCbgrTo
Pyihy8OupNs9HXSBF3LoBPKQVGnbBrf9guNyefbRBuywO2wXJf0J8ExjI/I5FsfX
sFKWOBnbVr2b0FfxULtGyKz0sg9PVeAzq2+vwCWDbeT6aKFg//sYL/IJTxbEmyV7
r3diLDqc8XgPIu6X/nBA0lR8SNQwLPofSYgWfGcy9U9k4U6LK70f6IrcEy7+7x+E
oyRXQqNmEJsC0yHLHIfBX4w/w76K7/vo+q2Ut/7DQIMBGnzioP0FE6fcrUZv+jV0
kubw13pHjluZPDAysY6M+aHYSr4meCWsB/iyQ0OhCU/55gm31iuuWZtIcTUckKec
dvy3sfGbQsoEgPWJvHvATBpskcKIUNKRZqY+2M7kvrO0LZjI2K+cZCbDIYVFhIRb
k4QXNsHAf9Ns/L4JKrmpSnTEjCrIpUrq4fWYSleojDtxhn9im4svAH44x7bWngh0
QWdbmaGnu6BvQWmbYQdLWukGlznN1mQuWYuJ7lS1gqRAUMEtfYmTIFQnF6dWBPMo
EcMCwlZTRgM9qc8I5Vqj9Uw82SxCuffRt5YROilkk+blm9sw6hLtKVcUkxW4+vXm
zqPvVhCs54Bcb6fWn9RY3d01pKNglZl2E7gz9G4Vz4LA1WRqukDdqVAGCqSzDp+K
vQ/OLaX6Los8y/mcxHkFOr5m05SpTB4mIrYSnwR1MUaP2kWDLcS7k9au6kLop5tq
5De1itPtzFUTZQUTuLc2mKZtV4lk5Zog1C3eKgcr0CuYUQpPbQbVpzxbGYxt3+KO
TE1xDl9hlwdeSpe9MG3Jdz/8MojOnslwERHVsyW3pHNne8NWK9kShxvkvIfb09EO
DRceLO6/Ji1GEx4NXjYniemUg68l+wXegL5tEvKXPQVhB5GUNjec/RZCBzUUvFQN
cjmXg2TqSrZfOLITwa+6I4b3M6JN+8iu3ylWgoI/9DMgIfMk/P2bEPWbHHrrJFU6
cGy/AtHz13jxviNN6LWBOkbScelPUsR0hfXDrAIAueVd164Kbzlk1qt1ZXvcQPi9
1TNYqQ/dkenqjjoY0Uw2pGru7ZeSpP07s4lbNRCrPv878CX8VNPLNxWFSvw+1WET
FqaFN7aEMfYCJjf69NPEgCXnwwS7bDvK9p6m/ppKH93w8ybu0UPfBKaIhxo0oAYl
ZJkQiJUkQFJScBXyyHXZycoQQ24Wu6FkOyuJK2453oElyVKEZODpa9kXrIwlqsgG
Ttsj90LiDis+9raxAe9cxSQqKwNJyDOmleWaY/QvvNQveWnXZE0NcIi90Fo9ZKis
1JrmPZlWKhm4h2qJSJz/PhRAWD+rAlMn2ieDp1L2BQvFqgkiAbwFuBB9We8FANco
94WXue6WYWArMNAv5jtsIoL2ujwS2aqqNMt2FA5KTOJjB0WbDUVlFwurgK+SHsGd
TRX2rv5TUZMRKo3MYRMdIXQ85VNmXc9Vg6tejOCDgWN1VQr3chJ+B49Z0Se9hyaC
+gYHQjfM8l7sWoJl8cW/kja2zgo/xTP+wJhnjj6C1YJLdEcI67YInmoKzeKH3Q/K
tIdimTjje+FLMPSXlID/Wy6mjSqLLWs+hBy5HgmIKSKZEA5+I1zgngQbqUT5ZGob
p3WYhEzGCB61kBeUB/aOQqnKotAlxBpRM5lXiUQO4iy5BPD0FCK973SwXpvhQH3U
boEF6zEJjtx2voEeaR1uPgw1xjl+VQM9ppzZ68hEX5meu09p9sZB2dqj3WjaZ4Ks
rWs2ltb6qLe7F4OvDgEYEp+dQX/P611pTy1ECHM5WcokckPpgHOEB+w6eYOs1BwY
fE+lBAE8PFISnKuOXUIDUQTXkhUHXoXKU1/bBgVMovr5ebBbjnA8r794TLMUT6Ob
MIzZz/+rkDShl0ixdaUrMCHC99rI7qgagsRPSKW3gLVbgl9Q35lbmw0i96bwsiLJ
cmiOsCIdsdUqUmdbjQXN1WNtu7SzFstvAmVtcPAI6pTQTh9GI84KFDlRAt6CGPKI
Vznd4CBBZFl4BE3I9ka/RQwouKeD7ug++VCiDK7gdpIX46R6OqXzSKx8KZWIkAtH
orItQ3PdntchtQ31UWHmEyd0l8++ZPD5SMxL+LqSxDI6Z6j7DLB6PkroqB/MQgw4
WWggpY4dPo4d80m86dMCCor/3bBTE9ctZKNfOT6mSSp29tlsBE3MRykmrXUFk5SE
G54F2pJLot/l/akW1ZlQcpDgGTR60tTTKpNOsa1ozv2P5R6T+aXstY89/vZgPZqc
V09lIryycLu68JO3+LN/So5BcrHZL1R3vl+EzUhp+vxoecfbTxqDcTBD6BPkIgg7
nNn/UGib2iwfkJCECEH3C8VX3Wwt8k2SEXObTQe8TW5yNfa6DN2pV/EYs90p8hK9
9gHFKBi4C1jons4e07Ke1sOUZWeCmGCHdg9hCM4bxOIiIB/NgGsx/EzJgViLyJQA
iMiYxGaulCNvjcTuorkhSZd10e0OxprqSENhDhul6q2BMX283zYN8q4xz6upwkZl
fuF87fjngaC0l6Km/JHuzKa8y3vUg2i+8082s4T8dWFucAphP/bhLkrXBR42ZOQO
YDrafXyqYnH40C0F6iSPBgqLynD01v3mKYk+qZ0TVKF98gPdIcocPecvIgUeFAlF
1sjTTUQDE6SDAaFmtIoCXm4ScGVbuoP8vdYfv25DHA9Cyvz07J3P6Yd+vGqmUrOB
5c4kVrqCgDkRhB/QokFWUG2ykcWBHUsqgHyZ9DOVr/rTxf31i6Zrxf7Q+nuT0meF
GQskO2Jw7QAGCZwfvb5GNSXVQbsnJMyH04+6E1q+YHAowTXKeVERIKsbXRYevvZj
LcY4gykpyCfIwl1BMNgbkPzkvf5TgJqdkT7kBq4WrlZVwok5DBjjkx8agcptQx0n
kGCjbeCbq79L3h6RCvBaQ1bPOlZh/Ubb+6uM0BfAUKdZc7khJA3LOsnmwTzI+Avd
o997/ZqdB8bnk9PjSCKQB+xNbQeQUNGJD/vqhux0hvWu3m5BrnUn2ea85i0PH5uQ
Tu6cX3atkcKPF3JGl/xyQabnynd6IzPEGAVMKZKxq2bGV9+MF6JWmBU+UxVoAxtY
SEZO8ufTQpip86B+MhIbFJJrjF+VQ0LBBRjimMaai7BqCl39d1Acq1R6eHo60iUz
DMZMG9efBkNbPQp+qxXOsMf1Q78OLfG5NgaTUE0FwQRLDpI7l+PYDHfyUx9YEXV9
cDVibbgeZWBB40r4AOXoF3nKWV30pfloBbTbgHuDLyyAxxGH/mBbF4A9fmcTKDql
kz31Cm1sp+8h5rkNR2SQOuqnRVi3NENeIgZxYnxJzGak0fNyeCSFMqp5pPtZOSHj
QQYc6qJLNIjyKfa14H3yXGsFNiKNgE1aRC9DeRGzEBbCGebXY8PviDZdtGCMhidX
zgPgkL/KQs62GQNBa4DA5nSiiMC3N1FUOW4XNaxZ+jruDDm5h3UFf6yIfzJyVwXz
5C8WlSI1wUdmksr5FUmYCQf+3KTp/eIIHWomzhfNBKe5zhEu1fPDLv1wL0pzVDyX
Ph4U81giGL5jAu3/RXRHuavypzKoZiLxaYzSGHj6R5igzxfl+d01bBO1I1oK5Q0n
dvDKquqODA/z1ywGVmPPV9mN44Uk9ZhQDruSNeuXAmCqze2AAWPl1L/etspD4zLV
mIRuxwrF+jHBVBPikOPQE2AKB+Zug5nxVI0xhgo1dMP1+M2TrhAVg+Nles9+UaE0
Ehf0TogplJ///HWFiper119vfw9f5JwyLg7APJANYMp0Mrp8WjSo9sz1GvJcD+KN
BN4SrBvxurjDoenNAI3umylI+tu3ii3GlydT1OUmPohvBHXRSJu4e5LSIpRHogPJ
4LEdaRMwMzyPN6DyNJtieeuvMyzSyWoW89AGq9WmsCXceaA+qhPhC46r7qI05zhG
0Y7tgI5hrZPLWRi0SVngclldY3EzIZ8MORD7WxtkGBBu501XMaoxNfkAiZh0Wt7j
7v1B41uwFFkGdaiZU1LSeqCaT3Zx7WJC5m2Jz810/D51+D3KKby2j3vReyNSRkC7
wBqyCuSkzUPKZnam413XZU2lK9bARgfVHxPD457IStikNU/zza5h4ytljYgW1kyV
W0i938fDdgi+p7S6h5QEJGUUgFvabl/ObtyJ8XL5dtm1ugLdnGVNaiS5OYeoaFdz
0rx+n22WHR6TPapU7sdqGGClLKKUDN9OMb22V5qY1hXO12q1U5iVDo21fTSiA52K
fHGOxxF00YaEo0oayNOUAyhx9RDDNXtbMWzvziVTaSgYpoEu0YtVK6J4jd7PUBSu
5XRDpdMUBs6ngX/ZyQ3gLOjfXtfFFCq6AAoNQuI9oAhF0+zW8VD2Q49i6Fhc6bXD
WA+usWCJC8vAjHpEB4+FrR3dIkfb6GiCCJzUKPINUIKDbOhfJrRJFkqhlE8kkEYR
Ea6spLpPMws2TcRf0/ZycTIJFPPtWfO46LDkMfEZ327jBVoOBNCEeeRsJuaMhwuS
GLhdauR+d8KNgTXhodd0qWSpvJbkl1JRa07vvG590vcMohtYL/uoPee6bpGLPPMs
d4QctcE1w+2ER7Oyoqr2HnIi27VPbv1bJmEva58U/BEL4voE+3aip9SLGkTrjOGo
w5Y7/+zb8BYaPE8AHyYQpD8JgFnFr8W+brWbcPmV97Gs6lm3e8fF6scewX0mRMWw
Cia1r61mkqFKpN2j41N+Klp3osP42OG4K3nxLOB1OXNurhfGzZseUJuSaooZOkV4
mhWRltIYQ9CMTk0uBC7+Sc1fUyFVlwEheus5Yn89GGvKKvcbozV8dnsKARLkiZPs
6nmSulcjS4w2ywmdz8uOaigX/TSmJ3a8HxOSX2jXemRGC6MyIvTOpJtcxmhuT0Uq
5z+PbD4+MMOpSTdlqXO+QulgfM1YrlHm6NdKEhxh602MukyBx2HVd3XaBzu+2zM0
6vfXoyMv9nNZTfsG97dgjqj6HYzHHIGBuiA8QKy8rVT1ZAqAOsosQOoC3Sx9xVdd
NJZNmlmL4c7W4nuDp86Kx2g60KsefvxDXZKvuZ1lsBzVzjB8Dh1LpvWIcX6ka69R
jZOOUQIqYr1aj6fDAOfoIrVcgMs931X0UU73wszBj6NpMMaIwOZZ7fXeQpy6Qvzm
j2gJdHzJpSsOj3UKbN/xpKi/vVxh2M4dfBHp3SlnUmc3XtoqH7BLVbZCy31JR/9A
AIoGIGB7KBMcNPfkEVTzK8eYx3dMUimEdhkAtaT2PNwlaw94WrEJrmZDAqK0uCWx
SbtFqcgXwKh+H2wVfbs5BN3UY+NTFOCUJyF4PvzLAYXB33b1zPye+BuwqZdTRgi/
CZw+iNhl4fbDPzB9223cNdFnuax0jhJ62btSw+KynwOc9kK+i9nhd+JuW/bqjQE9
OK8tvRxQP0h57QW4Yp6CRSNfpOnZTMTWdZNEG5wCjNVkk0b7ogdPHDB2geiS2pAg
vLK+QG2istBy6J0MhGDn8Ac2cevJPHCYowFZ2EDDTVqVhKRjYp+Ickf+mwFQ7/GO
FC19X/5yO9MfUbhTPiTYyMUyP5oxrKlqLi+cQSfX4SbZiCVBytAgUIoB6cqK1yN/
+WXa9709VJQTxdBvBSe3F1igZTujyfReaIAzvHgr/4Fw1cdPen51r+KFblTbq60v
mSP0e2qBTsvGGvZzrTr4vkXcgtXUsbmdMzkEBYW9nWYZL5nkIXOyc80+LRY+mYif
h3+DH9JBBqXhOTTdCeowbhz2J38+ktsTPAcIHcaFHI+dxLhkDo6jr/8jYBaMdujW
CmbTqPBZJazD6A1D53Gxkn8q7tcS96wR1HGXFL7TrH1NX8cALo++fdUumQsPvKlL
uVyjPp3/PXTryCEFTvvELA5v9kzgcPmwV+eeNYdDl+XGsk50SDhuCi9r1JJnk8xg
ijxhkAP8XlvTuPetU8KirDgpIdXCaWEVV/SaEAKmfoPrJMgwfasv4ah95QSHHP7N
v2IIpl0N92JBtciJYN7RUCJWBwLF5F8nkhJek/EMErZ5zSUq/5etDhf+aCA5LZ4B
Fac4ZAMCk6jszfjOtFbdDxAT/wQojpvPyYbYYHDHCeiWX/yt8Log3K/J/4ZCmy0Z
bXQBJ1xtC3NQV8LcO1M4NVdf0hU7Ml1O52lxXgTLOZD8AzCgJyyKAMA/v8GS6hzP
/ErBdcMG68xZs3VzVOQwCBgakE26LO0dmsud+OwPULHoLSHLHeH41ylg5mPefdpt
5kHj0rAKJM0jznDB5rdxuwM7GYijo0QGCVmnniKgInvJg8okDU3pMD21tG1gEpdD
N0DPKk0AyAVsiVJSKkNKCcmsnfu9yqmMwseiuQOxNnQ0Jq7TNfHAC1WMTM9rhoUo
S5FZgFHf7AVdEg8MU4ICqZFC1PqqvCrmeWF+XJ7hkC/UmbI3ho0P3S1XgmYFxCCG
kZ5zMAMut3Mj8OrYGN/lNSMJN5VVz4s8c6AYZJWT2emkbVXJrwzLq3tlB7JznVQM
R4uwW2gogNfpOfvXnb/xqf3ubuwRBnAK1KCnCX6bOG+5Zc53se3UsBnLRgvchLaF
k8eI+4+cY9aR5ykXEdFCN3S4f/OFO/xT/BRDWAfIx4JnU2Hdxf4uBN6M/vqGQC6y
cFbRe4eY7kO0hk/0A+ykNc9JuWeZSY3QwpFDfBIDfsqolsXLuKpMdmld1Bpnh3J6
EvCWIMmM3KO3boeHvOkY6NSRhbRyY44Y0C5DjnRqzgrfTQKUeTsJcCiXUfMYJxMK
NQnth7312p3qG0S2A7c8aRpdV9uOWgxslTbh4kaIlpvBtCi85APAbHgcOrpbXn33
pSEURXXWVa/GwuHxvqZZYax3SB332CfNJcTDuXa0ibZhDdYkzL0luc1roblj820c
A3DEJx5ygx4MtbWhMsbTususqkorx72gAwfameGa1UjN5EVdgavKJbb3q0qyBpnB
V9NgFqOCFZAv0phkILt/wWCtDknVZVNPPvbDVdtw2ssze5h+WOtOYogngkX3Kzoi
yDt2lb/ggj8/WFHWIUiHJUyvjx9UUr4ALAHDN5bumFFUP9qP02YG3q1H6DvTobTK
yc3/J2Q4/MDyyqdgXeJ8rji9OMYVUCR3KCTQGahauJuw4O10a6Z/pDrySIewW+T2
xGFsxrYqnAw318G295W7LDfesxcGskF53CdHCpKqwprLdHWSznYa5OeFt26M1uKh
oI1qIrHEwWlZKWJciA0FyqNy7AcmBf/iuK9nc7qzrqiM5NET48sMGvAnSO+JLSOf
trv3glm68FQw3grK+3dxzw/LLNETH1eqLUs6HXZ3tWdgoSUEPGFkjO/O35gricq4
5jgXKvVXj1AwxyE+NlWNqMbv5NwmbLKM5jrS2d6B0UfLqnOjzNUv+Za13doOZh5L
foQlqv6XAE8EmOWvX9vgUGatbSLs1kVgfEhVJuaMZP+aqHDl4wd9beFsxzNbBES7
W6XQvJiMM6VkdJAvafzmpXwG9RJGQ5dk3FU2yDTafXcJVRKXqiIR90MF+Hwwy3nE
8XRrY1GYc2w15FytmW7NsCkbAu1LXdZv/UCKlmg5+al+iBZmr8hYAs++rJ/AnsTs
VMwiSdtFSC9gEyArJEyFrqhMGKcLdVmL1AvcSKUlFequ0uycnxodXCcACdJgnXPe
mog8+AeX9OFmJ9r21f8zbJH1PFU/7RcRhnzKdQMFdNAN2uBKFKTu23wfq3rtdpmH
AOp4QFxwNAi4EHCaKMfwrmU4QXIph5rK7nMautGW7GV5OYYsE1syPkHykZl3mXTo
XzL8rGL5mPb7+bsIKQP3zvxNntSlQ8gg8Y0WC4LrcnI5/466wf64ynfD01zi5MSN
Wmfg+dik7xlApQxJ7y5TXhCLd5WzM8Id0XSCpFdtEmegnT+uV81aYy81iTseyRwR
4qNhDkhl/EqzOAZSCd97wgdfpxdPoTkQCHQAAa2mSaJAspELcpMRszaIlxbF/rLW
lkIhV+uWZm+NnUwzudAyG2dhRGZvHXWYYdMgoZb8dZ26n6C5hNXvCKJfdXXhnroG
7yvjclWavuDvVlhiu0jZvjXe2uNV7ZWAz6+LLgrUwrRKo6v/WLsYzvHj6lcSXe3F
rpPdYvmrwrh9ySRQkNPSF977BG6ZGqX/gVosdLyGO9vSywZEwBHdxHTmXcXONCjv
d5Zc6WroB1S2uDZNskshT0BZCJukXve3WEq7De9alzZ4kJtGBGd+OkKGfqtd+d9Z
XHV3J/OZHDEaMSg/7zCHDd9pzlvkJvDFdwN4hgyNjm/6pq91F/53VHi36pJmvPgd
F28285YOqPGM0PwVB4rg601GwPorxs8JdXRHXQ8uzDUauRMPEuz9vIa9Xr84jZCH
g+/y0in8ToxNFSD8/20DtmaFvSJ6zn9wb7A3MO1VCGTj2mD1FDA/fBWSVCYYpDa5
m52MyJBtyCdQirBdf4o5Mxf4RvozZ+qfYxIrOKCr0nrk29/9AKdbV1sgyv8SdhHa
nDO19W57jpsJIdukV3gSp7CIGUDE8FzJU84IPhrGfo8jPn9LvLACvxnXstI0DPQR
RiPkcg2VtgjfZvJrioc74D+hw/ujJioyWH7ccdlQvs9JnWKxKkL9fWDoJ9L3+9O3
kw0mt7DFiTovVskABazObzLLWU7+dfd5GB+Q93ulJ52PIvhOyj+b6LkdGQKLZwcc
K+DXpPedyQSBaMzvlEaTvGjB4YFuzcNIyLVsoDvTAnKA9+bbcLuYvNNqe8enoC+0
1Pv4ob4iSTsod71IYX1bS8hm30Of1KE5eYKjzm5u5eIJnukrZkj2iKg/74K2tJhX
vZk6uxfQswMN09dUO+JEmP3YLx81UKN40athH8+AbB3ijFe8PnCngukB4e3cYt52
wP6ozYDBkeknl/QdtlvjunslGpZmkXju7lsv8M408nHFP1kHDUDj1BRQrZn8tCRO
XoBdmQku7EwKqni0wHqmCqcENjF5KIZ4crlkvqCAmTrudhbHyb0K844PCmA1Tsbi
NqiQy4rVbhK4M+0HfUPRnolPz93aMEjhpsnNMetUzwc+Z5ICVKJOWeb2JN7yo+VX
8UBjywH0TGAuuuOdORcwY3fgbJu46SIqqFxJFiWAGVsKLLIa7HuwD8jzcxUWf6oL
CV2jfm2brCmcqmgzvKKN79PVNI5Cv65RxSb5Yljrr7vziVhepXD+VhbLmLlQnVJn
PwY3AHyUKP6PsjXpt8DGPaXRcX+S2z4wPdDGWeKU9+xa3Zbi/Xa6xwDecNm0lxT1
kNzKoz9qVXOf06LibvibGbH7fFcVrwMVfNK57plsWrUKYlG2pc8gyK2f2dJqg+9d
vSMaO/QmR3YiYMuI6FSnxTGikHXNYBONuEuAZB/EzYevGj63dtSuJDDZ0CUXJM7u
QzOMOQUJ5e73PVC0THtxQZ9ga+egM9eY3plCL5Jf55aA88kvde5aKzpS1l2EAch3
6Dslayq4DQ16HwlhRpzcjBY+XZ1t5GVNcabmC0Qb6wricefUY45zOAmfvpkOJyJ4
Kqgzdb58T0mYJksW6GLsjQbkVhgy2jaTXqi3zIutvAImSvg3/HxEPjwXTdrRIuF3
RgSwHBfC2cZlpQNcw/UIlPs7zPXQ1yVOFEgpj0O7PvdiHuJ7qjqh2U/1BJuCvYQi
3orxL67YiqNK92S5e7HSKm/V88vyGvtGVa4CxCZLA4hfi+zGBj2Hq5IRKO3OtTOm
Ao2eQg7Hh1djVyjtFD76XYxkCkN2ShnvnRDc9FBi+Cng7eLeWTfQf9fr6Q9UMUv3
BaJAEsgNK7a4lLupmasEUx+Co3OdmKZNfrxO8LWyLChmRlT5jmQx19Dw/W0lkDqp
gSR7OUAjZ3up0OAbJzi386VQQ7WBppzq5wUbcp6I/bNSYlueobJYux1zgXxs6xnn
h3KFj0k+wvjHew0CkBc+rvwYXvM7nRJqlThAlWx9nLM7d/7O/yamYHDudtkYNqEx
w35aETx3gqAo/tpkqZKG+YH+OYqEieJ6DhYxW6/EdD0xZW9c/7jJIKapsb5wm2L1
XZoiUb2uDB65A5d0HEFf6xMfQvfRkQTTm3lqc3nObslqYPF0UQmkP307pOGM67Th
IHLLx8CnDg9Ct9lXJbLIm71fHdGmbje8exomFCjFdf+CUyUo8qdwniQoGkQvEioL
b099WOxIl5gD/mE5yqeuGJpGI2eyMkQRlMGZ0FqCfNtzSbcUq5kNzdKW6dm+LqQ6
4YWpbC6DxTxx6vF6rGcYpJpVaca726St/XASWKOATh2RihfPjavEVrJewBuWbxsW
ZOmp0HzkYbiPnezqzP+J1195hMLRVdZ7nXkxBhwLGBBQYaFbvfCmhedAwaenskYu
BXSP4TzCkrr/acQn7mvqQIPKOijit3/iDEYgRU47WxOwPaGiTj1nCfRUKeAQKcEQ
L/I87XMRXdO1zwzKCpeKblGWSI4eNg9arr6Xu6XWhbCNLqy/xCmnf73NykQJQBXf
JrAAYrU/4wkVC1+xoV46EmhudxWsGMPSADsYKIU7DAgkN23LAxDATy4Ngf2m5X5X
aJVk6/lIMNeNEJzM44acdeDQ9KppNclx47MrEf4+NR2Xyumse0gvdKEJ9P6d4ueA
ENzCYEsWGSbKpry6K7Pn6W2R9D1lA3gL/09/PYC8VU3wyoIlvHEpabVf/WU7Z0gT
MONQDjEZt29BpNexa6fYZMmmXBUfPcRmt2HxI7oj897M3y99wu4eex7jP0q1jqdM
NPelCReqgK2S+2QmpXQG+EWG893RHT7nYGUWrlsWQI+QT+pT2C21AdNGZdo7XYaD
7BIKF/fyKFBzLPuXimHPu+X1aVVkjZ6eW0E7Fft+7RtcSp4JMZwEfP7zySgAMN2d
P+ipErgatZdHNKdImD+Am8nj01ekMrdPWQYPgLcy8Wo3+Y1eOPpeHss10LvlVACE
TQZyIPMMqNZY9SCxGX/V8ai7WF0J4159xS8y29DCvPuyQcNcVxDCglgyoFM2FTcn
fNmFvJRPLti77DxCZU3D+hlXKvSJCWNj9RYOb1JxxoqfskMqokMxx8G8ArIWTwQ1
34rk5RLtU7eHHH8MAa9HFf2jEwkMt61cqkwnXx16cddog+7VCsoY3OrhAyWUSZIb
wlXPhdTVCagsUL/aPwpsghypn4dDDQyOxNXv/b9SC27FLMwDN26o93fW+eO8kU5X
jgkakO3gCUEaLJ+wbeGDGVXK6ncvGynWDy55xBOF6zU/FqNvFBzRa7oqq6jueYcp
93V3buh3o2WIPXHRESS7Xb0PVm0FA3fthQZFqNDm3IkWtQl5siXnKpwOEZzzwrTy
hpJTS3wptTxbvg6nLAqL5XpDS/+9vJGI71II2hLxnEeb1LXBiokfejOJizlfjEUH
/zQa/TrHoWExpue4bufZ8FCjvoU4yDIKr/gRLhe54hEE4RVjCaEs9BwFOGNxsRvn
aW0LGyVFYiX/XQShNBaQYo8gE5B29yHLhKkrmCeGRab4h7anFLf2RSJXKWcdJcSC
AnJSujLIE+Jaczv1vXUclZNuFKZeOutB/oPd2LVxANlp+euaVobalfZrjLbLUxca
GE6pJo+2ZU54S15au68/rqfcp956n/35JM7+vsAtD/mR2NmZCY+EoRcd8rUBtEJl
lIRgVxIFHSjylIquxuWuhblz9Ovh5qhtQStp2wahwZET577EfHkWReZIjWMc0Y31
8N5bVb1v34SIRAUJiMrfBMuxuNBciXKIbPqQgrQlPPmIJP1m+E+wsBVxkSg6zDfS
EiiXTdxrOpXWZe8EGWA9275jkTsF/LLKf9K4K1kZ3JJcR309FeiB69ZzHmJ4S5zk
Ho31JgkfKjFZ4Y1++JcWpkYdrCf7wjfsJ6P5xBm11gA7292q573fCI45lItkAfvo
LpZ/y5OYqi/tZ1pBeoooModGZyAzRuhi/M8Av+r11zpgAK/X34DeWbxnsa355U9P
aKvIsOI7ERPTp4VWOsz+upTUIeXZSJhSwhanfbSXu0vjVC7G8ovG9XWPss65V/7+
6b0TrQFdcaBC2Au20gZSXIMkRFhv9etZUGQl63JtbwxQ6ZxrAx2K3w3l11b6aKTh
7cOy3XBcVkYFvwNw7hwKXYJqqtzWALbfe1O5D40FmsxTRzcbZGNAAmL9OBeTQvaG
7ae+BRvsz+qwKAWWVIC3bE6ImQ/1PnyaUk80wPXrUrsSIE0fpyQ96b9SOTs4uicF
0lSSazLrJ/ewn+4z0FUvfEq4n8sAeWzUvCYKmind32DTI29usYl+/qdZHREuCaM9
KO6R487jhigzpYngTOySfPiiaP0RzKNHRgzebIMTGK0VVhzidLv6UedO/K9Gx3qB
cXoI/eqtKRPz828ChaG/msOll0AEAwzgxUaB5qvm8QZcNO5RpKUR125jU6wpuK3T
A1iYout01Apqg2H/zWc4kYpPEMlJGuWzPVQyF0gAyVtrlfjLVDlv8oOICrNKLviw
meZwfmboRyEJ0r4zLoznT8gMbhEhZDmwDWBBptyGfAoFCzu/PgaU/UKGI7TKGgRn
ekTX7IGarnXj6yQnWqP0AoGh4Zj1SS5Gm1gTMCs5d4OEGkl1sLAk7YtzWWNVo+PI
kk+OIUoblkR/Je26Wa0HsGJidMDZXGRbydt0rImC0sKvXAS5D1vANjv2rLBukhxI
dEGeZDl+wXu2eZBpDph6Gt+xLvQ0mnbkT23ruJYd85l51+NP/7aaKg5RjxuiC2F7
ZJ8AUbB+69v/4mC28+6Ajd3rHD/ImVIYLzm9mV89Cdc8gZzr2dN8Jnh+gYdUPnBW
cYHBrNAxg4l62tnr8ASTBRpvfqqL+9Z6pfnp74ZSHy77IP8vycrOsQlsf4jOcQFV
tYZyqBN507Ens3RK0a5/fOMDuwXNHMf4GECLKgIr3AaRZrK0x+le/fpNsAXFZ5rd
cvXDwkTQODpLR2yyT4omdignW60fmd1URtLEPF/rCevIotRv1zaWG0gLzlYD8KUI
rhWcqX+ddo+FI98z4ASSKrMQAgeS2dAmes5b9GAcbcsCpf5r8oePvXczugJtLgSu
FO6vN9ogGzkKXwM22e2IFP8PNBZ15rg84nJ0kChecWf7PBG2oc6iSUwoRPtRW3Oh
wtmi3/dEDseVw49vKt2aGUzyd8g6E6AMebGlPvSqD0RckIbuMSf3I0o/givYzDLw
9NUFJ0B+RnVlK8G0xTN+LJRwCjT4BxVIRgKXvQSoWLgNuC98g1jPZaiThbXqYHez
J7n1YW728xyXjVpYgLW0o04E3STDYC+E3qO/5qrZR43k24ncpwmzBGJDkiy18OFV
5+uhFcnmNm5Njnl1aUdW/SdKdcsCDRTb0jhJ+49QGfZRayfvNy2s2+p40iRx8oFU
4juySAYOiQv+YmtMpCwClnB+H2Ew351TW4of9f18x8vzBxsmOseU0lw1H0o1Og/D
Hj4VV3T+QHZzAGVynKU7V16gnegpI29cIgr8TGu13LTcCK01spsouT3sDiaJSopm
zhxpGwixEx78EdEJM/7d7wgIXe6bm1nMUoD+bNAFMFQuMlzwr93t8dcCTKVgkRln
3B56dYnRuAUo7VPM0zWDwLMOE0/9lVcp+xn3iMEHHxuBbta3Su0Giguq4UCdZin0
TrO+r6JUxd99h/F7GUymUGLkfAgojMY8plKkxtPTZE/dyQshuPPfI1CfYGGdyzrW
gqiiL5SOduGmEqlMrFOII379bnUHADd5AvXNBeztgsQb7sHVH0Z+fklUlV6y8nko
fkuDn1gVmLBYpjKjHL9IC1+Yl0dtfA+s0B+sV/cfL3huFK8DZG/3wahZ66JsIfcr
Q4gbDXr1yhvCvVg1j243TkgQVSTWV8r5C38DcrEN2n9c6U4nGtJnFAW76UjkkPI5
oYnVHaXya06F+fllOkjHSYC+xEC0Hp421Dv03EVsmS+Azp9s8KpGwHekuhCV7XoD
vMimFRnm6O79jDZoD5Hlwof8sKCRmtXRezYOwjnQdyM/c/jtyTYwZilKhf8G05Yh
K5aUUpYVC6XvdH8L1XxhGVNi0flzzz6GNk21EanwzSILaezG6sfsZMesyQjmu8MN
FQ/foU7+hpuhVHpAW9o8LzZbIvY383QRG8Hq+j3Ynes85Rshpz+WSYIVLZy/zo3w
b+KNvqfOLPxsuTdHtZGKNqozMK0cE1jMpSzUGzDewSJSl7E9N36FLusUp6cZiARg
GYFeQH2t3inbRbyyX8+o3UeWhf0gmEU8lNxcyACVOHXkMJnj9M+L9QJ47yYHRnGp
79lmtdz5U5ymJxiE8QWc9mQQg6w0zU+MLCmiU9fYAYHS5aCTjrKn4Q5sVNbwC9hL
Ov4I5A3/I+1bWnFSR5Wjo2ufUzWcfWgGdEDyRXOQPIo27tdSOPB9SY96vtPmBYG+
qXnoV9L8JQKfSVVzeCG4qFfHUvY1uOyKzjzUaP8HkcizlNNrc9IRrCiDT8mpykEF
C/IZR0j9GZ0WexNSg3b55T5nJHIo+CVxiUfnVdRgyCWA/eqvxel98fHTnc2BS3Zo
dLF44IwobPxxDsKUMu9nL1RT4bYLquOZL5NvwPtwb1nALP+qmURlZCtOIOU1IHOD
KE6jY1Ni79TcjOJaWgz0vfNDspqX63ZpFELIO3P6GZm+Xv9ZUl85Kz8CCLl4l/1A
4DgIsDhaVP8evwYVxx4iC7vRbgLAiU4L0SDfgxD5AGjUVeiuE//iEYT/EBnO0xCP
znreMdjd9O+Dh0Ba9tXCDNoM4KI4oXaIA2HIJQ9XHrSdtt8bYnAzfcezwPuC7rYk
rLpcC5kt8XG/eAr0Mk06gSS6dAkatjSzsJVFBwojv9y5kbnlyll0GCF/x1fFHyuI
+OS+Rok/8C3zoGNlH7OQgmGOqI+vB6+dHg4+wBVv1OToLNjcQuG4ITvFmpGZmFjp
UIHi7CCj0UGYLlz+n+4pjjtdJrE2yhbr3bV5Vwl3MGWGS2LWkYFUgMPkQ5ScyjHZ
Rljvan21d02RQgSKenHTAkAfL4CFuIppeSE1aUsYFU5QfX65A/CRulpQZNel9t2V
+dfkCZ4nRVqMER9E2UqVfRK+Ha87rxvhyu2Ood+oOFYkmnvNqAZ46ZDxxDMJfHrp
xInntXHZsKS9oR7LPtxzondUR46AroKpWnGJojJtEobzYsvXbm1sIXJbg8aWTRLR
BJCP6bkrqS+TWmvdF4LcyWHBzOYljcXeMQvkovAn8475mjyuitcws1zitTH4LZX4
nqTfEDXE64dFr1JsAMGlEZaVy+WsJh+VJdU1cPfmXCK+HOZWxrY7Ue6zqX61DgFl
cxahdfmpifEjir2M86RKfbNTMAwongo5WtrMEI7muimvzS0smc4Mje5735kZFnFC
e3/+d2yWohEBWNVSmme/SVjvCt55Rt1EKBpEKpa2JqKrbcCRAW87m2qBNvaEQcaq
1enKs8YHZEdEkol5XlzIDp/ftq61xmcFL3QyLL8LMsh2BejrVDMYBzoeZsYPavvN
GR76us9T1K6GMswBch98SfFOsczqC80b2VX1/LIYoQi3F+uSVEPZcY3zFp1nhoGs
mB0nMRLoTjYxJ36j6RR7//F3QkLdPKWDP7Rk/dWMGPpY72JQ6P+rLQzDJf72DofH
/+8yY0wXdX+P7qYWYCX7kffKAR6QvXKt2Tvj+DUWxCcC6DZs6guP5c1p1dTpihJW
q92vLJ6oR5GsZobObAbkX72LKOG/t+tBQcXQAF8eG7Wrk2d2SmhzhsV5fqAYtJS0
44vYrFDVkJtbyQFMCRKrGS8quC0ADk6XjPCk4jHAubeAYzuHbpA2qmRPIlDnes2C
5SRuHupb6RciMEIKWUBy+mHzyhBkHrS+K3WEDSn/tsebEo8p3TLW2nC1e3UpijvN
6y7+swPyoOMXqMC4eYdG1tLXa5gh0q0RroOcf6/ZRuXiEnQVtzaGXetyn4ylbt/E
sHnTieRL8nzRcgWi0Drc6Sx8uofDBnvMPG4pHMT9wcZ9wxXYdMu1GfaNL28/lacP
1tUzLykge1+g4jvoFqjHLPSjO5b4Oebx1wfIUTuaMQAqlwMZxYfYhzwEjgwmS5/G
U9vJ+lxzCK/rWvo8LSS5U028CN67xBVz1vSouUBO5Lp5hxyY3JZapU3Nc8YM3BHE
GuEi8AVnBv+NUfVeB3Wo+hm+18UIuv4x3gZBuZzLB6MkHvI5OVtYVMw8WqmJfsku
ASNpHkTrXWP1R7vlNtjUtNl1KTRjEe/z/gIQpFanJjpvW9BHLwn3Ch2Cq8M4GNuy
PIeVtprFLVuejnP1Pxpf2j4v4MjDGqAs7auLJVFJt9xH16PAqS8vp383JwETZ1xb
dawglvjpUFPvyxJl+BDtQiwJU+kRtyDm7wdaq02arfSoXe/XCODkKFApA0yFAz7q
PbMbVtX/hNR8xxpVkK351A+2QGdufMF+8l4X5fuYMWBOIwRgC3uiVJ6+9xuHOlDg
qDN1x6EEdOsZrt/jL8vsFpCr1Bhoq9EiABDzvokt4Usxve8mM3kVBvGY8Pe5M3mk
inAL5lvHkAzOdQZDffVFBhVTbJhfD3onykchc/0Lr4MJtO3TK0uNVOjHtgIv/JqO
vNyJGfzAYQOU0Sx/5XOl8L668j21T8wiiFLlJoP9GGnSW06C5Y8b9Pyga5KBUqv/
3DTn4bD/fPLMKiUZJjPm0waOwNzJvFYSaxnQtICCq/K8kdRw4qCKuvB/FtOG+/9B
IhDgUu2X/XNMtk9gHwpHvXMn3tB9LxgxFxtPjoVcaY5qgE3X6FrmqYu0ikdeRTU+
vS0SG0eAM5O5oUJx8uU9oxPFT0cMhPX8Ui/wqQSLNfnpoI3OM7zPRMuB0h2+hgBx
vGztRMloLSu78XtQB9cY1AFhnbDjcT4mSfxlfW/++I00KhQHe7zkwCtwdCmaDC5K
BkDHc+QGlKPuDRz9YR0zw8/JLLhtR19moRBNdr2L0S0MOoi1krvFHt8LBZPt3RVK
Wn/genS3tpOneXgWg8RYAZV/FR3p6Lh70idNzT1jIjsRDCmQ85mvWtzstmzzPB1Y
qy33KfSwfn9XyKL0SOrVxhSJM61z2iN0pfiO+u2e5lOpqvonKriBzLWPyptQFp2f
/RV8P02f37O8DA6JAmlVXq2C5FyvxdjHVZpe1jgZCzYjde+Of53i3p7XD4CZMCuu
quYVxcCFoZSrheEpSKyzPDQnNO05PQ3/p5dyRpGzOClEZY0rDMm3qZtvK0WVslky
vBGmN7zrOP1PSRLDbKj50hxnIpHLvPLgNj4nIGJSNyBiRmo3jm0ZjJIYKi/jCC4V
hoDAfkuywIc5/QJD+/IAgb4eUpg0zTZNETsvTuwclTu41zjXMtJnWTNe5W8LPozH
Sv93hT1inEiQqg6NerMRPy1BPLJLRkyDA1tX/RHDmbIBTdY78BdqxeAcoCxJOV6m
Q2zvozebdvfSTG8O1kAm5NrJUUJjSHUomekYMRItTbH4MJGkeT6jEvLTQDos77PH
HCQLHzC7UiT6uZxFIzeETSRCP2MgI/F9sZlQlOcWjw9fV/0RArvEKuaG1y3eFZj/
P6lP6TSYtzIMmOUciXOCzl90vPwXuBalFvA5SdlvLApRkgQ/tNDB/DtG/WtGTKVs
kUUng+rN16B0FW1tF0A8I0dn8oUr++uIdc48QCgVm/w1Biq43gZhaxncVlggiT+6
dMJ/zfsuo/LhMoUPfyp/TddNcqT4QIFr8HcGlyId37gLSsSCAtjmH4y54VPHcWOC
pgHhOptylewA7XkHDa0eFZqcIO4OD36fTO0z/4TihLq0eOWmkCMv41hnvxGywX0F
VenHFFmaASy7/VzTw6gvZCUrqnHJZIJ8z8sl/6g92ci0JXv0aDlXSvS/oaAXd7uV
a9hP5UgPOJciwEB3wt4Xfa+Jqd6EFas9BW6A/VEq1XDMJC469hZfyfRF8Gd2MwJF
XwXr3URtliBHzlG2ML9uhvbpxZMxYo0s7e4eqVz940lLj6ZUSe5yMHKXF1YrMXQO
NeYH97a4i5nhCoC7bG37vBJFMNQDlOraaptlD1tUkScXrqhsOZArQE7YHnDdnCUy
zv5ff3g+VAi1XMChL8asRhkLX0/5Bk9NKeujl6NmQy5Ghf9G9/YEYudz+mxGEQgo
SNuFnHp6a3PUhzfESp9mLgbjumTdBCIChzTHZDh/aHKZmGsINNCjPIHgNqulB60K
Ip3L+lj75aEu3mol+gpKm+62RlXx1XxdC6Q3lSWDloCFCpK0m5GmQnhrd4qzPYi6
JLaSvOh44PynU+kuRxt9bNNRhNeDeQVFo1iaFO7Zw3pU2sz+h1oe+h/Kre/QtTdu
tcXAjExOztzr75XrnwOAVx6A6ByYkmGdAcF5Dl5T7W9UQBCNcDY6urWVaZvtqm24
gxeEFtYc/yMexO5ztkmyJOpnLoAj0s4qErFoE3znibHNMqRCCVuBbke3Cykwwl5N
wou+MHj1zsmWjw1nLyKoBSj6EjNeqihcWICvfAFytzAe0zflV5TnF8Cz2tGrWLj3
JryK3To3nR2+eFdd79YcQtKR9CFpS7Th/xkxvE227XoKErhuw6ed5FoXaM1cmMOM
9bRkn5dDDITk3z400M2kqUlorU+us7BtbIy0faPkG8yNS1xCzhbj56ufUIh9jZtL
pfn6RvkPfOAH53WXgNRk0sKS8GeVQyFBzgNDkQrGxKE5H+iWVKzEppfeP+73zgTk
9fE6w/49ibYsFAhnvOocYGnIoJ0qCC3kzP5KGEVAJ6YKSNM7NGlUFIzOY6Tmc2Mr
YFi15YGBajNVNlvfMhnIl8Z0kKAH2jD5cZ7Ipj0A/1iA+VdBuMFNmdc09h28XXZF
+7I1E6nGGQyp5VjDMPNp0nznXr9d2KuPr8mAraOqm1V3MdVpP/aRhuHMuDr98CmH
YELADAimWMCbJl7HNgxW0y5yXZ49HQAlLitv3a0kyzZBbdkeJvhgVb2/I/h8OCfv
s9HxfXWu3yq04DpTUuaHrN+rQYtBxFUyOItKdWvirM/bwo642I6YWpfS+BKykDoF
ixQ8hsaTpTXmHn6ICNCyqf8BdaRy+9bP3vhKF1Q3fFc8VOMUXFe+wpJSxWFPKy5v
eGXZgUxeKPdft9fGAcCzEwXd36h3mhr1vz7+kNWciXAtGD/jE76oxs5ZbrwT1rQo
HpfqqvTh22ARHnAFXIavDkq8sJtYP/b55SA3s9vmZmYmMZTjUrqo0mbYx3Uru8w6
HI73lVzmcLCqDIoBY6EJrT7FW35+P/clQ2O4eybp2Tq3yAvlaFBkaR6lTR/NkrBl
67qxSsDACH30ddwRTPXnVu7PRoDKq94qDz0bcloJdNHtU4Cwxbotaqg7aC1bd05w
8FGThZU6pX4Ez+l45AQ246fQKEVCQJJl0YdTwOSLzvW4xY6vk66+tolMNwMtLsNU
xcXV3rOwlYqDQQRWs+MoUvC4ZIzOH5PR50bUjwoKmMuJlHpHzPc5Rdfwufy1gnIA
pvdEJtNNKBEvkdXmneF3HyzEvayI7XKdU8KxIqIAPWV6RBPTqEYcxLM4YmaT7snD
Hf5v+j8w5/J1QZpkqsbwaM1VolVFcF3/MagnANK2+GZay14YPWbnGVqfhA4oXXnA
4V/VGS7mbuVNimWU/ofsW8Gw2Nb3myB6PcSvPmAYFcU7XH7Ie2QaVASGLNKyad+u
HIOsmphLySB8ag3LUxMJoegjDLVhdqWFBiYVnHyMLzyqkK4vgMTgHH54bqZkEoRK
X3PNKYCpvUo9B2B2R0TDpXXO09dqgNsMHwZOArJIJtGkSG9Qzf/271vYeJO3beQ3
f7mcP6Gn8ujrJnFHh6P406zbZQLuFrPQaYjPjgQFxTxu22tdM3GZ8f7oy3F8kZJS
zHaG4jWU1VR81Dg0zdCzdkRxksIZWrIiLeTUxM52LEFDCGQzmSmmhOJtHSmA8mz2
GwSyAtu2cDOYgFEP+ly3lY5vcC4IIFDxm4HZ7uhda4agV9NFH6cEMWnIbEaZy2Qq
S2Kx7xK2u8csmo6ujuPoApWaUd+68y5w2O/geB74PME+Lq04WPnYuGz+GaTvqYVe
Mc8SUb93JLpERU+9rml6vbn8Ub5pf9QjEJzMBUMJ5aIvBmYiOJZkMmMGda2+qyr9
dWjeTA0jszSpZZzY4FncQMJaZfBoOIJFX/a7ihHaSKI0YOC/ACHbYRlEHMRawCfX
IE40F7ODfQ3J+eQPrn2NAU4poQISUV5xULg3RYjG/4FbbT/xge+rVVdOA/pNE/e7
Pvakq7lHoiLGGXd2pgkNmP2gZceSN3n55J/qFuzcSJ9OWuoE/cWxZ0ZvtrCBWM9z
5Xu5i9Sy9bT9//6OEwOHxyWVYmpRxB+a+RPm5IvsLoUEP44FKlqg9dKkQRUIVdBz
RSYTyK9zIFbB9CRUEqPeJnZzF//DPfqZNSOO3qWTwAkMIcLAN2usuosEP6E1eDgc
d1dhWWlbFewoWNPL+gEQMabwExSiz8UwqPit/chKZPC2ewJShuqTL5M8h6EFL8tu
OkVsZgwaO3mXFbZQ11LeU7eoU5yuvTX+6Ud/l7bSg+k2UNmGZ8Q8Q4G1MMmmKnUQ
bnZmjz4lANDcmuMgMa3OQKMNTp6q3qTLgiYKJmXl1A6ijyaibtk8NnMCcHS7mfbZ
df1Z66Se0FDHPVxxMlXUDBcV3WqrMn4wBK6Oacrw1+dLl3gRVEt9awmIU0/Bnjtn
A5GYOJnZl1DzRkaZ55om+j86I3lN8XePhHbJLHu4L14wJX6F6niY5irr2fGyX6Qz
a6prFmh/5EkDElzo5lOtY5D0F1jKQYrPatIVZK3f6H1Qcu/k/6/zL5u0gWgNsfkS
+4+ETVHv6lI8ZBgIrOjIhkNefH8ZGkbSdjDBC4J9axvaaKcY7Fd709SBoVLZq0so
I3OJMAHg5Y//bbn1rq1C/2muYqRFd+/9a4+k2lPAMqHQqjFUNtiSMjWXALLD7OSg
WAm038GqgZaj876ILIl9U0aLRk1ZuPF4CD5nmRm/MyVrPa7SAww0iDZz3EC+D2W6
1B+0fi8spFDxJGryrSh3JvrX5Kn9sWwjkox9KOyW/eGi1+8kL6OLPQP7CE4SiSuC
LfsiIDF9JzcGoCXILGSVe6eY3nwfsMc8K8somNVE3q6DZPKCZxLdMswFarOINDmN
PFE+c+iS3NOjlux4tGcjgjCZ81lwxL8+hsJrtLZS1hM8wWRHEBh58wFSmUbsC64/
kpGwD9jJ5MwxePhHeYij4SyEpXCLPfPqb0Inp2gN8zQdb1WmqVERAiSyGhj/7ktd
uowlBXv4bT0RABjh34IGdlLKcpSaUWaSZv/kdwSGiC+4dul4n+0uI2ZdOjo0bvS1
c4wvC9m1heG1CpaBYFVA8KOC+U1KgYJeree1JUiINaIF4KA6pM/iS7HBKzVSNhZX
Wbzpbca4taIKMmEXa+0GlyfP/eymu4QukU7WfSo7eAvjmxSJ8iwm+EptHo/zotOK
zwCqokUJYvxzdwhfUrL9YGS0edQIvkKD04e1fmmKXgSPdWpLmW8oz8uEL3CtOAWY
plZByyxh+ZSVlV8KPEC03QEQ2IJUlnZ2YVnHTnuWA3Uhjw7aSOoyR28gWde8iGYR
VfGluSRZz9vt2YKZqam1b9JqT+e4QxiFfr3baA8rXO+9lGAPuEYDYpr+LAYho+dU
RHhmw/VnegtPAe5IYQtq5U1mCW24LHrEAoEcx0ma8/7Js7+zeXnYT9jzupz1oWLJ
rmi4oHWkMYQAXu47np+RJPQUeisHIynJl1Qe2HkqmemxrvaICdhKKtIpBCInOTXq
UMexvJnSNPC93MuSXc45ou6rs3BSe76lRiskxMrTAC7cbw3ofkM//CIOv2njieKx
saCNqaz0NDatafGoUMyp0Uc0U99nY9tiK6OAlxbmPnEb743mSgqNXk5/0ts1MftX
It7mrLBe7uHoM5K+QLdLd9/K0esekAzPapd/A6sAzp2K17gsIqpvYMyxtGv6PXv8
nElN5dpUdxguxdaB3IZzp0tkDLwfRGXfKRtZYo/RIJrxKqVQzKdn4PjpL9gHll1G
++2HC4U8J1je6dhmYeMzsYDETyHuuIFATvcmG7qOiLGO/4B81+SEF25E2fq5Lchk
Ewf9tBvrRPCErKbW3qHTC7pqTawFWlbRHpDZe/hTSPSJJIu6JKrdYgO95ZbQ0Pwj
8YWWymu4m52dmI9SfWT74AwsHyOa8uIh7ih5n54k/Y1UBBqt1wIkPt5aEKaxZBCm
lBJR3jK0/HWqREkgF2RwPNeT/K1lrFoMggBPvm0/1XIAeDMDhts9kMH1LPQNpfh2
PJpVBXvaMarOgnn4SOoYVCDF6kddj5lTY0z1GmuNRvE6xUWyvLfsBwy4i9ZOlOS+
MzYO3ynVA18/EeoRZQ0xg6t7q4uvuagm51nKSzFhA4nTwDIDtnElWgpoXGr3q9rM
DaK4M3kxOO+TBX0IMiU+pxdSIOI3tXtqeDWvTgDe7ZED5CGVfnlqao0DQ70ZShbb
ormXJEuHmUcdwf3E2mL5/XbxpSduFdv6lc3i7QQ7WgsA1syut2JyKv1+3/iXQRtN
67biRsHk/fVs2fzMobBYYxHvWC5Pq+bGWD4fGQKYk1kr5kEkkhd6jkYeus2ad9lr
4JBK7JqwHEMc3/t+CAXlltwaXCoDf1lunRxzqJDXO/OXVCpYuVidnze7TWgxFGWg
vhcBaceBTMKW8q/qBQiz72a7UyEbCxBwwjSxROF+W0yifxXpWalLIMpyMO8RlDZy
czM+TBu87kM0HsdBbcbuURR/nNRlmYbv5T9xA/Yye7w1ven0D9pr+0Xb0hiQqaUs
D1PrdhdQggrnM3dO+F0pd8y+3sIK24/9VxAMEF/OoOdqe9bpQRD9w2YTHVrA1eBa
yDOhpxKiEld3r/cZMVYaCFKWaNLifulVc7PGaa82zftFFJI+NCHzbqtA9ga/tDJD
u6Eq1A/C10v4KdhLqcNWfg76OkhmymfUE/clqYznlHy66ULADl3curlOmCC8M8Kw
7zUkWXIjqvQ70EL80PBL1oz8Z7aYgOpmS/Xk8mihGLU9/g/Bg6yX2s1gTkRko+2u
Mqcl5wVsKEMjOS3SEv8X+KdHRg41v0iOrXvxmCvDMRBgAzQ04UCrng6LmESt4wEx
Mxs+L+X+IvKE+B+RteQJ+d4sZqN54xuvMdrcUvagxG3KEcgJXTqbb2IZLzXvf6Uw
w82YwanUnddI0n37UWvhzlzQjBPfyu+0y9aRF5znKSvaklWVqtWdjllDQCOBijuq
jX+oJf7R0C3P+cbiYxdByzdZAbM21yK3CNJspe0WMbzFx0hB5LWnECdSGigElVAZ
8DDBRt3DoDwUOkMgOofm1h2pikOKlth+uSpIy+GDhM8JH9oaF3Ot/pzVt+/jCdW1
NosZLei4vVAz1ohopbge0xARhxzZ/MxdOa0d+Hw6hHGgQ+X8eSkjlgRHrIZWoaBy
hV56agUn1FSZL8abqLv6Jzi/DV7rdrrNnF+kksgcHk6W+ubjsx18YFHHEb08Op84
hznjsjUas4B+LPn+XVs3MHS9KaYueHGyVwYdEon6/gm3t0gyJ6mGuaomGf/K/L4M
M4f5LS15/mvI5SlBD2AG5C4/t968A5U46vvoJ9q6IPdKZzSPmba5B2v8OOKxp/AF
R0pU8e9jRR6Uy522YjWHs4yNPUrwCGaRB3M+2BdcabL8ynusRZGtGJoq+ntFJunD
wQdVWuwNJwpHai3mxYOe/9oQ195EyFKppEqPGqtV3QpEH2HI8XTVOFwM2noFaPBY
EBHNW1B1zavMEJ0PzZ0vIxj+z93HMPC0mOd1mHquD/6fIq7qAPniiG8ZddFsxh8c
Iq4X9fNvNKnaHr+329+MYfEJSJSIuklVt98jz3NSV9yb+RVLOA0zAFboHq5+WCfC
A1LcAG+iyXKFazuFoWemgrsEcJ7VRtsPqYmOh59dcT/2OaNVz6IH09/VZPa+JKm+
P78YW7Seympy5daIZCyAQZtvz4baMwXKKom5UkWfSTR8z//rRmsD/4TgAIDm3kON
cltAaS9hdTxNeu9YVVKOx1wPKY0H28DoegBxnfEur/tN2Z4M9Vbb6n7vV2eTCfe7
934jYQiQiHBRiYTLUlSuxKpKPC0DTsgFJ3Kb/OtAvRWaB4dyl1bQ34X9cbxI5JoH
A0NfrpvJS7/RUbR5ly+Parte/vG6DGwRYNP237OjChzUlEqthc743wIm8f/3+3AR
DH7xakYO8+Y1cvwOjWszwaibY02PIwQ+dGB2VgB/drFzo0m18nQTuGUM176Oxl3C
MCsUvLLpVHPaDxY2RLRoznrtxCPfnEBt9l1I3WNqBFIVqWhVftqcRsUaWOAG+Sf0
cJYCM4Tt7LyD6FByMgaw47kkqmjpLZP1hfRK1tulolTlUzmdo4Bc1PqTAsqmLa9w
zG4dm3Nse9Fu3MCjr5dPwSMHirQnjIrt8iwLAXoEBP7siICOxzc8NUcUMUtF/f0W
WLo0UWgjR9hsQvASSz6nIoOcbCMMFLTW27sUGE94145IAWZ+3QUMMMwtiY1+q2BK
7auJf5wiDOLkmAMaQ5V0XyBAmXxRJ+vZBwipBVZK2kl2bG7pI+VsqvWPVopSoGPq
dOsw+t6nwUDNDqlKfsgTQOr9B7kG4/6g7pcSuXWJwro+jsY73+UALuOwfy7U7kOM
08Ynf9je9SpL6uqP0Dw9lRhzj2KodH4/YQ8Uk0+0wazrPSovXSii/VREF8MMO5+j
DctH+hINkWVYkElIxaQgtm+V8/4rHk5po7tkQoVclQtH9CMDgUmepRRQzq3YOxs8
EhbYyDtERi6bGt38xToqp1TN/KHOq08nDogf35EBXb5x7x/p29zEd/m24SM2zGor
nhkDcluDrRTc1Ie6spbNkWhVxOFxwxqrbTuNh6ncK+ZEdoq0ac2elqTlP5PfsoWa
bRlREqFU9Jo84Gwpxn8e0sK51jzCZFmveBU13KRXn4PcLlfcyLuBS9p+puArSxQh
dyKKukQglJNPJOxIw27cDjFEd5ShDhUMEqVSLCFfYYbbBQr/s29ALRYHll72t5h/
FFPf44QNhjFFaQ+8QQn2qwhUYAnl2M+jRT2wINl6RFLl8c0p50XqvTRL3M0buwta
u4a/anqf3m9xgf+1ZlSqE3cwT1dwP/MiULJhZawkT95kN8ZH6ZePeXCbpEjjo3r6
iXLHDJENjQJFHLCp7sOvvfVPdreCdV6yJ8iK6th8FUyHToLZTeHkbdORN+80Nxdb
fUftA7UL+1B/DlrhjOH18jy7zfaYxTMOv08fVigW3ff+IcSp+fAIhof2yLfXlnbJ
x/4ZntQ5bTeaJI94lJSyDlgx1b7y5VrTSTxuM3oDFGCHJPunD/MEZOq/ijukHHM+
lf/MsnaeNC24I+pw0ZC5XPIcnj5H4lQpgxo8ku+pS+68YAkpWsuuZ73SzAWOIfWZ
4a6dk1AKclMb5lhkrekdf3MmA0OnQ8T+QIhVeOyoqTZx9Jv01XsvCs4l/D2cdRXO
p+VtBGgT9oZfc+1bEyXnugSerX8xS9BjTwLaqz4UJK1UQPnZ+4cRZj9U8aeA3epX
o4M+8da8YueW/8hZafGyC126DFJxllOxTUFThd/XNAGMePphqnV6M6LfOwLq1aNl
QgmxN5OPojbjJ9lDi0t7+Bs5RwZXce87XczXSp7C6Sh1v+Bukz6zsFnqruVQoPMA
dpAO4FTrqEGJVYya/lCpXD/J6JrjhVhU6rhAdgB7B1XUt5drJ+aPkVX6M8rE9r3G
G2+OaBLXpIZOrC88dRMabIBL9RvmBXlyKAYDzLo/wrIvt6HrlpZ8vsZm+OxW+LEL
TFC54AwIp/P2CmvBwPFR4PY5r71fU5xbtv98Ufi/5iCox1QjdqlajHxrHfqXZoVG
QKzYM+rwBgVRouvnU3/rIv0E/8MwmPKwh36TBGjowna5jD4DWHIalCd5MSRCwKA9
0dE6vyMjiWOfTDKmZQhse/v9D95VEmFjCyOjgUY/mMuRLUDoSIjvxAWrLVTRO8+U
ehykb94K8EQgjwZPUTJkH1i9kyJrvp3tGRyNmVbWt5C/RO42uSv5xrJyU+Lak5Y2
f8/lfv2Hsa+RAdUvKaBdiZSIkRD7kHOrff7O8k6o0PYfogWi+VPenMcKz+hTSvcb
xRICu6CnZyJBX9CE2m9vzMNM23dkK8YkabeeMZxAxE/47IhutKbBqlMON2gGBGbd
c952e/dupdRYBFgI7+1Hrw7+jfmlbKcY9MkSSgn+BA+NJk2ju97gIpYdfTuOPar1
JBegymAqtmQU7n2wmcmmGg+t7G+63MZD+37wets5mkR98ZlbCitKkG7TN4xFO2kT
LPIET7AUhvyKL5cCw/v+6wslf3RBvGEjaOtDZwaQX3GpEcJ3DI/k/vScRDcmB7x7
q6ZoV58AIzJeoUUcwTFObMrAdab0nJapYMBIWYCh/5VhctUnhKwCFGglgvJpoBC2
WGmaEUdM0o0Y6enpt50t+pBEkjZEFISauwWIFtu3TQRW9jG4hcb455PGHpMtLDgQ
PZRcYyIyw5/pSj1fmXiXgo0LqEAA5O9xUyIIkH9iZM0qxll/hRG258OGfw1DxKcQ
zvyuRCkSipmCdPz9vmattyG4w2tl79n0rhwq2O8x2s1BzlUfvNLQebGyv20+Dptk
qMbsjke0jGSsoCfHsdJuoNnMF0BDkL9eWuxnjZNrM+zQonlovoyv4AoGSB805xyx
bnLd6Fs9LwLlHgNi0iJNa7fVp7d2fsujTp6/1U4J5EZQke4SPAYnA54LuyX1QmpF
pPKgP0y51seZqCeblvScRvn3jvIHtSssDbd2gkNliA/b+mDEjkW5wCWVxORsA1yn
WvPCDHcAGisKaL67lRT+jEzcmk84sIJHEztPzBa8+PtCooilpxzC0NgczUqag5lx
cIOcGtv8z9QoP6e9wjbi77ELh/FlxY/AdtYP7rYppZ7sLzaBGiAbcdBfMQadXWJa
yOrJerIe6CDCXZ040NfJDNPlbnzVNtGOKwyIJDtAnPeL9+YmLY8c2He+mgnng5GH
FshZxRBua7lFvuh14GMRT7CZset3iDf1rEYXtFNdbPZnFUEOj2R3bwQR+Qp1Dx+5
LLUECZa+Hr3tHxfbUWGpkKY5kckM/r441TL1cxKKovyjO5iM9Hx9q7DoNiRHh6UZ
F+JrOdbKau1f3jR4M2F+iV58vpCZQLPvcQg3ZlVy22WpMZ1qCKUQEtdgi+VKGCjv
vMfMA/Bi8isGXS+anJkAeVCFmicnIhJMth0wWVLF9XS8M8hvU1sIAAqbCcraan1L
Oe0ReLoGSjCT2Z7gqGD0uJX3UE/peiEpNSGvGh7aDMkLMV/0ylcY/mRoDQl0gfLi
9HaepJhmtnazuAswqtLmkoOBmK2xP2Qewg7vsZ1vQhAjyq3n+wCeEGtdzU5wJ9LJ
JpWd9uJKeyVnJCYrjVuQD5F6nyYxmw1vJaR3/WlIlPffrB0OGm2IqFxsMByDg5+S
fT80y547gTr0Bw1fDnisA9FWFdoYKbuFvLbti55ANHCn0taNx7fAebdYxbt8HanM
WfXBXLRjWdLntA8nsssKMYKNQE/acr+0SBPSAlzQ8GcfI22ZnLuAWp2TOXYwx06o
nBJI96kGqZyW6B+6qhqbvyhsD874dyY8ylk8trH65daGNMQsl4fcfsf/vdxq5oZK
8jZQtO3YDbvfNP2S3MlD84Hr/pvLdYS2q9Fc0JcfZnKjLwXXN/ygRsAny+fOTV77
dcwxUZbVNRNXTV8iCNQldeaGnEfU3VDIGoQE1E7TPuG2jm50wZKGkYxjCyzBFUax
by3HVxMSHe33yw56mqk1XmAmRXjvlbE/FRSUl9iyythPuuXvrDnB2lXBA9AGpwyb
ve9qh8VeATUd9BnfYS1J5TI8vvkzS0YKepp0hM4UBivGPPlStAybMPb+OCF9FB+n
ChSVZGI912scep75C0T+GZQESzOuGbsYsv/rlihCmClFPyy7LsQNciUPWpprscHP
4qLtNQ5sna+Tu2Q5bzm+vew942gEx86p67EYCXnE43QiXpg1kOyP4xesha8rhuCH
Q2EJBsftvQtXbBkUmY++stBn2k5Yl7PWUfjnSauZo11gOaxDWrTZdDgSb+YRnpEh
mr3k7+D/mfThVOrSPwM+uCRA4ArEULC7T4ZzglxaXbOUaiFhAeGSJSQrMVBkthTC
1iTRiwKJLCLfqxiGWy5RIYnICWbAYJNokj2VXlTTBVefEN2TwTG68IalOPWTZR2q
IJfFzMcfF15TZrpq/oy0OsTnTT0mcFyhPRF9wixwawb2MhFvdR8rcaoQe32AJe19
Jmw9i8BFyt312XhEJJ8Ox1Aoo2TmJgP16Nbi7DCKWgR2HJvlNAq1CTm5EIOpocCQ
U6Q5QbamE7JkFAH64dqW0CJcyZzJ+uaOI5A2BS8jm9EnK3cy4yhqH4kW/IA3zfQB
GjrA+P1Mlt0MDSQLU5TfivX2+pW5HcQmc+ZOwuOVzKdPfFLzfRPzN3PSm8vef9ZS
BbaOl3OTnHnJXvQnb9SK9935iZ5+wjFavH2vi0qEpZqur/nFpMN/Ue5S5E++b/mA
vPM0VhdychK3I3nTyn0mji1E1uEU9+tb4hbM3NiDVXkvntfr/0Psklwyw+EqL+/I
ICbyX0G8cU/JeA/5pLCKbtcXqWv89tAE0oBAdB1Oy2kbCcuOfw1DaS85TUyfqOeY
hswFkDMpa8fafZ76wujRDN7SU/IS8h7YZDA7QdYgHrMrn8io8uPiu9h8qlAytaUu
P/YwFTSaMuEQnxQti7VMRRx4bZPlp0pM8AXW2JaDoKsJUWyt+HJpfQZx036giYmS
NgORtgAQn6SIddbsLQgxKbicQOXBnP5nlna6JDH+aFl3rm844QI64k0DcC7dftsQ
P/mxlnHj3ZEt7BKScX7v+IR3cGsWUkD9h6e/vdu/Aun0f5gRCLPUf9PT+LE9+VSS
dpABwxkU3OjKzaVx6CNz1uvwXIBELnxvHA6jRJHegXNuIQbXuWgxGcEIQefqmkBP
v4nMeM2NGUTZp4e+W7uxf8LShNQ6IKFEVJ8ltUWzotblciw69xZVZsaUJZGCS6Wt
WiwPlpUxPAxtLvSItJsB9At7lemlrUpS9Ew+fTJs58CBDgPDGDntq5RPaTfCIuCw
3vJ6FKP6gj0gJQ/BA94HexFckNRGBR49vRS/2+fTDsgDsfu4XyEdLzIMbVxibli7
+tWj3e4mDm2KlBf7NoeELxd8dOA3LjvWqOcCyf+4xp7zcb/aDjC1qvreruXa3w2x
hnue+5wtfKUnfTYUOIgSDsIv4UXfQpvcoYpUYnp2YOg1fIxC/kZM9WNRCtM7NIbo
Ocfx+eE1JLCGwwycYY8GJ41AJBhiv75bCc6wiq85g4bgww/KLAAo+j4KEGxDI348
QS7orkyc5wYhmUwSQmOoDkxFmQcNjnLXH3u+UtChYXdxeXXC2ps8o+YmciJ8AM7r
CZJGTxIGSvqvDSO12QyWBMi0fh/uYKrYIWSam+YIcCEli8epm6jyhdCy5RqDl5w9
fb8umPL5PBGUr4vebHBLEoiMJ1tUX0VynAnbqorQx6MpydQ+m8grNauXjJl0t5HE
4c52rL8RAufl7m1fDEElbTI3TItrfmGfdCT+rHQf4YYMG5NuglLZOgIWWBTD43tU
Y9SjnGXcbAgqt4cauPIhIKpTJuPexBZZVL2YVvGAT19XHJSywID0InJldkewd2uP
Ce7vxhEmpNFprKsXKdX3lDp/s+KgLvrKFpV7mYYcl4eeUniT3isO06JzVFrjScVE
NAlO4rTKfJrNxVn60BEvZq6XZ9MAnoZuEE7CKxR3TfJ+bu7HEbc/mhR+fMNyZ9bU
NrY+QTHXeWRmv6X6Teie8lmZNCA1F/N3Ij9IkmIDI9Rs7l7xDL2uUp4+3ls0SkRj
99HwmhDlhcIdK4Lx2bnnlwblOPUzZ1iOI4AiHliIr/48SNblSTTvki9xkMrhsrnv
x918mvOpxH+egM5PVEza48cJEGJKTjvp3E+7tZA5Id/gdq2JVmjeUtDRYPJRok+P
0roExbfyhdtjQJ4tIhvXrU1yYFbzzwcvbBQEv185LrON/PSbzbRuwm63GTq/SEFP
OatPjNktG/Ogwh6N+vwOiRynUbNqAezd4WV8tVVdUDOHR+GBlZy1hSO2WPf9xzk9
sgL3pDTA9x5gENQwNfpgxy3LWMosKwSO0RVqxJv0G7O3iPEoU6dZ4juaimCbufkB
/IJvAKH99lMwnFU9LCgN+3EVa7RgxHHIU+DvfscTULIiCUppt3sGk3jzksGcijxF
PV41a5izYtne3oScV3+uvSGKwgcDXz7C9VJ+nBTvH51GHpEz0LzH/5ohohC8IG+A
0/zkSgU+VK+gMlafhk+8KWqnBlV+AttN9UCcARSLI3q/NGa08rMLGrat6a8f3qLX
vJR17xFJNifSxsoNB9lzn+EMPl6nkqKGBC3aDttpaZDJ6cFmZJXN6BgH2W4ASKjC
/ln3MNf7uasZwcAtcLjE1MEngUgXNNzzbJpARp6g7CYcKkrPm6TkUPS+lHnFLgoR
jyg4p2MIpbkaKIMtyCw0bnKZ0eFDkrrn5EkonZsshSHuf5oCr0+zvnkYC9/gDS75
s4IgouJ76kdchXBcyTxd9nfiSAsIQgNFFZFg42gtdHROGCZos4Du74ZdzMxT7iHU
7ItlCqEQoewdes7bT5PP6hFY6zkt9FGtPBodzTYtBm+hM411BkrJ2fnXany02Kjj
2vrTpRIuWPvCR7QTjjaL4JLPvgSn4WjZvBScWt3n5l4Viq3A0NVLgHhXXTIOQF8W
tBnZI2zO9hBEX9pXcx0lR/MgRNTfP81zfwSb/hzmD7bNEjTAvzx6Bo0NOKpmv61B
jMT7vg40e9inouHwhJFcA4txFaEzSETj0yebHfFnYEsGcH+v4HqT0HqJpQY7/30i
0AS1h+0H4XrIDp4SyP6qBPr5pf9UTQYXeM35rCq4WRo7rnH4S6Wb3eQOc+q52VaY
Mf1uMTQDcm3s2G5S+tc3xtSLb8+bW3dOt2DjQu+ro4Uv13n1kpNB/by7r4NPbdeR
v2kBlPevkzobkferDWoPeoeVMccT+2En7Vn1tFtvv7nfgM0ieZa/6Cc6iuzuP9i7
LjvJJEn5glsONOKvq4pJt0YBAhh5TkO8zjzSsFarnKmPYnlaR+tq7Ro3i4nVF9PE
n1P5ApaA3Cf4NMQcYoaeJPQFjX0fK0O8gblFleD8sZr0wqBX/3dyRn5wRtYqaeXO
J6sOIhX3xJmp55OTbtCKlJVEkdRtxTZmWcyfEVqh2Ps7eijc19bLxb7gbTjPLZZQ
qYzoplIj2FAipUwqgMbw50Cb+X4PuFLoFYZj2giN9/H9LoJeaXN6u2cmHtt/nGls
sdtedLew0Q4vV5VamPkQ2tebOI9UyFBi+hjxHM1S6yb/iWqPleZAv3Ro0wQNq6wD
57+iS1eQ4+soIRAujfo5ZDaU5hkxEvTDX4nrA6o3jYEtsXYNbk1c5GIbEmFB/mO6
PPcM+mDx0EsGtiVLPh9z5OE7maIQv8C4EPYWucBoyQiuKPJEYtjG5q6AFvadAw03
E6328dVdJTOXFVM8wi9WOdTiPuoxCXsXVvUvBZSnU+RFiJ33h5heDJiSqG5oCkwn
Pkxu23Po+yKmqVLzYZT7tUtyBMaYzy0k5s+GPUTf+2VpDx2WXAJyMwLnB0kJbnOL
Y4fHMZCZMIE9NKKXq3k8Rxvkd3IyYmlFDZx4N5qaXjZIYAYuARh8HCWNht08pkS3
Lh3iPqZ4B3mA6IRlzk6OcSFWhIuNZC3Ix0JnT58pjv15gJ2r+qRY3dUo8wRdM7GM
r2r7ULtN0hhazrrjl0gXwGvhm+22vMn5ilZ5JlkvIQBeutGS+XUKu7G8aP1iRwCI
3hP/kc8dgNcMq/q9ugLCCpHIsgiLRBG5iqZa+88UGs6fhx/MQJJ2wzXDEXffB4rq
RIaygprhqQEl1tb3xzlbrw35rhO+pPljBjpxxGF9WmODiAzHxZP3JKbjKQfdRm3X
q2lyIX58win8VXojzGQ87O/VSbq2Qb2U6t3WyALQcBUq2pakmYfIhkxFSTZBzU/X
ZySO8roGRkR0FOPIS6yav5tkhzn3po5tDlweMCbmc5CTEvK1rkV4bU08SqRTu5lF
rszBaxLNQb4Y3yQKvcHlscXiZ1mRplGZj4CuJj26mv0+81QSG6Blj+oX0yNzgdEP
XYDyeFZzrjP7Q7DodRlv/zsqqTXYEh+90eNVuWXfLyRo2cZBHH6K34uyYu5I6tu+
J3myxYZY67v2m054J48EYzXGFR3kbeIrEYSR9Edy2y/ZDZCjAotnT/e2U9rr03qd
ehBAMPfrxdet9UzQ3yKfSyfSabMWG93CozP7bpJ6hpw628MD3bSTQwragDIV1iEs
6ZcW6BC1rOpkAMwYHoMdS89mtsjMETFUNzCt/v4Fc7VYLsrSyBM2V9TOZmxvgU6z
I2jJhr5yxAEd19iKeP+WgMXHNZw7T7ss19hyONtWQXhb6KBrAkUqDV9jrRBC14j4
R3lFkj0y1UyeBNEGAVFcmmHLHgbVal2r3BFbgkwIrCehagS6H/pt/NMhC5pkOWcP
874MB2FMuvMLK5QxEpWhzH+FqOFQ9i/OAIOCDuEf7QZRVPtQM+GXyajZndDNLIPC
9270ixqBcjXMQFvXUSZgn7Nm1dXatM7sHeW9l+LrgFckXWTOm/7BeO1anNkj213v
BXPc1+aT/5L2qaRvJdC8wWR1koSM/pVGGq5cjTrQmuw3ZDXj7axReqcIIuWmstRY
Il/u8UV+S1VMsynF/gKSu2h6IEg4CZwb1ON1IFhVpeIy8DD0/ihs6nGmQp6TmBTJ
aZ2pojzFKi5+/SonJG4IPIjgnB1HAjPXoM5yInv375OKpm4oNh+787R2SeHGQUZo
za8FtuwXG4npL9I3tGwanlGdz2JtZy5xzn863yo4bjrnZMm1foHK6LqLrJw64RlK
5FcjEqWBjsPi8V2eLGk+DL6GxuARAFQo1FV/vPqKMjr9gdevqBOJAUZ4+jzKQO6z
PerAxwpNKYswFQNno+2EMFODH/1UkWdqrWu6QxeNv7UKSYGQfZGpZ4/maFZxKnjf
amaVtNNzCW5T9NO0mpe5ulX1Jm+H4BFWFLYu1sbiCVSKWDwg0MMmA1u/QWJzw/iV
EmVWxYBGvoJxcXiMY+1+mUnfdRh0jhxpTHuSu5nlETTf6rjzuRR5RheD5DtVVwPa
SJFFZjq0Ws11Hp0BZv4C+Z/PQbn0zXB2mYU7PlYJ1aZT6t7CW1xY25umYO/bUUaE
Dn1Q83ggmVia/TLT4Yp/oSXk6S+SP1aeV8b6yOw9gr3AuGin0AAf0CoUAVLZTekf
akt71y/emB05v+5b7mOiQm5PfWFHZ1Om+GmoX0gszMbZqhrHXAOM3SuEcD6tuI/t
DObY42LhyvVGH0EW6fmO7kQA8eKNYBkedGnYlTfendD8GFjXvx/McJ4pEdNAtqaX
zh9eLVVuaSDcvleh8WURJ/gXagMPztLo9kADRM8fnJCjO8Bd1PlNgN4LaSs7gINE
ffi5b7sUUQBFquYvfPorlNgkh3AsrTS84+W9re7wDuh1qOTxlKffj70TZMtuyN9V
qBK3hmsHf2vWk8jNjYfK/K2NAvdCk4rpMHRavZ6XlB1jyep5wwgite1yfwSTaa88
ZzX8WqIII5lx8pE2XXHmHuAUpk4IlasVUK7TrlhYUTnr3s9q7O9mIcQhiTVKfLhr
0hE7sBzgf6pQpeLsYHU4UlamIxYHz88sLLmYIOXybuGOETaI+4XVaGBNWi73fdWs
3JExv+K3rpL2Xh9PTmyyoKggWpcPTz0ddK3+EyBod1wMnxuwAQcCMtTxMf0SQtlh
3a8xBGeBv7zhFyPUafzvR6FPkcy4lEkUpCcHSnEcGYMooF4vo6oUKWfvsdbSeTE2
nQI6+sN2/erCBNpybTLsOu91/O1n2tGj8QAzkYYIxJWPogS2taWvDIivmSsjeMhU
9fEHq+TYmd9BZBCyJzhj1GdXuogKFQlgHwlpm0JaidRg5q1sJviQbE/sG9KHXgRr
Olpplg22YrQNG3WWHLyBe5jvdPiJ/ulrPueKRRztMJcJtWAfz1GUUor/UjP24eex
W5fjGIU2Cba1wdNDJ6j4ErQg54Ke9CIuEoqZMwEpVJ8ysZe1e2VKhQVEzDuT8uR/
Se5VVyyIG/DGYj/89kV7/V5v1XLFHE5SrBT3EWwBWFg3VKbDaR1iyA8Q8peCrH3E
sEB+lOZu3Ah4310Gec0L4Sm1tNxGrnBiPi2B2Ha80vUSQ9YMw0mXywaT28JbQKw7
S/UDnlLRJCBSLPuXcfUiU7T6kppVKPbzpwvjcLFL5A89KP7ohSdlWhjIrYtK/DHE
8iRsf2buVE5jpcTrwwBq0n1WcmVRsKGUTjDc8YBLmSEHHtfKyr1WhMY1FBXPQP30
eLCmMLEZJ7U3TtfB16+T4dMHWS+CG4KztUSRTZ5hZEQsdudx+RmmyAcM6jt085ap
/EK3DBmo9z6mAXa2sX+TcQGYmQTVReLrImI5noVX1abqm8dgxC11b9ruPj6kWy4o
F3yY+MZdFiLtcdc/PXIgk/0687aEyXDLvlvAU6G6QkLjponmD3yikf+t1F9VoSYF
un5mDRKboHVAfL3C9iWi2KdEd0H2jU4Rddya+S5hj2pZm/fi5fZ5hacwOtBYwaoj
AXv4Pr+CfHcSmdjdQV9OBP4v0KoXe+d9be5CClwWG6bSy9c1qnqwIV2MOv5TWFZW
04+vRvOHnMyQOaGf2RBb1SL6HDBLItjfUqtaqTHrwLCHZBYW7uzad3m/7mPwPJu+
Hv7tAfJJi4HZT8LDPYQxDR6th1AOaWAdl4y9lZUkYkwTvWFjtnkSb1SuhB9jG6ml
f84mInrMcxatny9LxWcXXOmPQgkNRLbfBfTtbMRyOsY97zjTjSXQixrrIvHhTnlH
9/pWG/Q6id0F6gqxtJ1SW4t4Gr9vDCGWJpRu/oEPY/Ah13WXeZI6O4g5i92jXDat
47Yq61oMXYECZLOtfA4ITES/CKrpLuSCk/2Q2cTTzRhGawNf/bKiRwkN6WX3kySm
ZNmlfBm8QnHUTVfKYqcGUz2mYjrp/ipYRSbqAAPrlO2XZ8qu3karpRnskb4ISdsf
yEGftlO+MKtjWxRCiDR9ReFHVVjILxPBorpI3Qirt2zQGxaJBirnYqFRlpjdNH5g
YWKUtjeFnqsVPapck98xneScMRp+5/uWQivC8grTztzCwgoT+43RteUEV7GOagWc
PYcxVWehqcCGs5dhYjC6MQdB0hL7q2LMv3o1JSijqj4GzdHT7+D2V4icDMSAtiva
wJ13n+P9U9RNw+cCRb2S636gL7dva4DYLtb+XS1XA/LfcnOthM2D7DMlLhZafrbo
2+mSi1gJhuBnlRiDK/Yj8/zzAv1l1VeqeuaTzLl1NPjE1GUWVHjvr+2Y7QycyA2N
XAYtI8llUzGQkK2swh4LEHkiq9AV1g4eHakhxC8liTf87tH3VRae52KtX0BZiMfe
aOfOjP/Ze8fjfdqA8wM7eMWn5FTZJsp+DfTc1lQVSxiqjdB/wGLIbyPSbj5+3Lx3
39427EUF22I6RsRvzsOFwas4F0807KaX0DDk104yzOCTTXTLzKlPVu/a0sLRKh/P
g0/Zna9fok0KUBaGiGxosQ6wwlUijM+3l+rZ9t8SIWTx6DyMSfhTiFo226XtKOBt
kVhMSUs21KWa9UrVkyvFrqJtrc/wwe8uqkQvyZc8s/G8xvylKtWTeeaL7rfAihXy
4Q9so5EDBssVPJZdLj1e+GiZWbQM2JTpfbVPbeTDHOYxE12n0B2FXnvBYiHCKbU/
l2a7mlPOpJFyIWzvebvUASFZZQKK8fEbMG3s0NY+PEYduHp6bxoYYkVC9qVZ7fmu
fRJKmZjeVqq0GS5orvQnclDtrGIOMUO3hfOY+CEChM+R/+FDKCrdi6Y6eU1b0h9D
6+Sg1hiwsSDpconEHHdfSW9LaEgytPGUAXBMZnvYHJnhql3GR4fN4pl5eJAtSe3s
oDwIdM1cA79QoTKQNvIv3NnuyIkIJUEYwjGQ7022pGJlwvHgcgcHRIe9SA7Fp2f8
DZ9DTvb3UrQl6p085UnWhiV5vBzFHCVivFBngEUFDRe8W6316kzjX9TQH1fJ/f20
84OZENs/pFqPW6APnsHGbq3ccDNe/syuTsvbb9x0cKA6QHV/xzscXtuLmsKPFUxW
N7njixptzQy/s7r459A/Z1LwDvNehgw7eVpONqlIhx9skOSWbXZeEgNwBsxpo8ky
WOU2EL2oZdY6UIjUqV3M87ocGKpUZ10UDptYHEt4j5BiRwE6SIPd/9jZU6U39LJH
/XmcucL8h7Sm56eACuMsf+xe73niKyjNdWKRdJ9cqrTealBvF0kS08DIThpWChNM
Kg72Mjpban6zObecZS2n2HkO+Hmqi8kR/hCPVTPh/dEv3crXCEOntu7hbpjwoIJI
LL8IVDyiXt0rutq8H0FKIHpV52ptpoKGsLQV2ZiyuF2Y9CSHxtkp6asuhk4EQVlq
dGnRk1UxHJGm6LMpI4H8AdV6VGGM3dAuQlfTFY/HElQd9UHoGud7GkUb+NYr681u
Afwyyc2ihKwlNlRyDI1PT0jW8G9kkAEGXv+crwqkDZ+H4vWISzibZSHheWi9WOEV
YRImVR2jTzoVTlio2OPch/Q+vURbRx/sx2uVAYoQNBgar3oUizsGUx1J+CIllyRr
9u22jpli9vhXcgX8glMYBX79LFOqEGJ/P1ognq85OymPKq3FNsM9gA171xhJasyR
ZyIoq8d/RUiHY5+zpMDCg2l0iQpJP5dhvZLdElbPaAC/k3jZ0a+qOZuD/D/ibws8
YyW4pSufi7wEu36YwLXhFUz/gSnNPSMm3+JfL8EZpQw2O0e28lxiW2CotWt+Nsri
HiDwpuWBvld+wd3SZv+0kMnVpSK8ynubKCtCEsfkDDsqVfofU8j1OjC6QqcDStmF
76V1ZFTbxEIPzqvTlmQANegRzVZNMZWmUBSVXB4z1oLNbnyrN+UW1TYzy3rFSBWB
DJmKEN6pt89aLnrP2aaZ+psOCylJWJ/w/xgrJ/nUV4nu+2FUePvweJ8pJtVELFmq
6caNTSdzVtBzgpImMA54UrwOlKKt/3YD/ok+kg7LcrwSGREdN2/CtBWznVUS1iuI
DxAtdo9HHMwjF2OJEfDKH7aGRkPpSZ4LJLjf3AU+ksEPt4DC8qmhEvqOT3g4amNx
8twUVz8DtmNpXDlfT6xxwi/sg800T2SzHLfEnV3ZlPcDdNN9fUmeJkTBlcgeh2h9
ZNNAWXb8wZFv2cPl3CwaQxwTn60QWte9QVxnO6kFWni3lQFoBBbQWMtSC2gQF7zZ
QTa2AVlTi5zm+Nx19Q/OXL8Hi4u87l5z/C+7OcfFZK7P5vyPn3U6qLd2j7IJ1VVr
TBEjQxat4xLo+C1M0OMm7I8CgESPet/QFY/pixcufCYqfdLRAWHs6ObHGS0Wpd2H
PeE6WdnpBFLSo8ai455BIPHNmEIaiLupqctpiajQQcr/hWj1bOw8pEHQ64MSC3BX
49sgsW5Z+Ruc8CMhe7v5spzUfgwGSjnarUiduKb6ADQ3k4Iufe2eJcQbpQOlrniP
gwG61A6DHHlI2BR4EDz6hHBEwP64/KAQDP+B6fw41RTCzIFnGIjMpeQ5xXSPom7P
MrJ4K9lxtIcIVEt+vZh9/W46CQ2rhkCTG2M80WhlrC1O4TokKKERLSFj8QQnzNnd
nuRmrNHAPXpE7Jni9zL96a3JHKOdUt54/kf2RN4qCmBoKY7OmPTWSd/IflV/VHpT
sB5v09lymfbM6gt09e9X4qp/2Aub8I2g5muV0o9VJ7dqX9EeMGJ7PJz2TUSq9J0G
v+6WzFNAK9ao5Qks2re0i6Wpc4++UuPwz+kL9aZak4h28tjIS478K4iRboaCRsP1
WIfY8rocx66mTfSHsaSSv8ENZaTHr43ZU8XyePQej2tOdcyJfsVyLn8ytzSw6fFK
VIfq1sybViJ6uSaZGmalwQ9ZgMa+OFLAjxYfdf1DAW0f8GV5Bqb+o6J8yTxm2Sc5
wEzqRtAXVzwE+uI/4SI8oMLvkBoyZK6rcitflYEDzcpGl+vS9aHgGUSyrm9PPWgH
ku0XSxWVclHZff0jK+LZtlJjHEpYFl9pj3XIycEj94j+gIaxTn+FH8df36LiDwdB
TkynpnYIvh3eLkocUROTJWH0BYFRgh5qi/54vOEpvsuGgVr68SFso6YyHSLPzYEA
GgjdGyPQflYVoX4W7EPkF/ox7onz9F254Ft2D5Ue+Xk/zpknhWuilxvNUeabeaqn
u581u5IMXfwKZnHofA8xbLhud7pW6tXbPp9++hbsov07eG8UpYACmr6VFROWlN6U
rY9cWzoTZgjvJ2qBF0hyFz4DiDSihZ/MbrPVFkUeSkbRRJtvCeHTZHQL+0/TGSqZ
ZIlmbxpx0R4cix1nO9Zl7x5qNRxRy0+La13OZiewO6+wk7iQzsr1NiUlHmKwZ806
5BsWo3WvoXDOLxFO6rkz8x12hyD+Kvh/gAkUIMLosgVm2ORcw7orqR/Lwqus9EjK
4d7JgKBF2PTSrzNhh3/F8qrcjCI0068Q5IZd6ueQ9yP5L8uAFPuR2BQHGMV9BmXB
4j3ZMdE2bcFrk+guMjYI3vz0V+QGHlrsNeQdKutJmN7/sW/iMhTPJH9F50kxfghX
QoL20/ZscorFVgmp8mXNeysdOpfAeAWnCSCXq/WCTsX8v80P5KSN6EWVZwSIHpVa
O/15DzI1nXwbWpXMFvSCYV8oImFDcXSkAZfv3s515ZUaLFVFtlYByfJK6YmIdk5l
E09J/eiAlWYCWQmbuvus/dURiD5+TiYf3bZ81HN/BozVBk569XXwT4GmYuIllOR7
d36f/XdI0CLoeTakQW0Rvc1aXrHC9jos+3msaUM3bTdlPnh855CSHRn28wT7TZeu
L4w7XuSPeAYJ61MN7ZoVwUr8PCuF4bct65Q5GFvquJy56QpjX/YhMTfJUS4nfJX+
D6yHBxgdvcL5TADBa+ZQTS5jCWWDipGzm1jCcGMwKrMIHiVbowEGxhdfEWDnKgIm
TsIMle4n2DsDpqvBmbTmL8pJjUXgw7HdcHL3Jtob/sK9FQi/oc/3og2XBUK/QYcx
4Cl85X+tLguAyZtqsmRcZYvSZP5B6Zu2chDHTQcVLn6VWFgc6kgApeT1fJmS+i6w
rE9qg0YR8B8RDHvc5AMI4ZZJjCElYJgDRYZcJgF8w0FgErM4EUHdeZvkgx0wDPCq
HUsPKl+A8QGMCg209tn3GM0TYwAB3c6qddLRBzFjoVI+yyS6mZDEInJla69tRx78
sqDtgdCm0DQesP/eDMiCKH7uiS2NMhvV8zi4ERf7A5eLpKhVKOgAWybzPyEQPRJv
ju1AZ4OSzu/Rm4ickF8qJMXLo//2YTRZmDcYGWye199BjEVqZS8F9BL85d9OziTE
mlFxtVxDkfX3LKUlgiEkjKu6dcUeqDFMDmmyUHFTUpu0G5zw9k1t7gK3uYEYNSbn
7Xk5GBurA34x0tRfQEKAA6e3FaF0ICuVRFIEM+7obHvLc7Kw7/3n6yT9uIZKn/7U
Eq4+LmDjhqF/k/3VScaQyIzKRSHfPWeiGSjT/Bdd9LwBgz3CpiVf2ZYk6N3/mXIk
BS+pC1wCvDfvvMXeUM/4HgiFf/IjP6KWVM6Q8BdxtgZ0+XmRIQD8TqtP4cXXe1ih
W1ncp60GVeO6LxRJbCvRPmb54xwfbn5jDuQhYClL4DNvqpj69ot6B2fYP0TUuBMJ
SqD6ojwUDwP4F1kT7iPfAfid0ri/iyoBQkxPBMatEgJAE8maVCTFWbhhU2r+pnrl
aKqXZFdyACaTUicwsd2MDew303r5Q4bBx7hwfLfP/zs9Q8nIdlf4fAkZ9UsN7Hse
ufKTlqI8Ql11sssZgIutmSd7RnovGRO5QH/qxKD3ZOytxs768rJFCiV+arW/gTqX
+2PvrydIcRKxOp20Y1+6Oae03+fmPEOWADyOx4jTQrcMXK0unMRVVhEggwexUS7N
ohLHdhJVzUymWmPTbUveK5nbcjZOU4HNJGHdtUPe8RDWf9ogZkzDshV9jtYLMt7k
1CMHwf52T75X8HOIyocLBt1zdIekrfAcB1m3klIEBCkB8pzsbU1L2bg3I5d7cno+
o5RxDt9jmFTyt6DuAjLm9rFf3S6gHeth1TTNNYcsm/96YA8476w9pSRtfNsvrXNC
rC2sHqC1oFtTZJ21NRBuENmbqNkaqJoMDbE0YXDL8lZRCbs8IRCbH5Ghj98IEHlQ
voACsW4sHBI2NbFqMhEuHRy1fmGDFH8Opg5PlLnbK7vnvFAPke7BeL+JUfCSnXxe
DWuzdkZclzsL88HQf3EIZ+B05Vg7HCzqjIuqnQoZ2881Z9UQzDe0S1y1DIL7CSLc
TPOOKuORUg4l3CJcAxfWBVikaeHvFoBYJ6ipP7CAH81qHMCk54LK+2QWHh7AuYJB
yfxMP7wTdDx/YPXl2na7L6nYopwKUemqm6maHigo+0d1Q9KC5FW+3Sn0nSRT/Pwf
BSoeAldQdJ4E/tGu1SljOuNjaDik8Dm9Tv3phgpjqid10uILHWjGDMyWCM9GY+Km
QPIObvfDSosnTO32RvSiKtwiduiaBCACtgMagCzsrMw92Y/3zwWmzjlWplbdqWqS
h6ouDOFUDPvdc6S442Sazu/5gnWyvmsFG5z8RY8nphPLUNQ0Nyf6isqcvbmNNo2m
QBvV50l2mx/R9wGo4GN8vRBCQ6Af91cfVObj+gDMNr+SbpQtzBp4yMG5J+b+zXdL
+FRr0RcMkQZQ1I9WtS/RHapi2mYE6GwfwDFtGxBdCRP97rlQSqAc7f9cuUsi5Eby
nYouGiYgNKZdwVAiQQA1LudlZJla1Q8WRgkNh/lIHjTF+XCKZXOnVw9kYf/ZQQmR
kb0I9VciGjhfNENRsKpxjSaTfYAVnV+vRW9Csl1CPRN/xq4GaA0+CdAsrmQ82Uxk
Irq5/6oJK493W/Dsxi419J6SGxQBjZVWj3/9ON/TwJ6LzsuoZgvT+jnWvZuMqY+g
2F59J3EYCS75NVTtYfsHf7gdB4VkR8kQgcSw0nl4VQVuJe+mOSaGqvaNpuChIZYH
rQH1s1FVNlbWiGpH1tOorrImoSsHdzpg50vNORnmE8HfrGl8bXxE1FGMVlHnkvgF
cauVLOo5VgNrxHExBsSBphkvRTnDsmZLUaynhd/F4BsQpaE44sbpjO2JBhQ5RYJg
1Q65idQEM0IgE2Yha1iV0+HcXfSpa5fERbjTW1dFi04hUZXC0HjH9JmcKFoOmBJn
ZSL5WLiAaNigEFCpPP2uuCEntzShn/ANZbQnPhzuS1TB1EsLxEBF5qNCFiDtYRA3
0UMIP+21kOzvO88VhgNq0bOHPK+FBuTEeWuU1jNds+mYkaUMBQBgUo9QA/P/45U/
hfRyg27n1iP4G1PtJYi6iQGQotspyHfWJW1I39RViqeOIpC/eISKiDoYnvYlBSel
BzrP6nUNZJJ+qw1M3SHDEg3yzrgnbwDBprmUjVLsordNz2B59Qk1bolUKbE6mF5v
+fd5x0aJx4Zr+bkDtLDjAwLQANMNY81ilis5eFpLlktHzFfCQAXQJtNlzHHHV4k5
u9isjCroOqSUrU8BpsDPeNgAqKIozkimsYTfPy/5UDVJ/4E8xDDLTGuIb2L8+R0x
tR38o5yzgTlPJMI2QvVbkIeN56M1webnN5StLxjFwkVmQoDWAOq0YFx3KHU4iRVi
vJw5pAX2lyxLKp4qdU5VIuORKrE0tiS2xqOoqBTl2QKWKl4JQw+AuyopB3+nnrmp
rPCDIFodb4yu6JieXtoP9kA4UOyFYxNujjxuMHslT5fcEdlDBNusNHtqGQ1TGXQG
X+b45O6X6UbRqMmpMLviISZOhEtjqGPoipGe1SEQrHWh491o3cOw2emyQX/W3Esw
cPQEMTbjnHHi/4NPx5rwfL1jzA5kt4YFje27SDN82nbo6sVPEHr6FJ4Bt7ZTW3kU
ZM+Iw4SdJR8NCJzIRTQxjO/O9jHDwXYVY+nDoG0XD615avd2+BqFBLQe8Fefmq4s
hjsiEwi0w6XIppv7CSVN6cL3ahyFiKm2Dqmt37yIXNYmsU1Pt3NqqEZuUo0Zn+TH
H3r9C54fwtnpAe80z1pNbcXhI60cnQbLvhkL3QbDp2hWauHkHcZ2XUob2fFM2GtI
f6em6HfEgVeSuweX3dBFKqx5GX/U83RQWxpsXyGXqkqzL8ckyl+g/vWOcywlRLGM
Oqx1a1QUXPluvz3YC8xGwrI5DpDG6hTOumx4ZQy/pA4+frfg5VPHhrTyf7EtX/ks
sqlOP0G6jTnI+mKasuyQvMZH7P7xOTlI+3lQjATwf/UDUNOx91jKrVWwcvQ6/ih4
OCuZntzr+VuSc2JfXeX2qjvuE6HGFoILgVHD4ostXRj2tLwH6EZskm1WmKIyCcrV
RblBIjYzCTe/+OEhNAq0xMwllDjM6ASlibdDXILI8/zlk53JjrOUgfWwYhh4PgYC
h62vRdCJ/WrD3Yv0gjh4vvFzIyCB7dJaTvlTLvOdw4IADHBinM208o2Yni31sZyD
5juRGFqn0vDfJEeAhDEFV0Wo69pfbn9/cPhj8t9K+XUz9am7TsJZANikml2eF1AQ
TFnlwoy77paHrNXrAeyBkuRRg/Rh3fLB7Tlz7OivXgJ84mhnDx6AaQ+oqUYlk8h5
A/TuqM0rkdyHyQo13rCMY3yctx9oIQdIPeMiOrpJSG3K2u3lz9rUBu79xLFhCQK5
VTEAB0X5OzwTRYmg4bXi6QhLj1Q/FA9kd2wMSK71MXsTuQH0Ijtd55umdSOEfeWr
Dkq1gXZCR/FAnlQRAdbOaK2m8NAhQxNOn/yMn4/h49UEkApONiNbB07UJ8BorzEv
lLpt4ero/rgIG6QFDmweA0fnRwHQJTP+1h3Kv1uK+129VNaFrX0r/E+kEG/AZe5y
Wrn7MsHueKieXP1habZPH5BbnAD180n3bLUzEFOpQzCz1lljhPgvCgpO+FjZkgYj
wiSi1ieDFvJLpfHZ/kHoaG8JHAciEn9No8jzRvpY5qnUBbeJ6uFlCjppTXFj2sjs
VZFOVvTZUZwwIgjTsDhRrvai6CXLZdy5kGk0aiz2U92Arwc31rvJosrzdYqLGvf0
WzRWUV0pblLrzQArWOTBMypKYDcEmvMhPqBWLXy0L/2VHiSZfFlSac1fTR9f1ZkD
5IZB367RqV8gYWLUIbDcjzJSJqwaEJ+wT81HU087WTE+DNauPtcwXvknRdB3W4mU
XqRB5MqmrVqY0zhj8gYBhx47TfVUIF9CHZnbjctkPUC8yfzl4GTF9fdhTLBGy8fc
GD610EDrhpgu4Pdac5/l/4XE23g2qtE1TQv9Q+ghsPIGFLC/SgXQFKL+m73rUoCC
QY+s2je6htKuLrY3WkHQFlIlmezhUJXfKAPErQbPhJvEd7WH0CXcr1Z7NreON8MH
9jRgRDVU+t2cHyQrkD2eMCth4yLYoIIte+H6MsBTZKha5d5FDnkAq/9MCepKKAlm
7WMKhonR58kgRrxYd9ovVR5pctItu+vmKWuFDSXy5Z1SkAgKcfVE4lEaV3PKy6Ns
0ro+56U/cfkw9tCV+pR0jSJ2vC4tEqCfAWjPn+KKHIA9XkPI1XaN7r8HIp/dbrMi
EkFq7vNJrhGY1msePjYSVGrF2H6owmVlf5A0oSEeAv1TA4m931nvmoPBeREpQEgR
sO8tr9zkW2PD19XI+KBaNeLlUVIIUI1X0iLKKktpEnVADoag1TMvTzT+PP4OvM15
u9W6Qhox9Pxcqb2fud0ZvOyvXffv6v1oboWTTfyKgFn9zNlBFbfZj5rKthaxkEhs
eYxPUJG12OLhVASvDRAYyNn0d+ZgBdK7o0rWRQRU5qK7CJI4yn4RBkOb+ubRYkRl
/TfW1HQeNVpN4Tjag+hcH+54bMZ3SH29iTC0OQ0af6OwiB9oLQVkS3zcIIB2JRkY
HnAPFbUz71MobFHhBNeDo08J+HQbkrQOXwuiOBXQWSlRqtZmB8LJ3bPF7qgadEuH
hntQEQ5+rt2/AQLm22gjji4gi3KH6tk8ojsp5gCdwaqYDyIVKUAFKO53Pjk1fjqx
t1d8RHhQF4pZA9hKumi4jip+i67ck64jxtrJbZDEQUXUUes0GQNUIKNMikO0xTRB
M5+gkGi/3dX7p5XYVp8IYc3GDYPNUK+MHG0Wcg9pa7NuZ+9UnQyp0d5sFO7J+hCH
Y5bqS1fEqW4b7TyZCbIyI9eAEoWQsNexLPRqzAmqwoZV0D41If02RGwISbqIY6KG
+2iRZBtqI3WlafNPh6gsAhezz+/TKfAYkVtryomclQaqT/QzlghuJCWWUnpcaMtB
y6cCIIwgp+La9XHcUCu7ilR3hqAaTvotJwfv82Rvx4QzwT3xMo9OjbHjXAb6o1+d
GsGtyCFx5eMqNM22izYpwxiEzISm/HP4Kwmrn3i5ZH2Zg4zsE+fgj679IvgQJ+MO
xgb+zBdODD9LRZXUBXPH+o4uurZ020oUzUGhj2jJcpFhndfrU5JUQQAOTJnbPChL
AJQFdLm9P5GdvJis+XXcpmS2mU7X3HoNUyQB8sJLxvkkNr5qV8sOp9F/wLghArDa
RWVCaJflB71bYOmjSXK+CBwfcvSfAFmBB6GzrxLKEJ6IDbTj/T4TrTrWpSCOoiX9
Les2e+9kCRBplr1nhQVuha+315+Ac90akaKrHEJINNmDUa7R7a0Vz2RF4j9hZ512
5GfXY1J42y+lt7yO3b9cPflRIwwOJlqLVnsg8SkkNiKnECCqMRzKj5AXe447E2s6
SCEwjFXzMlfVbxaEkJmLaUSfxXMbSl/6XUbXx/wpZwqaVe5ALYi9GLMySIXTYiol
Lu9nHaI5+k8tc5J37OVkBzdS7BLCh18G+N4UDrYLMctRewY4BSQMR+ct/N4xZIX6
IuVET1QJDv1qq5tfpA2iim2JDHoHzz0V7xncLocNTBWTn4GqaAATGOLc6ZwEGW1B
3a+5jAf9Qm8ayTQjfYPPHJ/mmFY7UiSXZMeuWnOvclCDyfMNFyr08kXClpXBynsp
ILxQA/bCfA1khvuIBwbHgtiiEnNRkfvQkVf1eRESfYMQ6wd2St1K5oEQs4eA1INN
JptX+meVW9v4C9Vev/EURSOhdTtFvnPY7WKgtgKR7MbbmxhSg20i57qOudb15T4J
FprouaVTO0fWtLMWtTKLNdvZHFLbl76RMurt9MsoO758KuFOzXzMWyYWO1RLxD3p
6a8SGbVkfHeoprGIHgiCjEBmqBjzG1AN6ULuzD+RoJrNi3r4jXU5GJoaBNqJz9dg
CiWEtOD65v2X/Wb0+Z9AWeeWWlY6fSV7y+DY7ncwz3rnVrqufPZiRfNfn3rBW3e6
j5oh0rjcb7ZOCZqpWnpIOI+RTRCtY7hK/bMfle7B/vbkOLmnRTkNSMYXEEPcp9Ys
+ayNTEJ+/PEl5tqo7SURTqUbBrBfO+Hje5Ku1nYk0ArGkFl5kUkuTaS53Uk4aWuS
bjU565+MKoXCfZFC/XbyDDOtvmD+za2jAYDzTRp/Xmu0PJTmeK0FOrcNzyrxzULM
zkOI/mqerQZrOBCjBdZKYp0Q/MijE+wjgRVb3Ab39DyM1erRBDnOgqn2W9PJrBL2
TWy8unOGl5wZtIQGLVKDL00ls2/DbKRDsqEUza2isp4d7X6Fo2CAAFYjh2YbRDGn
VhN4VnMIcAb41hFnabu/ad8cm9AkAzPNSLizQl9g/triNoYg2+cC1cYOU0dL75o7
xnRPGNE9gwHtMhxyc7OrwD21arrhO6oUywNDTEchM346eosA4Bu+qU16UBiQdbyl
pYr/tuwRASQIkIx+3xkyi0OHjIrJAb9bdfZo0ZXkS63GXH7Uuk0Q15ZLbM+kJ+C1
vqFb/e8Hcp6cYzSps5thHrNO84YuLeXC3DrLEunOeYAhP6zn6G3BTgHxmE8r8ZSM
kinTLJUnKg+PLS41zbJ/Ff0Zv1BpNHBxPj/7KRKMR/f03nJWmEhvXU9zl/gMTr5L
gUg+ZyVvk0z+ybETdh3ZntLSSWlMIs0/J4iu+Jzh6HKUplGJZBR4Zqg1gEZ0v+/d
4HwBKlbxZ0iyug4B+4L7iwfPaswEMZBNeIGMhSSNdPEr+8+pC9lhfM/XWU0SdUK/
GZxI7kyWJtD0JiCOyJjGFXbDDUbsI72SqO7MTMWkN1P/72ijNEdgV7tRFQo052UE
DUDwXpUSyNhmv9cQDaE0gVd/N2SEDtbK6DD5/0E1bAnTKIzCKF5P1zgHI0KtnpmB
POd4yJ0siJEivb8lL2ZiGJdBO6ZqpdKJQTgYmoMCZYxX2XC0SdaM6T3hHEptwQNU
dRnkki9Xa5cm5CFaPiHPMoxKOkL4qJp+0mhV0eksr6qtJvNXLNPOupZRyWiW6e9g
8UKFmuL4sWXSDEAHkEofwf7jDriea827NK11HmvS3iddHMhAxCKDhoLVdtF2oirI
beZWlFsuw8AIXgE31XfC5/VDCGHAv4q9jH8NLvjLR4qV2m5qkQShlGnhiIb0+9cD
MdFOsu+j8Om0XTYXWrFAHoW4jPqMdvBBzkXJfXr6ZzkW/KDOyEEn9vR2ltSh+aKq
36j/MfpnWOTDKRBIrsQBE4B1tebQME2zXORRZQbXJr0YBv8GEMe+YXpJcctuQf3S
JFVGcw4JHzcbLjZpxf7gzU+WeGqjATa7zbBjEReS28mVw1YicRwwIfmQJUzjJxdP
GkJrQq+e7JSyHHmVC/e9mOlNRmntXWcpIqjAb+1aXxV8TVf+6Y9oBz3cbt5dF8Sl
P5auTe7Yfu/AFLhxEDeRnV7T1BT8T47rGA6uOn8bgrGN8fxfYnCIk7tXPKuSU2PA
bCq158zvXKYZjUOmTnw/B3Mx8xylo2ucVy4kK6lxMiL5ESeegXxopQSkNbVTBdI1
DNAeL/8H+doM7GFnulkW5YFdXoQ+t/NfBwct6dehVkgYDgwztTr7duMCnHJuu/Pl
BacLX39D45PddfhU+oeenF8xDww5ABW3K7qCrviaCFoY9ykKgHp7lZgmgJp3W6us
rkwQcjX/r1WR7cpfRtUfwTkZy6vuV37/ARzSLxvN0fJz5Lv0IlLZ+KKksyHrbP75
KwE5NaKthsSKlgem84etBbCn+DQ+T0Z1VCPf25Wykw3Cy3ugOAx8xTtoVNvCqKl4
jPKZhxRNcUMvHja1sXPVaZi/Gbk1nAwZNuWm/xcBNuf9aN1eNuMxwHWtEEI9kKNx
CJJYGqSdxeAJIVEanLyUfRRehU5xi7L0nFq8DNblrmtZ6Zl8EOEJU/uBb1wc2GC0
rgispmKkuFRrG/dsR0RoVZANM/XDu9Y3JHNXpKx5XZurbCsYViZW0YL+t9Co4/aI
+XzkyKpCK3NX2DCgCuJ3TYJthRH33ebZ+0kZkDsMIGtXshv5z3mHpckCJ8Sq3jee
/Xo+ApXOuHlAEbyl6WnpmPGjBWYKS1/L20GLEH7THMPhglkDRZ5/lDziVd/YQRg1
k9Qw4WSEWFOcr01qmMd3glVY193927cdLz+d4pPSXYtKv4rIJ8oLHWMUIr6CrcKb
edbd3lHOXm6T6N6zxWGmaR5PP7cpCRYtNf9Qq7z5TRculR5klQjaWZ1HBxFkXuFP
VWpbzjjtwv8ERTqYQ7auNkOoMgU25W+aGq35y1CK0DaxEr6YO5H5txsA3g/NkUYb
b3/f+3zmQafnN/i2E/jL8x+eWnrqnGsR/wBh2yLClb1Bwkmq15dI4RfxF7ebfAOD
McEzeSMHXI0f7Qn6xxo8M9vGA/BhabKcEGUZoXEv/HMsEkWOQoKd+dsPAfrsSkQD
0en4lohM3moRit3ToELYhedjkxi24Zn/HwL/z/ORQ2TeHzfDDqC/ROAuBF/baldq
nVc0tespETaleJFdHpgGRiPemFj6zSFomjnIhMQaDWnfK0BZDXLQx8HUDNKY/lJv
qQCEsQY4Kh6+RxOYRT/ypT2AEKUFHEdlljQwmeRT/Z324t42qFIJDj3jXAWl4LKc
MJF2ZC/mrxXy1zOJy8K5/Tdt8fmGjqL5dyyjOJL+3DMMFl6sP/BvKYmAQDD84YMY
nk/XW9mTdk+TAJ5qa6lgtOsB/T1bnAyJ3s44wPK5ntAKlkDAj0qvO/xd3s8Zpvkp
fKAsCZwCGd0tfCy27rLxtWIpYZiz9ocDeDgDcBYyRFsHqD0bwoTb2cttd8xqQIFd
PO6jvPk/6h3orjYQdknXAqSWK2IrTxH3jUKBTrZDxWjq+YKf+LtJqdydKiSdy4Ug
1YWenonjVzbE2oMAd/PkVUvPugvfb6Y6XBI6nybfQjika0yvxpkboyAfwtjxqvz9
xJS7tN2TSwufSSP8VMYV1PvMh6W2k2QPLuzXOhvO+SQaF67oG1X5mvflheJpUFu1
KUZt0GFb/VimOMKjcW/UyDi2JLmIIEI7uANuEiGpspCeZ8bUkR0EsP/VtJqygN5L
FcrDXQGouWk3Yd5rYnqKo6jJmKFNm/cys1ZYna+1nbYLsl6P60Abx6VeThUhIr14
n6B3GDTTD1ZF4xAluVFdYnOqSC9jBcqs7QF2bBfxI49DS04FAPJsh8avb8R2UlUp
rs60PnamhfJ1WcRbabzyzV8P8UmObmaIcjZZdb9YuUwj/2ux2Xe9rr2zuLxIkm5Q
cP3txUoEpAaRA7UVPbWxXAhTRV3ZnRZ8pYzalzodaUFvUGMPHcTdfuxFAGoE7jOg
DK79MWsu2jq466qx6KuHSALHjhUIsbM3LV88HbW+YINrPXVWwxD6sE6+9vv92MFH
jqgmfiGhxKC7V6y0u3fWsNlgDgX0v9iMLHaZANjpCunVxtIbgNs8hN1qLubMk7qp
r5bAK/VN8TthRSeq7e3fV8uMlZhKifBTlJkUFsdPbOUtCIHOtKNVtgEhYy1CN/YY
nDQRuIl5ejY731XnVhYYeHoFGBOwTt9zHDjjNJfxjIcqi+yQiYn4uUX43XvTfy84
3lkOEwMKI9FEMYLlpIkD+zDekMcKFYRs0H9Jdc59Tjt2W1Y09tTtSk2bfkdzPzTx
Wer2UhBxT+Sda1NNA6T7i4Ceq4F/gentssGaa13ejad4fqIafGHnsIs0MDP2z686
1zLfXNtWQkstpO9F8E82K2I6Rz8zMH/atkCqLLvb0wWRX91MrpwIlzplnghPbHoZ
J2gjh5qNJu/Xqs4BaqZC6VIG3LNW+zxFwkWyrfOTV2WhuRiWhiy/Ry002YSea0dr
+0VZya2naH0UQIX+sf/JPWHTi1EjFhV4cnUW4mWbl4Ti3k2g2mJJanPFuCQ1B1tz
PevDQnMBvH6P567lZgA5A58wmOeHGEW8k9FPpdwxvmYnLpPxOjpk4e0mK/V0nYqb
DTXPKl+nRlU6/pK93cRv4ph3nIdPrqwfU1MdcvsIhO2qgY5GsL1HDh6LUsl4E3zF
rSY1ZQrWLCqcIExX7dYFfXr9PVS74pvKe1n+BK56i4qLTGDWIfuK2+5GavCrIDtn
2WRyriyA9AvUZTbiZdwTByTVz4p+HTGT7c4aPoLgq9o3vWqkFn+Rg3rZiSlKAViF
9eA24hWCjyuHEHxTlfM60kABV1NOyz28z+5/6TAfrd3ulahOSFxon76UVaERP318
GA0bZY7jF+lNwU16rtfoncdLoZLH5E90An4qZegQ+I4NPrazMH21ZCyo3YGYCK+p
CK5y/paXe+yVXKWT6QJ6bm6tBtr1VggmtrxPxE012sLBm1QA4UsAMdepFaQ1tBi8
eOFJUBu/jkdWqLJgqMyAoUOAUbuu3PdCUZeGzJ0FAmVMHOXra9R5I11scHLriJGn
nUelePuNoOwcvERjLbIYNZKcXrDbocArNbVNrl12xpyztjk9wrzxQ422utorZtVd
gnciGXoNb8Pe2nWBQ9M9RkFnHgla1tb+GWiz5iUOlpbP3FzUKaqtDnEZYhZqA0ig
g6QwEc99fjX/1R/SpH4xOPoJ6pJmarzhvqAwqTM806TLjIVVy6AFoHycS5N7ILkb
katUpw77LH/j6shZvMgtuh5o21q2qp2mE+VvFlkj9efYwISkH1kzqL9lp1FT7A3p
eJppmUS6en1mD7dQj95TuG3dmvz/L/RinrRHVNCT0ABLr4MZ4OXKUeEXIUudkIZZ
ylQ8NCLyahDofS/jAEXf3sy3z8KRUyZx22p3nd4UyZRJZhryD1Q3YiEwG+Psim+G
NdCTuJ+CKqkOpc5JNeIsiGeB9JghDllAPJV9VA+W6U6lHZHhrV7lpTUGQQANSpnz
690bVld0yQeStaAAwFsh1sr6SyKwG85wvRPNDW17iz2gjEGk8Ev7P4Lvx12s4f8x
tgdA4IRKO4PG97vbfAMHzCnOyL9i9sPvUPnDRGXGtldp3oPxXjjH7PmhBL7/wyg6
0yzaI5vrUH4xpT0myvKFyqo1sjxSfbmKInZxVoMstvRDyavm09r8tkLXb+nM+2YB
6SxnT/gROP9yLmVof2RrD9GPKEJGqwn40o4Qjoi3cW538UGK04ZDRL1LQcdYNnEe
D6xhuW5+HilydD4OHu4yyZoARCHD1Q9QfFc37AfBm0gbNBGp7yVF3RW5wZ2hhl4n
Pt87EfTEVXGEM2386CYzATOuz/LLSMuJctO2T567HIW4tnALzfwWqhiu+ffz2Z/w
Qo11cv70x4PJV2tQ0KE6jIdW0fyfsZVg24jFOSak68esmPKEq8dN2xsoQsruaItA
ZkZXy39F5YMH3hoduKxdAii5BNFA3PbrMjrJNW73yW8WzVSnbwnVXYEZzHNzoEN9
nfmuupWXMyV71FrH53EfBJ/TN4Qt9ogNq3NvkEjqh38wnHUMuLK3Yp3IIXEjN+G0
J67HOksc9fa59JWZbFVa1HX2lt8YYU2gLxFh3DPByNGTKAZ0iPSOJd7CHOfqy3Y9
JVMIglKyXgDz0EodIsbO2JJT4QNeVYecp/1SFahMih2TtqGOJYjCKM+eJxNnH9Oj
ymmDf3Km4PK8DeXtpJJyjeVPr1IxT0P5zjDROrFasRrydCIHmXxlfHetsbJuWbjv
Sj2TTx/io35p7LEB567Mb/G1lH4VerKdSGiBxxQHtWeANYvR6WWvaOEpT09aj8IY
RnbiV/95uO/tvX91msVTWrLEP6Gvta6KPt4oMJ9dRcefFu63eDj3m5JjD9R6L+YO
t402dlWdTDzA9/3pYw580hqrQGM3nst8LqLANw+/6+W6ncL1VLS04NYbGGkpi9C+
gFLX8Rq9OdVpdHCSbz4yOPoRxmQTi/ZKsef09Tq7YEZ2CiGJgXzeLnKh84r+0wGS
GFUKBTJSw7QoTHl2kbn072rPUQXiLyb2Rth59geBzES9lzSMKpY6he3eieY06kzl
ygSdDWFJ38ckU1s4N2DDRD3wNtEy9UeAHto4vZNa+sMzqgbMGLH9rT1cwMJGXVq3
FrzVhNi/6b5r3G8e+bW+oW/fglzgKjfzlmrTjI1++6XYm/tiHHkKf4VGFPTFDip3
6hauN4c02h+92wE83JHJOPBZCoNHPNCY+KoMPZGMlU2HK4aFYzh7ZPHQXXDitqQt
awFM7i9vylY5geF8r39aEoFpFAI8UHAJV6aw80zfMeulJWB5dcIr4ZCdtUI0DWdz
H9z5zoSkvcXS2+WFt36t0v0PHsX/VBl7QopBfNphwhcqo1lSJlm5XCYTl4iMHcCQ
X0G51hafoq4IXZIM7udrayg9jaOFwEqxoWG+/GIua1DiHpb22CV5xq06akyhpQQp
qvHv1zPSRQkTe0EX0Dyq6hbFCVTR8N4kZT2QzPVdOJwP5ZaAZAFfoteTevd/drmO
uF8akKwaYaKeXNTmVD3T7zaSumlUhJMJi5siSFcR6asK9GXqcIVT9fLc61z+6KHE
A7+3otLXLQ/FeGC9OR9c56KAtd4bJMHemqrrkK6TNGUYW701dhU/jcGsqEEXu8Wm
RYjLO+MoNQbK5FG0o2ChjzHMNNcX8qctn/Is4xq49cjGLNZFx9PfWN/RfC0I0EMh
HpqX4OiWCrInNKU1vrc3xcGbdjE3sTszLiSE7yzDaeu0eOfdBn/xxYYpt4I2lcJN
3FueTC8TdFr2lamKXrz8WfM1TT/Ry5Oum7057WAXzyc1cWpXurgMfU8JtXnYqS9k
uDy7obH/aRDUZ4Kn8cG+fdK5If5sc2U/8MjKHX4YQ+zehRJh5iFTBfsoYzY7Xn2s
CEvPHlQeYUu+5FPJqZimvLV+8thUK+O5M8OWWVCmgb8rORS8PbIiI4qmZxdbmYP6
qE754i3LeETxQ3oJyizxeeChpBlAKOA/Ll0BcD0I8OFaoMxF5k3PdpvLXmVvD8Eq
GPr5v2V/c1jbqwLCrTeRM/Jtxg6Bt3BVvnMwgeZ2tZx1FP2TcKDMQ7iqnN4Trt/L
VSeU3mCQINwPx6Nmcvl7UgquIucLjtZaOc/+dOE9jECKoA6wKxcS8SHyuzsRCu7m
/8XTAXxe3d2v+oxJ8vWu1vFW7dnx/yl5WdriUDU3cI9wZjmsmVBq8zlca6S02/7F
OLzE2oiKXKXr2Tst3wNWFTGNOdzXEmBbs5rmOAv99TpJrliMtN9HOOiZ/P+qUaR/
GbQa0tL7UvJBsJrt2/5zedkBEnPevUIkoijeDzJ+4wX74ii5vGivFW7ylO6btPBn
ig8r4KNfI5fgmb06PJzExSn7T+l31pkWKBB9xkOx1hfdLHiDOvvGanNC77otQ7Mz
cN/py0Y8ywifx4tVwNY8gnPDCG7EV/hR/NRMEqPuhFcCcadPHpu7T/6oSlHgTt2j
bDuywo+g+nbkMWIlKdSaQopg67l+t5wUZq1fj75+yh/SROE/Z7lgpRskbC71MeA7
J5P+QSsgGvScsdp96NvmgYuambaS1BRtGxWuTKu3VObba1vF1bwlpthELx2/YOKe
mKGPgZ6nLYIxSc1m3ub2rTI/7aAHao7F8D/OHcuYFrIUbt40+zq4n8JJ3XSLQx7E
7RdIrmpRwWgGsVo7cwfCC/AUiWCH9K74cxPo00+SkxQ1z6Am2erffcC1B8LJ9Wnv
pm2ZvxZlJzt/evOx1tneeNAgMwWl8ndI32/x8ftLS8mtU36fyeBrlyyK/UM4f/GS
balelXHiLYsQf4X304H8BrlRGl3VnhdeVquWsJWx0UzsbhBpBjeEt83qIU61V6x3
f5D0i63LN8xl712bivv9HutlTI+fvLsP7sRdoG0mw842rVVElmGJI9CY68L8N+l7
+NQxvRLfPXzI5iBOrVYy+4ZK9WDj4KdVSRI1ChYuFRUiTnk/CUihVbrbPXji5pM4
BWiClVMF6TVO/PBKGhuY2ftKtuA5M2RuQLl5nHsoXMPkZfcq/YqphaCyzk8nVVnI
nANQ3epLSvUSL1/iwMDAbUdswg40rWykgT7O/qW5EppSYF+Vt/EXJTJVhgNwQnwS
TyXxA3x94vIwPkkzccwWFW8+6KBjR599T8+dewtgWDR5aM1x2DTV/D18yR9fzRWh
OJ6b6eK95C2fGrqbtoquNC7SJoV5kQG/8HqMDB+3vCMntcCYI3NkEpt0kPr5kAxh
8dtgQwZB4Sh1P3NoRPxpbFezghVTK1EU80/0TwVsGENTt29zHoYp/IwVdtsTKOQp
o9VIsqdvv7ty0zN9Ofqg4tgtx9cDVhttGY7t/kJEayyOFNoIdnv6qMjdUx/u4guB
4KVkzf+fN8jorcJ314dAkEgj+Fbtud87u8auIncLRGUHCwkWCpEiF42xjDQDlQRr
pn4Zw2/AWpFOt4hRpEwzSHnDiljLXO2v8NdX0y08IidrDNvkA8MBzyobM3pa6a8n
8K8hSKW18C6gnJsya4Tn60+rZ7aCibRwbRflGoKMGyr4DFyu0m3ozTwX5MVnROrj
xx4XtVi5egxVECv/Ed4peV5CeegsdTvXAmMdUDENayD1lgVTqLTWcXI6zGSxz69l
fBHk4A/X2FxYjdh/3o+m1KzYqB7XDLlkPu2wq22F986wTsW+KLSfW3usp2hLLfxb
STIq0TdF0Ew9NHsPqohLCE54E0xVZuWC82tyH+5QTNpzyhAcjpY7bLm+YakdAvK8
OiqjHL3fd9sJzi6jY1HDc0lq2A4Kfyac9m+Z0+WIBerLgPX3/jyKf/0l02ngzmAw
zr5SBfV0PekjvfpAq/KHwCsjHjbInfNd1vDIDtn2zW4MrNODrVTSx7cTAjpeLA+y
WhHl1sYqEBaNrq/qmINYVhd5X4AEAjDoeOde8eqTBP01YwtFOEV45V8tHWwIOU+k
d+RTiW4SwNv2UnhQjpvtSkYHwwHJKOnpjXjn009E9GGx/P6El93Cr/mCAJsBQzP1
A3Cf0BiLGv8Rus7KUql17SRNePKr3Ex3x1vPQoyU07daNqoi63s2GDs+xDFgfVKJ
t/a+H6bLxVD/qxkkEVkCOo3yP4YmxP7BBmTMCrPJiewyJjJVjOyaFRKOufg77clg
aAzPWchLKk3O2V+ckBVV6AzhGFRXn2c1pUje5bMzchcMHXxG3euJjPQNu9NgPAcp
Gqr3vyI1+ZFNdooRj0sJGJXWX9kBtAPqBYA8N866ARSycBgUI1f7V1v/+10CJAqd
sw1epe3dPx0cFrOYEghTZ8URI3r9Kxj9ogz3XN9Vcn5YCIvSO08fb/d0QiTQPB0K
ptLC7C1zdurAoph5I2M5oP11AJ5Lar5d9Da0cfc5ed8k7fUWS6gugUpUM3quev/1
Sx09NW5s1JDVNrTyxScjRiSINEEoPRitR1WsqFSe9zLMkgROGzOzAKPrQClnxAqp
UomNz5aQjEtBSERO62F3NcpzJ/NriIPLwUIo3Grd7LmcSB+JzxllJ8OckOa1IAb5
a1zTorJ7ni1I6xmgnKKFSGduHuqKmdugliPBEMMHr6xkJ/Fz1aS+Z+/D5D8przJh
F++3eFChPa9qtPTOpdIeDsBj/XuZMckvbnlKC6YnaAJeaqJfCm1VGrwN4ps+pH3e
QVSIqt5MJ67/8qaTOnAAq7hE/Ad2VlGW4R30jrTKiLyZ8LmTePWqVrZsw2GowaPW
bhcAV5JBIXn5rifAki7hxPv8eCP262Y6o5tXOvDWrMdLlmW1WuWI/ppSQGNptEiO
aSTrXmk5g9Imv9tk6IQuZqpMBG0XidpUtYcglYN+pvH7a+PWkeWp9Q1F4gKdkw0z
DocjwXm32z3Tn/FlXMkH/1Qe+9Kgk++gi0JJDcSp6MOPK9PKOscAtHA2dJkB1ByD
IWgkeoN8nfHcLhm68TglK0qydsIgFYYbDnwLyTL9gh5jeH8qlPnOdji34JA4L/4t
fkrNGhgCcqHhZ3laQMlw8L9pzQifGqgL85VtaK9nuxpRvulIuyiyFhATAxcWK8XG
zi6vppY79FflEjJcOrA0u+WlYZxwl3ESl5Mxk0FoMctTGHqhRjvjSf5qoBO+cL6Q
Pgm2t4E4WJSJbBg7OarRXk1ySCjDXiT2D46ueUxYvoeWLiHTUpGWMe5J6IOKlfsf
abRx8PDdrXzxuASIIjWffVxJbIsoB6+xWutCPkQ50Wf8JeG++XJ13wEApwlSk9QX
outGYTxPqKl8zzli9JG6SPkjyfIi5dT+O/la8oOeS4lgXnLCsPW/LDyQgyb3RZAC
7ClE9m8TDT/yLQtILN0p4jc7z0NlcsLs3s1kvy2SP3y+HyqtSDbGBcin1Q1jjt/h
DeEqRujmojLzI8Y3S1Iy5YgQI4LmMRReSZM79dJllVJjb+19g03RU59frtC3GD4G
BH6wn2+5Yq6o9WGaK7Hl+4D6/aUkDWEhCKhV5YU1V8utftHOgXftLSDRBQePshKo
zDgwSmd59OFb/btQ/2d2jFhoKwvKVJAHureRUqqXFiu8QiHMLhpm2RqEeEzalEfP
1m7CH6KObInasdhxSaHRrxD+JbKN7fwzHLMsnSiRzCPgmFxQkxwnDffr1wv1YfAE
YaEEtcAIJ5MJCdYe2Baf/yKmkG58bZaTePPDROT7iZY4TU08BCAKkTESnjasEb4W
w4xXfdzfQiTqGnKSTJqNdAALxdHGwUFJTy4DBe+aRqM02Z4z6QgHoHBBqnN4B4I5
YmEPrHCTxsmF2mBql1sDsWPJkOX2d+m1BZmAZst+R8D3mSkq/X52/zA0TUtLqj8o
LcpG1r+Mb32/ohyKUNuHyyORTur1bww/i8dISkTKqD5UG+OoDYQ+lFat3P6Fwv/j
2W3k1MpMZtSZkj17ownv07MkbBmf+ilB2PNhB5ja89dWbu+619GENW/2u0WQPEW7
bsT0/56YMYIDvzHld/qpYiTbcSKoJEROh3wGds8v1+dG1xSJc1M9arqkLrNeJnsN
pFFmOuaSU684YkJ3wAYDbVEOkJsON2uTMieulCGtBSSe0c9ALVA9zjSNyXWhJpT2
OS9Qief+6D7sRqeX/r+cYoaQQ3PpY/erRr3sk3Y84X499cFJs2Cxxi+ulK4B3QJl
kTrpXQQcaWBBGYQp9VE0egrwXz7nR2uY1watEKTN+dVf0GTAaHkuHMNkPtKmnEQt
o0qlw8TWvWINsnx0nb4ZcpeFZwV8cpMbiRHRflj5wvuZm9Rm7YwMp0Le4+Ld95km
IeGQonK3XrCf5eQR7NxhdjRZvvnMt7D+QlhYJWx4ig76zadb6bWVZmfUZLRseRcv
9YbzlAQS4vKy7ivxZGVqeX+pDdeWu3RQf9hvZnFr2CKK2p2MDlSy1/zWJKaRZiQY
U/AOWEAK8QjcZmWwiZZFm9jDTsbj2pBzHkA+kuj/23u+tsopXN7WChKRRisl0G51
l/+Or62enSGZlbv8tMW/UIceHFroToAos6hpfvXp/C/nOScoJpHZKVjMqHbxhAlo
xCJ7JZ69j+a/d4e1rOFet4ACekkAGD2Ev7xb1Rih0T2ArbTyVKfl1VRchFudCI0v
Gtwze7Mmg0xb6jG5XsGwK4KADo9gEapetn2CsMItK6Q6nXbkD7kJwWhD55NYKivG
mhFFwSVh/IPHk+gR049PDjbFmTwz5pE8LYhwNa7C/bawmHRXG0lvfjbLJ2yAI9Wn
OBvigwwge7w3+9bwH0EepobrpteYQ8dAaE5X0UwJggSvby08E9V0t/BDOoRT2VIv
NYAE5cXpwJVmOrLRfQvbI8NAgytXmBAwIlyG6my+k6DW+842URkfULolE6SBJscI
Dyv6AQwVjmuNGOX66WJ8yRPbi6z8O6sTftFYLy/FdJ3hyDG0mtC4dh3U3QTnskiy
Q3k+ZkpA0oPeSGHJn7XMLhJ2y5h25F1A832YPcuWP0pbJ+kcoxThgKQ1U2UdS920
vfxt5jN16FGXbCLUykCJ4l0MN+3RDX/lMn9FPQJ4LaiRH5XJViXwb4BrFvYFhK3v
3B/OAzgLbiufbvXUsAV0ihcp6HzhYLr2saSFfgT8jbDV0guEjd0SAR/+qz8ooqQW
xfuFofKmtzpFNOznc4KIc2szYH9+lVtShiFAATHHHnTXDLmDqZ6DsavskBNiSkF4
2w/iSn+tfesLJtgeSDhZmbpljNTeCXLJNzJ5OIr1jP8wLeb6DTzwXyKt2K2du/9O
swqVlSImo9KpsQgOjQLQJvxGyiSGLrqDasJ0+16djpnJ1ka85xgB0Sn66IMTv+6J
iuctNw43KwBkdM4Qw/5TB9BIunLHsz5XlgGZPBCKTBctFvg7W85sULf8OazVDObt
T8sGuH3DYjJSAGFK3U6wwnYngJb4Ny/SRb1U1MEtw3TYBKx06aNie9r6TNqUExS7
SFVY96Au60p5ZH98mFd06OI9GU+U9BRg83x4MLZeRfNrZ0C92LdszSNYMP0IzkQU
i2xYEMaIaM+NpB0YtHHBgP1Up1L6Cctl/4UQf2xN7WmKNaJsgD+UdqxdS4dNrLfp
NzeT9xMeozD3Zqy7fE+sjv2w+A3YBI5y5uLQI08s2pH6QIidDREqb66GxTPyyIOF
kNys0q4OnNIHkxoq4VFL1GAVjvJt2b+J41hHPHxnZY1/MUVdGFPEpVwSw/ES6V21
H5thLaQQwJDnKWchIgj/QjvdLOpe6Z1FP55T4BEhz5+rjVerqHHMBMPv674hpZ0l
7LbOFWkmo0+v6Un0u7Mq0Xyf+psWgvGiiLCypDZEmIbJU5OuiZpTn13hZf0Uq+eR
2heSkSHs3DZcqxJNIpVcLnFlwbL4RGLrRnuSgDlzFTgZcyU3ErHRhisp4Kb341+P
H98oZrYgM/c8gyZG7uNtR3k2iNR+KD9AzJFM6AK8TaXrlRQlbuK69qIyTmGJ4dBr
IfrS4hZRHyARdpdhTfa7n07PEmkJvvnfdVTupg4gU7k7suvAlb7tI55RndxVH/6Z
zCc2MwRDCOseemj2a5jCYKIOmjS7vgv83naCuoaCaFZMbHRIiRBcoEYJCu+3FMyp
nHqRwCCx+vLRrhPdN0SAIsWjpGVzpPCNyleyp583SfvJiQij3OQnYx7WKbSwumj3
IAkpIiQg4H5jqOwrYlPsDRva7liKEl2cMtlIdilAldXTiPAOwa8tl3RbcdS/wHzO
X14ZrNJRrIlX3yJ8rq0SuSawSfZPMhGsqAlzRzdx7rQ/3Ukzxm4QX/hgGVT2lTU0
dfyYZAcb7Y5YqERW3PEF5LkHLH2gJnaKp4XCuj9nuTuoFVLbR5cCBA87GqenSFY9
P8nOKNVvLUAC+OKgEl8tYDEgGXuXZ8wC3zuR3MZvatbsRMAv4CMc5z9W84+Po/Gy
HwsBwdw6JHcTDmv9cUkvMKnSogTp1s0HqiTPhQecrtW/oIdy/iMqR+/YZjpmDeqS
+TgjrBZag7WKIYWhjwREAY2buwIdF1kIqHGU5NgZg0cJylblkQR/s2H1KHJakMzi
ZlYTpJHegwYFkpNeztd/ydW1HbBunyD38sd8+KmYbA2nHsyrRytBIq0wD4yYhJw5
kg6aFb6fDBUuArNh3P6ykeSwhdX1W5kI0ZSrdE41vIAP1bbW9+l0dtXix/Dg9gYp
i8CaszDYZ99Lp/zpOLBcfJZIr9WQ4QKhO2LWjIIUiig6jFSAzLSMT9aZMv3v6z8O
DwNbEmKv1J7qTaEd3dcU81IvBPgUkRvrP76oflJ+7N7OfME4xoWpmX63+U0YQEVg
dcZyuRYVF0bmt/9s+mfCX6t9aTt9f7Aa4YeeDT/IzI7rGDLfKD9mE+iGDg0SKao7
WKI06mdExEnelbmUyhtwb8HYcnbaD2+azJVhT8dK4KBaV5pKOTczGl90lPK0GGtM
JC6TyoU6Nmc88VrWcWBQTNEenTO3Y/X87Z0/j/omOR3BSDM7jjfTUPlbZlLJQ3Cm
O7o7C6rOCT0A4oj1nZpN+aCDoab19l/LPgA9LI/CuLUoThf2p7ah7kLbdo7KX7XW
N6xzMYdCIZ//OvciOEQQoeBdlDe5A0RCYWoTT0VnpL79ENUDAdCXrnylFU08NdOF
ccJEchJnh3RtnfuDKzSScatNvQFcPevk9leQOX8zdGno6SHthunXxXCQZh5KWfxL
lIc9FxH7iAM20RJk4EGOeDOGJKhCJoQG7xjK6PGpIWVvaSw5srPwQUm6HdSjwllx
0LVygeUUk0BlEHUk2g9wJLm8DNpPO4fSKNrtiqVHtFxmzC7aX1icPQikORY62+zU
9QY8IIOCoQclwatH6DZTzQnyRGnrApDpSqp9EqMg5LugEWnb8z9jpKx6WcMHq9Dv
MxlceKqOKHI/ndHLqhlZqlkLFZrteGj5WMxOSXvQUiRuO0Ywn7V27GaVZYx2P9pA
1MRa8eAkCrGilP3h2t4bjTxtvN9FJVw5UwXWNeuwOQmNLSgvNUdi1FbFFnUisS7V
fUBcEADxtg0htIwt7+3XprfXIizQi6ZgLyw0jGkcAEyEccIEn/p65GnUjKYecyBK
Ws3UsTQo4EI66A/eTMxLt3rjd5q/aez/BGBzpg0sWubX2qrvDIqZKnxnoZWLjld0
yjgRpShTR5ByM+itmMcBGHuv/EA1K1mS9H98EaeT6QKO+l+ERmymudqS7surodmm
oo/hgw7gz+pMjdOjxM9XrQBgvxMQznj6ldQvHs+ty6Ai3bWkyE1RzgcoXSwI9jja
xQUzvVRUvt91n084nHnvOnDeVUX4R/08YymPSbhdbx7vMIYPF+QeR5Dhdf+gngJq
cFf+7oofWp/fl6sY7PKMZJM+mXgx+PaK4FULZ++rE7hLSDaoIt2cltQvXzROjU8X
YB4qZYRMz8r7pWKgyyXA0n5eMD1QhV+4agr7SCodMbFQc1wPrYb+iQep6DvYlrMw
5hlhcF3/LsiMhK0wlzQwJwpDGxWg4NCfH8reqpRkyrqLLLBLUWzKdYAqT5cQGSCv
atzCuUixsWAkwyfN3qjxaLFTTA5TEFdgx07mJfTZJ4tPiFCHnweZl2wDtVNNtlnS
8Yxdk1XI90fvNWJhTBQ81a7SWOACNw68EO6+fvpXlqpyoR7Qn6sNvdrgvHyLUg0+
PR3yTN0VP0lV0K8Fi5Xgyqq8/QxNvSJfAeb9qQpDFBFwOJvQn0097neS5UATI3M4
3MXOkutU59u0vGpTo6OiFwJf7q8V/9htAPDcTEuuY+gW7xbxBPAoqRQn77r6eRGn
Ib6d6lJLazNSe/nMhIzVmfsp+fC5MtJlROjEsVY8RdaEll56LfcMq2fritrBTHuk
nHHx/rq794Z5FWCz4NHMRMW5gfX69jRbdmO0olZHO3HULeYynzw0twsr20lBaoOc
NXOtW5rRI5BMvBxgjh3XMWGyal44q7KyecT9X7FswKUXQbloqVLqdtk7K04G70Xz
n4QlhOrJzsSnx1teyGg0/GW5pkW2lIpAfY34rLB2T3Q0Hl4Tx/iffLflVv6djDWI
435UMLaYJCeNaEAzGfW5PiZXvZqq9vpFiJvDt4+hJHvDSrTf0Y2KBgxwIeCOiJrd
SOBVPN8O1fTc14zTOOTdc7nENcfx9B+d4fqIFAQPVlJQR6uj+PPbccdT6Shhz6p9
b+jE+VlotRQ3i8bbxkmUbaenM9vl1FJwHf6bcd3xwd9X+d+v/pT7MgkqmwfQlQXJ
CBFKupHaWqBxe3NX5exOyspSLebCFIiy+CR/HFwcWx1fKV1WkEUQKqgpb/A7jbxP
TjGzudNJ1FBkFZtIM6etZZrMk1/kUudCxAqrN7dsR8yVuKea3ANqTflwotabohVP
jvQwAAscLlZdXAT598Tb7mJ0GtpBfA7duykCdeOxRKvAeykSLar787tTEFCuzDjy
VCSuhne5VyF+bQ62kAsPditTeHpYqNW7iezdeHI9w8K+jG1jpM+b/yt4MdDfL6U/
RKlidmLrbuOYM7HWUTrHt3XZyzwXFjAmAsVBqldkhrjVVjU7N0aibdW+HLVtdDAt
TA/oortEf2Wr3ol9N/l/yWoUBtYTCgHOAzOYltqfcvrPTpeZIAnCpGSCZzQuSfY2
3K2P+Yo99eCUYNbUtK4gWNZ7aXopW7WIgVzgYjnSUGI8y/BKwoD8hcvQeDDn+5xJ
h+nxM48qZTVBlqd0D166ocLEPss5FXOHSFp8YGe+mAc5ijKgk0G23oefTZjZcK08
4VUA4SCTqu8ityjT4PbZT0YpuKykO+lAl5A3lkb2Jc2k8kBglaaQMH8xuFoURUzZ
4FPsoz6wU18EoipwyNsscpRTH852Tl7CsrWfAFy6Tib8ClOIkEiCtMXTpL0/+zFB
17qRJcg+t5urSbEuYZYaF8OpQtnPpHJ4rUgg4uIerPc/S7sHItVeTaJFeOm/JsUN
Ekpb/0JjeDtTH99qk2Y0v0oeQEsZiUFY8jcwrI/aEScxFEWkp1+NUCadBX9t1RWd
IvDWeMsmmSVfdEMgUN6/sg2ph7qAY4sNdaNSVrUM/IPRdunDoziJMASufywvd00G
0roHtYaRCAtp5A2It2/vnXhjtZHpAZyvTtzt+9RttAgXV+Q+dgdUoHPvjhMVm2OE
GUZPuNRfBDQ0OcQywbDzkNZFgkypXW9q8romnVBeQNK53sLaehSH1+JA2eeT6jbC
Vlk2Rii8xp80hJUvUKn3Cixz0synwVV2P47I+/0b0ToRWc6judjbVpXxmvuRAiu5
0FgK1N6cOadBx2fqOGT8HMp0nbH+Np2Jwl42RdmjJXgFUhLOie0re3kJkcIbu+Sn
oIHxPEXe8Kxqy/V7M11aMZM3B/op4eQR3drB8heub0EBqbBRMRLOERrEBSJhrtNy
9ySXyUQ/o9YJ3RAOTtkxlj38TX6YsHaHd+0EJTF2Ae/V3WiKr3RyuDtUfhaGGRZ0
b6PH+65uj3gwBFQBh+CpKDTlQQNH1FtOGOqUivjqMDwWw6Gg57aCj8EhSYhg5ZCq
p+9M091g8dznK7Xjm7vNhbmPdcM8Yv/I+Tw4uC/I1aco1Wdxafh6/lpi1sYO4QyI
KvPdcqs0L/sXWRXB6GOtHZ/L2yERpuOBsUgKrM5Y1bJCQFV98BHcd8M4P3hkJz/G
EEMPMwQtWmhB6OXdacuikiTzmyi47oMFVQMg81Ec/nsq7h9XFIeNRC0uRKN0hAxd
31hxF/Rzr9VD3wRuGJyek7DIOX941cCQQ6dft/ZZeR9/A00VMHz9Emn1qtJK05Zn
ug4pDLgIHcCCDY3UOZrLByjK+EI+PqXMjy/J0nUde2wtXDFtUMOAJmdoPbXK+sdy
2vNav+DxhMRazljbGRT11KG8xYSnDQ9KviSH6DV4dUlSHXOc1+8/B4x4qkF42Bbl
cHr4kJu5RlNML/vCYmixB6g2rQ83nbOG9G2kxfb9kg6i58Hglxq7D5qVp+ZLXou4
vPK1/bOC4dex5R2Me9n3DooZQM5RmQEVDwIZsBPHOWqmiVPQbOcO5bWrAnonMB7e
njVIAa1HFjxF/BKEfsDxjzphcJ1UmJdtW6JVd79l7mvfDggxOupAHEErNNb9Dtbu
uUmZi18rRCUBVAmVqGFBDIwueSWFcrU2iwvbu6Ue1PsryVoGcREraFsfapJLwqoX
2Ql1Xze+7JIVAACt1zBorNwvSyeJZ7QZqRxWSaHeEnIStAyzndoJC9gJVfytLZgt
LfHsHB+9XUE1GO6os27gxMcSRM9ncTvRAzZYtIcIisr3J7gFPmHs0AmqUYQE07wM
bVXmUSaNQzrUhU7pnOhO5VJvxwLbQup1jK+vg9Mx82NmNgtTdxukdmgNAgI3Uwa5
B5Cobf4u2lGxCH5rzYmH1Sz6Y+iyrlaI1qkGfveZRk1glr3iPLk5bJfreX8iAXVz
+6cp/YsUNoR/gvoUuHN9OZxOaPftCakLQKS8LeUjwezgszR/WaFQ75wrna5hGs39
d1zcVjzXXfiquBC/jANM2fJlNJyMwUykh1zYmJgamZ8uZo5CFBEX53RtYbusH0G6
EqknrrshllfPl0sciQQz1G3kOe9IJWNCLO2a77MKlY22lV8LaOcRlEjFkdNwCHI9
OPT3LfBWIg70cxmRWYgHrF5FiKFka/aIFKFk2azNafGIEcBG57JaAZDCx6fMs8n3
sbx+3InmchhJ9I0dRv/dvX3K2mt0XRIzTbq3eYTsZQpRt7uXRbGwJHfHRY2zzbMq
orzgASJEFv2m+hNncHtf8rhDUnlHf3z9F35Q9UtCWSm/R8x5VNqXaMPFAMfGfkiT
H15q0otepIdyGta6GAkzAh5N5S5zO/6cYwCEzppaxCxHzXOOx1sKD5XL0PPI3V8W
M2xIO0xFrEhMZ8BvT16dVrbDstWVKY2aFGIQpClbw8jFktYK32OFaZ3sE6VFeQJZ
jt9py3lsdRY+bQ0/8tP35vhxHotFkl9IwB1xZDDavgC9OwQoczHW8zxPmS16KYwP
mRIMErB6FgrBqWVdH4+j8E7kIsdFRkuBJwtE8Swh83UyPVf2JOfpgXKt9r05fwiv
5Vc3QXixQIlAHZV2N9h9BAvhO/g7dL5jan78N2Xp0EMbpCudvVUjAuJFArIkGp7u
uk5QzR2P57GMUSnPNxM4nEPAI+2R5/vCEMKcBUIx8MKZS0Pxqg4CsFwRToGFxsR5
2jVF6Yd2ERYT4mAr7eVcy3ONIHCqNWz1ZUyVQPGzNVRV7vWlbygVaiIsBrS1l7f1
Zb3j+KciPutj4I47Dgi452oZOJQCMN7obrtCENMVd4x/xZGSa9uCouoIHA96mLx4
AQYUZHAx8ALJA6pAFLwfXbvgavxSPB3yHQsWg+CMMujWOtx5dgT9KuiJbPvy4Zo0
xN1KQdvqDtiIi/85E1dGibKU3q6FIdlE3Qp4qgUa30XTyzts1RpZAKwP44Hr5Zp5
V4b3vaoS0xdlG16+Ouf/6SapICflUw8yRG8Ev1GVsthRbOyLFph3AOyo2oZV4zjL
oCLln3fc0ttGFFBXCsEF94AnZ+jzZ2i7+rZOCOJwo8wvuISqCMAqThlMm40fYgBq
G+w1AcTcDECAd0tD80Cy5oy87OWIaoJgY4M9xZG/oM9zNsX56hWhEa56x967zpAm
2+csUlTQTPfpcgDNw5NuviJNfB7AxJd0ghEB44PT6X913B5LRb3dcafyWc1V4Uau
UPkuV52zPGuBbe8aNPVMf2Ne9m51wVaF/ksDwwesVLuKvS4XUjGVIQPLAx9kCVCV
JbgaYYFdelm28vJRKxkFJhARqgeDzrYaMgRUoBWD+E773LVNEvzXR9WWEq/eJ1KB
tJ5Nuni7qK/yZrpH3poTWYX8XBM3096jScQNSPs2Lm2hYJdvGBf3jfb7GVCBGJl8
YkAfCUCDAn/HJBI28ilFnlSf0d0ux4Xc6HFLSZqXjU5EBOXftUo//heHbpGEOg8Q
vqQugikWdYlDEbtLDLGqdfju53tmhTaeCHZhl1w4Qrh4sXrsLumeT8cRuCE1SxOY
OttNRaLYELrMjft3MkFpjn7f2oyJQevHXSyimSj7q37T28HLOLsjjHY1fvh1p6GQ
eBPJ/615BWsGgUWhnsuE49uTrOsxJqjNYQq3a8UZOdpoBTExJ09Gbo+P7GPKaJr+
q9b8IJo428NfHemSNZGkK7/cMTk180L7IWSuEO+gqRtJ6cukPMxgNUntDLtrJgvs
+TB+XeyIGgJs1yeikniqkQql83Hreh66RfwgjNS/as8SKUujdd/Cx9UMp7yjMjkK
1/ufzAeqv3R3yg7VhwJvH9HLC7nS7uhPyPtAuDd6uLjSqNnuJh8VreMiHUsNLJn1
zAoIOUMvOC9mBsr+Ck98criuiZ1WPplO+x4ZNZOYo8rmZktYCAe3BVUG//cbG2d9
NMos7UK4OwJh8Lcblvn60WVbxMC1MIqIAo/VFLcn+DRoNhzXP/PDB+PKDDa8QRx/
A1t4j4VQse32SBBP8dgeJmzCYa73FjyZNQwlZnpiFWNc8UjmjjpB/+OUSZEkRcIH
ZBUb/tlVi6brK7fhO+FEnRe6IINNqrYtzgNA7GaB+rjs6Yu0Z3q88j2GC+D6iFeW
DFwaSyzCSiEJ3AA0uYwKyoVd27UnnWxbA7NbN9VbAzASo75RJXQiXa9tNqg3hHkr
uA64WYSOuYNme78Jhs19EiCKYvjVu+TMrDZFDB6imTsjaNEXIebfz3GpIF/u0pG8
DkVZDSPwgOPrjsiv1aURuE9qZVFQ1+nUQK5FY/B/GS93aqZl12/ENQbxqcbu9g+Z
LB1rtCE6ufZf1HUwdt4EqThirH1HB1SZjXpBMlUD+GzTCuUsoxo6V5kVu6k68Xed
/1GHAAsDBRyhaSvdDwdMEoZC50jo9CFZ5UtLqCwawasdgTrPctvIX9wpFokZ64DL
6fnzZzBM6I7WeazOzVmjXuVpozXiALupojz0raX8S8Of+yMNIlxfPkACLkcRXO3B
tWWrXZQ8f5GAz3I2Wi5zvnptO/jmHGTuBVPDin8Su4d6ZSqTMv+0uvvSOYjotOA7
ukFFFKaOSI6SwMDACQYqTij9ICTLUc2ZL20lKJ/KZhxKRVU7QAwqgJfeR3jzcV/B
YXaeSRF6pf/snR2oDDGBJafc+iEMBKaCdsmCeQWoeF29O+LDMb6jGmh0aKOWSomi
/92P+hTr296Ss6f0B3Xb0SOC515IfopKOohV8kUi2PnwNqfQYB0Sppd6mlkVe1ve
lqYSQOo66HfZuwdiEwtNdTQr1xx2ouZMsWHR4nydaOKB0j24lwIkiKkG1x8VFlvF
xR6nSWFnxfRZ+/yTRfB+2URZGCsPUy+h6zmbv48kdrUYKkgl5/RsMle9f5LwevPJ
z4kMw+RBeWCIRs8x3yNKHTNBe7tEU1bsW3aOjzMrfjvTHd8UUH7ZWRyEqx1qXRZF
i8Ij+vrruUWtehBHokE/9/TuaaXaVXyxyOwgc3iDyqcyYg6o5mqsGZ9RpyB5Ux1w
905sh4Ke66apNdlHUhuIXop4WcPU0mKQi2z1s0pHALJJg4d2r4E2vorrWSK24bOo
Frlb45HRL3Db+B4rkCgi68m46/3/rlJVuaExtfkh6J9yFdAM630+VuTo9o8K0kaX
DTGAtde5nFP9CzC4Lx5ZrQvk1OBV1F12k7wkcZ7ccoFJaOdrLsNnHXdm7fxxx61/
jMFXdm9SQZKuLcrv0En5sCywO1XHUYcxLbO3e2XxpkUBSpmTFdynoQqG4+jTzeJm
/VaRezLhMAjdOdy91CAMXCuKJ6KuhLu9UvhQ5qW59uRcWD0BkYmmalZRdkH5EI9C
yFE6vUc2F8W1kMeV6TElVQcGGyRGuJquGMoW6EwvBVO6UIZoKjSbAjv6Gb26HSQh
k+9NLw3u4DxntcjtsepCQVQuYQt3fR31WDWScHkLzmnKdf6OJfLtRTZ5+UGOO94H
nRotUmOaVoIvPRI8obUze3yUQCymOlYkCSQsyFXeaTCFMrZi2eeaz06z10qm3dxF
QFH+SNqsoMOD6Nn7TDThBf3TKDnlC4EdAVK87Zv0m6w6HDki2AI5S9MRETANOiKt
KhUvcwvcArCZywZExZm5Bmx46497SYEd30mj4tazUdlobe1SCahkDM29i1Q9dLyd
fQ8Fej+eIgaWCPJNz70r3Zx5dRBLkDnGTEdXyM6LZd84koFelDaO8yMDs94KCUvz
Zqsn61+PT3MHfhdl3LMzEnX+po1NQFIVbFkkQdA0gZ7PZ5x5N6aIavFLG0JXNCRn
mRauwns5IN9SqI7WFbV11aW2Vl/GD9Z7K62Bx++qt+7s9/uB6SwNYBzBLr4xPzhv
VdYIOaH4UGeLXox0A4TQO5nGJHmj3kUqiZG/289lWWxo45LjPLImtFuXEv0apjR7
KuXTLWvfp7bMwzbaYm9LaAVafTn0fw2EolRfvjtwUuS0sgDipRHfIxESqFyRX8Mv
44ynK/qZCX0fDO5OyCm9+RgrLTqplYTBf1s7FZGbpcRYJoixbAifrGnR9q5u5gl7
hBdNDIo048b93MbA76f4NMOhbA+ryGbX1pwUzrifpJ/jghGDtdnBqJIUGGWCz0IQ
kP0MUKzdqxbQBSmmRLo0D+OY2wn1OgnqQif7U2DqWyuFg2hRqbxXrUpcQXy0/TN4
torEneaCeb2WU9jKxpAxEursMfyy5MYeUg4/cAWXi0hau0HDj/qNItfL08LY6twO
ktqMex97sSJjpG10iXUN2g3OZ65JJBCGqKbCeQYr1ftW55XT5kEPxNojP4APN2aw
eG3Tz1TDxXUWDVjczyu0BqKNp83GKA/2hOxaPp/3GTlPSiHZSX5F6Y+LykJ6YjTf
BiqvQNPoYAf22cke4giw1m3KQEGypTNGyLKDf0XAFKUMgt+5kfE7HDvrBB/uX6U8
q6nJIAHzRoz6d2K0vLQ2J1daHu1EsXmRCBtb3BDooTuNR3+H3Y57h0gJuhX/AZju
A4EpMaB7VQJX576NOO3tANwf5JfwBZpqquB75bbAt5cy0jzYwF5iMR1QjOp5TSOe
R8XIsJOqBn08MpffpGeq4dkw7/ZO5JSWOFLxoCHvgAokXBnz/aYD9UAGrerQmdKP
LCFKxQ2v5EjwpBGMxt5S1TSnCYjpme10ppz4xjcsuG/l2868ibnHsjmf/WzMzDGr
SfjntXeE4qQMgVR9ogdUF8c1kzxM657xdsV0+zKDWNE9b/vyLFfnVj5kuF70wuup
5iai9YaX/VYu6vOzOfgn82zPPagz2dyHVnPiYqWfBJfJI93enJgvLjc/QGTXXnLu
pLmEQ5TSZ73QxoSp1ISr18CahLsoQUSADraKaIi3K6iSnXSFlCwU2ENi7cF2waZ+
j8FpR4OlGxZNIl65GYJJJ/R4BbxjMjx2S6FxW1KTuRFuGfQ9Df99wxMUt/Y2ZFAT
I9hrRKlSAKkosax1tnF2wqMF/8RpVmYtrhHw6bhXUaxHJvFZtbKQY8qsK6Ifysgk
Vn3THXHrOjI510QzffWEivLAWzQPLgz0OXxVFbn8GbMXfeqa6vbEzG3u3jbo25ft
e96PQ+IjMrX17dwPlCkT37k30cb1OY/f/wX1W6x3UyPjIKkGxzq8tbO1AdYOemKF
IJW+sTUvvLebhBw0NaYmyAv8CRCfrz1CvCb3gkclc/mZJ8XuSwED4LYwHsbIlsgZ
L+nDY5UzopXdXHCenjMa/PK2nXXIRL1UXVnHDGOvXnV/PmQnNJ3/3xg7W5kso2SP
qUzX2O3DhIm9r5JUWbAUQ8vu98q8kj7P0ja4IuTbmnpqgoDV1IvKJTk1pErbzAcb
7T4SoXHO/6aAHrz4ZIkhlNQnGseA8Y5DJctP+lBp9HLb9ajHld8/hTdcghbefBG2
xqRGXvREn2XD7UBR4+iN3FFmE5UgBSrBiOf7sCWW5Oq4vNdanCb6ZL0dFPVavnL0
Mwixj9IKPBGlG5GhiVED1XClk3t5keWB8PKkr8qpAN79xdrW/0HoLblb3X6VD8T8
jTsjCLBxplfhn+Ko1Kyf+0Pqj8XP2qu+vBLK7yFYDDkYGaDszHzA8yHqyiodYUEB
fhaZ7UGxDY7t03rVAzkhFvDSRW5Ncd7GWLpT6yiRoibb51eXF1QINYgbyFVuWxNA
YXEVw6rYqRTp8f5I2wQqvlMugRejgCX5Aqt8oDYQxvffXAhVJOGDzV0x/0X6tYwh
zuxeI4QtAFE78+msi38Mg1yJdKTBWHvMFWo7gE6hFuMA3ntJqMH0p2shxxii4zBq
EY+FSJcEFMsdzGNUiS5X0VowfZBP52WuPpRtpxflEAnUPlBTS5uS/nI/GysPmTaB
o5G35geEThodbuylABNIK9bNBVWi9W6OJoS/JMD7G3N9X9hY9xRtVcNzFt00Leny
csOPGkKabFiTAZp5jRdGio1e76PdlHqSvlbRvGrXUsQTwzgnodTRawacBlrvVoLN
fp0CB1tWtkozU+16PoZdtRM7T8wxF/266538Z5HkddTzLTsZof4xDwuSq7G3NafK
z3s4zteZBQ6t5t89qt2CBcF0TEBwLNRPXNUzVvs8jlK7+nQMssz3y164DMlrNsCu
s7DRCnPOCZSzqnR6NFbfGVz7MFlZSs1GBnDhWUgOi4kgY1j4bh6qwv4hhOOs7Ctc
V8ajvvltWuMR8A6JZc183JLGPXfjnzTQxVoDLuLPd+50Qis7kWsJecYpaRCrTGhJ
GVllE5sUmL5L6u8Xskn3vOiCB0rkQzwvulb87u5GGRD7cEweioBrjkO+Bf+IiYcV
6Dk9I+g6fhlDCrEtKKig7GLcE5UoQq4SAAVDCH6MkKTXf/2bdlqc3Q8sqOxF4OEk
cXroYSCJFlElQ3UpumCIdYbvUm4Rox1FsgxzTI4YoBBopUwbYpTe27E6wt8qcxVq
BHNQAD2WIt+mkV+0flH0qFrji62nN51jU7dzuPh3cjV7G21aRn42MOU6GOCXpLdE
wZUVRAJwyhT0Sf40IrgWwfLs1VeTe+6QF8D581WCuhBXFeRTcssRylf+IBJnI6eV
mUcX5MSKvuDBhVsDPQL1yItn5s4ycGhzAB+iqpfowV90o/YAH5toQJO6FFo7UrB2
yoRkc4LwgRwc90sHV4jzmZZSZUlXnwzR/VqYd6rbiR2i0FIs09TljGOBg2K6gYQ7
oa0cMfPmj1XfJF3l/90Bbi+9gh38NRFbM/BlouKYe6dFX5yBn8rgxmclOQ4ApG52
dWMV9a11V/0eCPZtut9CXxAwJ6zwIS/pJimTsOCQ1PyxIxQsh5m/mXDBC2TP+Gpn
Ol9Zh00mkFYKYyC5Km8OOunXN67uNWdsqqlcGMa6zByk3bBPVHbmOf+fqC41kmAO
A1Z9b/r3fmmsrx5LQO95Tme/UOMfNeFHxsC1mUHX9w1JVVGcjl1W+mf/dGHxCtwm
mDmct3vQmn7stWtdIAIMyA8dKU33eVEIzRAIc2/8jDta8txwmKpZWsdmVo+t9rlS
w1d7kayKzPvhpAZjxUpLJ0nlkglZtmTyZeQbO2xA1eoA1Bxx+IKg/30cz2T1OLXW
cQEyPKFItlAKQ2opN86ZegA0AfT8beSz8VoyGTzy/9TBi+OHuBIJD2+UzbLQE918
ZbcSrGIraV1FbEZSYRTYQhsk4cA9Fw17dbldnJJ+RpcMnKX/MxLgaFBcAuQkJzkC
gzpbAg/62OTkkgM7zJiUEdBIHyfmhWqaRtMqnZLgHSefJSldUiSU/xfoYS6W/376
v2ctn2audCeu61CzJC5pmD8sEsVlTuiZIq8J39+/f/9zm830SWBW5ib3wR5B00bV
VrfAKQWGgZOE4TrkJjjwRzCxpG34Eav7eveas47m2nQ7J6oJS4W8Sc7glepHmlRd
JEg8TmanETGV651dD8TJsrrj1LErth+2m+2zn9Ge9wDoKtvVwcCMngeOr1DrsOku
f4XfmfdSiY7F7qc/gr/Jbf52fVqVBXBp9omW9u1OLOVzGyvc5hCpTQCuHR1Pkxc6
o0TWv/ymIjNIdC6juHiU/bE/fne9hCkfFMecQvr/jUyc4HYqHVAR0UYHiz/uxtCR
J/3I2I1aqUY6UBcc43MjCFYyxVCJnOcu1to5F82XtCYRDDBN29B8HZAYwXp9P5Z/
vK1bHkAFfGd51fpWcp1IdnQmovcD2vMjkaMWfbmwmr0bkFyq6WP1EEvWuME6fUUE
0hRXtlOmnocWJxR+jZplyJPydr9pOvZqxIhs9R3D6X/SBggRTo/C8A9r8obrWn3G
VuQdnSvTwletMAeOdzNChiMDK4xL0x/metDUei4KdE0VxSTK91cIjK3KJCimTuFI
LQ9z+i9FuwhK/MWyBJBua74MKjRUGI/MUdsxPrtWxvfSGbH3QANWrd59Xi9+dveo
7i77KATeveJJi0oX8DzOthYMbaMKdpjPN19b2irjnVYOpNr1k7wHRvESCQ+8eeVZ
am2N7Qb06fOtiFlYfJjsESYhWlX2x2fJBibWIrV9b8faqqLTks5lhclXJcyd9Rlm
xqHOB7UU+L9ry5+H9HKedvR1o7kZgsAW8VXSWDdyLfdkKV8A/FfOjGRx5/ggxyN9
Mj1+amjdDTjG77whfzltPNnIiP8STilW90aPaCOAfhIeKnPSOVUXng/RUVGl51xd
YuvVN3Gi+pzinZBV+iCa2yeLMPIuNUASLmSaKkwhvvzHaMM+g7+sHcGyGzDvZ7xJ
jfAft5s5lFMkTShZ18GkUe48Pm/LTBHzazLv4ve2LU5ytGi7AW0b3ItsmpEeXwNx
sHLnrP79EnFkw/L60Kq9DouaebLPAE50x1mF9rzMmx0o9wNCtdDJgQiiYfgY18yR
7AEgmi7AcK9lUFejNKc9oZ5p9DhJlZE2aBQL37uBING22AgiMjRo50KqIOtPJutK
mLg4Cwx2Zf8Fa1NZtoMiSp59BUk4T7yc3e+HpNjtYQZdX2cRZG9JH84SPuNXur4n
t6n3k9nOCmP8zwVrVDK88WbCCGM7RXdImbBqHfFLKSPFh1BRpzrdFKQdAruDWIkD
kPEeCk1W4K+gYt7Zd7GOL+1meKWlHum1O/eV+q92Uf7vaxeHHVJlxYUIPxBUPtkV
drzh2xrRgYeIJq9fRx/uw+WOHDWwqwOjZlpZIdjeuY6tZSw7Ofgcq6wmGjaUYd4Z
V9UKFz0T4h9Jk7iO5y6duH+baXffx1zpiDusXTthTa5kly0+AzvyFY4eAVonikZr
a8l/wVI7eYFFxGQSlmzmvu0tHkNFF2q/GgIkDhiCqF3ib1RulVj3i/8rvUc0j3hI
NGlAOEoypkAgae6vmfyHTkOL6CVEQ17NaxZX0MqX8fCITbLAYYMC0+ezFzbzWL6h
qCub0FAcWCQUvh36enyuAl0NY0ejrcZuaxDae7FQsb6sVBBtQQ0YLRPdRhs2EIw3
YTwb0l6WOITyms4htuqXXJxYy96MKVKm1HNA3a4L90ONHCea1s2Wy7T7KYgjGQFE
AaEeQp+k6xcq75+8wgUZ82vu8l7f1qdd2skrobW0INDLVqpdy1KyZb3LiYra6z5H
zX5+B+1KeHGaku7OF7OslSFEbEDy4ktdryp2MNnJ7//EBGL3WQ601G10VPiPhR8Z
DJSYZY9Rfz32kawived658T1kO/oOipTP6BNq+IX4ZXXAj0RDxd5kUE8qi67tKjV
m3D77ITU1bgYDyO8QhXlshOzkFXzjmxmKaZufmAIREQEEddjSycJSHFramK4KjUI
ICwdBHNsmpYILhMhgJdKmREGLREj9QLtwtGDV/VTEKeJbZ0cUh/hzsgXwsabNhrw
jErseVEA0MmRZ0qTTvCtSJ8BeNUdb6FZQHf2T3sR22zTdTDfY8Sfq3Atdb5i4+kC
vR6waOo1wInZDZ0JM0DzVtfM7V6dqeAIaLIcH8lnL4UEJ49jCoq6MtfIjwU/YKsS
v4H2LJ1phZHFighLFqlEP8t9ct3UK/2ePABOFUW2vRHrUzzH1rIlBZZqFPuQT6jV
+MVySkgwbJv2Ak+DRNIIJ+pv4T3rzuxT5ARsaQ/xuuxyO/sEZkeIk5Ib54jTowMD
NciyD5dwpgd6tYMVvoFUQi4Op/Yea2EBZTlUMGlTCxwBIO9mKJES3VrnoJGzU5bX
MAVDjkwvLaQc9DEXKUOaz0FCmXFYur5C+Rbz9/T2J9VZAmRpZxKPmYoL3Pk7SC5f
rv89fgHLEHk2x6nuegGKTiW5U7cXYzJieavdUK+5NktiyH/ACu4teh1yZhrTBV1R
GBbBL6uKX2erzlNNYXnJXMPmzLSQ42h4IXcr2mpjxSctI74eN1Y/lOvR3ee5iKZD
5vDxA19UuJAnMYM5gbpiMMJb8/zdjVEm/9/UNz661Z5lU8xW7a5iijQTlHnO1R4h
sppQGnB9+cz+K7Li2Vul0d6UYrcHK1kklvfH6NFrT2INqdqBTF5TA3+quspcx10G
6oYPqxfNZtoqlxXZSBdeobScQh489EdW5Zs8IKo+fUO+5hB632FreRTDmQlabvm1
i94vcMIOj17LeTmrVSIKlQxW753Mcsioh0cgtye9sEyA/EdwAU4PlquyurEXl3UK
sdUTaBLqcCuPZ5dOjvC+yOECiQGpCy7j1c7yMkWV6xSfgqenbQapqsO4vlY/N3nG
hvcoI+/rXAqE/+EASswvBVjQkTmhRanB+u0C2IXx19hBrhHGUYJRBUOyw39zFLP8
MjnspgJGQKYtp/iUZocNUi47x6CcTXmq+MxA44UUBwRWHt7+uvXasTPVd+YF014l
NJ+TAAX4HVUok+1PQ6pek2Hem7o0fwuZw1/Ln6j8h0LJeqWVLw7ayApuHRhZurey
Bxq6aq380YITxnhxU4LCCKBd9kkNRgDEvzzDSfKwLEbYJOHZXs/N0WYjZNHXf5u0
/T5r2kZkA0Oz3Z4rq91TvtrdrxWohj7m8dHk3OneKWEHFUI3/iUtfA9cLtaCyvkO
+nyBVTYlS93bMn1qTsVrm5dtPV9FAHKeEZLViIjM/9G/sZ1xEbYEM6YQsn4lv86M
SKMxVG2fmqo+CmWu9xkimx25j/HpnssSvQyvtyEUpCFlB4hMs/wV4lJgOUaQevVO
NOWND+GrPquVtBGcOTSexPyAOkKGP/oBwTKAsg5MKsSXHHTiLjIvbyY0arqaZTmY
ajVKmJRL0onzvi/v7f6JJIpWS3vrnGf/UrIHZ4eK1z6/bqi7D3byKe2c50PUozCX
oYeIATGrURQG6fTyZZcZwYmzsAOgDeeJovmffkq7VDv7zGd1tZeqCAgMmNWXVL1w
4OgCxsdewOOWIJQ1Z1SMf7O7A2AC+Iny9NjC/xaaOdfzBIOpn7VgMy0rqm4R5WnG
ZnraNK630EyMi5CrgbSUF/rrfDkUKneFiOjaHOdgim3jILLvWpG5/HY6pUzyGVpR
dQNL/9fKO47KherMBI3GaQM9KuC3kjMCPXxiXh0haXvLw0vKBwPAp6CHfIrUPER4
SzBXrrnGz4BervXq4aH/6HEf022TYHYukX94VzCtJ1vO55dLb+D0LP1aWQQf+h34
iadqXsQdljYTZN5/orJqoWMYLSj5aAjL2gqBbaICwBo9mtCxTPqAt8WB/j/nG75K
nBiITD8Ob3I/vZ1pbM1sbLkOR6M1BoLsdD6yb9E1G6ILvfOI5VGr17OR+vzTVg9v
G46jqmjAFnE2NF/SBF8oT2GT9rf+eTQlhmt5VC17z+5nQEnPKVkcLtGP75T/Nfm9
++hAYtBQpBGttRAFaUUzcv/3Ph7W68UBbOG6hXGIfKMG5wYjtaj1YuKjNMTrvHIo
7K+Qm4JHbrisEFW7Smau0fTrShfjk81+txr+g770fPPCHBbD7kRfAWDmwYnDsV4m
ri06xGlEGDVMaZ5APl91TtcZKifWJSr7JfvGt6U0lztnBjt4p2+FFijFfqVakPym
mVOKy4hKJYzznkkI/fMI+PKUudoe2nax7he+b7XqAPekmeC5PqwmGSTpHo3ZoyZw
8LltfBZ8FdLVfOl7WFcOP8CO6cCA1n8wpXOAuPMPFAKbh+f1xgUa7rUNThYw1ViM
I9iLzQJYxiJQn6eCXWGJw7rYvNci0+y4HjdXs6rArXOI3lXXUiGAOQGj16JYfPkC
O/bd9JX/TQnRZz6xzFW7oUqtRGgo9KTdkxLKb7yzhqQ3g+VXsd+PrEgcfuJWPu6E
8FORo8K/kHSvOUwhgGIna9JigIYzuMlt3MIdaC5noYlp46S0DA+fwCr4gycPRPd6
CzNfrdVeHyf6ZiSseUusFLQPbXj7KgUgegj7Dlw3AeTnSK1aBSsai9N+Y770M8xR
ZNFrA2JwkwhF8r5auR5oaNVYwG+/Cn0RBbQ2uo7S8PDECpNexnC9z1/jqL5GjjkF
CjK4yajSqsnMBYEaBsYinFfEtrmlFSN4DU/HahUFMAL/MXVHMhBFFZZxmMBMPaeJ
pStBkmUPaHKCtLN9/T9xXAgjBFqTXjbs/IB8i+aUzYu+i1CHBwY+5ljorG9PjDBn
nfurqm0OX8fn5MYdZabNuXVocBP+svqTkInebBjNxHA92HhBp+2YMX8zzGAaMMoj
Ruvhhi/o9YACPeWN08B1tHtCFTpjM4ubNg/fBEua0qjK3p83FsPhVoA83JFj7lqR
QK01VB3rPfXml4/HRqhVcbZYdht/Jh4c0YsIcOQA8jlZqaHgTBOPiCmcC/2HKiBy
htzZk0g+6XPotAPUk8QlwGetqC/cDr8nOmVeabIXZnQ4uG14bztOxpGHQueq1ajF
3yFBYUkJt0YYWAaBKQgHKszcs8McmVRfQU7w53GnK4nsGhTI9Ri1H69M870er6g6
8JriS/yQ/gcF4kAl3YxxvPUPLHaDxf1971/X6z31875xH5PjEvyfgSEFP9ayGTQD
z5gLv53N4aKclf+VfnzPjZANO2BP3GC5CfOWxJiy8LCP1DfoT2BnTGQtfHQ5lj8C
WTK1VYnjiP9Rd3bPOFnTXuZrDQY4sQsedXD+Xpr/QE3epqoLVhoSiiz/IOlvhH32
78F27wZWF1xUcWFWaWrGa+RnK2quM5XSsHGCxG3rtmZ+LiEhlXHFVkUyrUtkObug
7sE6Wk4lH6brXwNSTp/ByKfz8zynOr3vUaHivehnjAcgTj17yQX8xEvZV1TxwMgO
i0387lLb97y0CdlnsLaKNnHXVtPzzn84/pN0rdyQJEPzdMVQabqQmCCRAB8K+Bat
2RfQr/P+sf/zfh70xJoQPXTCOL3WHc9ms5+nn3rOOES2CVFyLIKfGcf/1Fs2ZDYL
T3waNpb+vPHa1e04ow/CGX/Ubzca0H5r00E2a5dk+WOvZoLxCJ2vKfbTm/qrn1/M
SOrELczEld7Rmv3z+9dc7ZT/3TsMgxzwAdyds6eNwcrRZh0wvAJcchZR5ajQjZYM
eHxoPM8vsPXUsYCOeXG+mz9KXZBaxXJa3Bu0LOC+bsQs7bqKkFBgP6dpTqQCJBsJ
3qvGGJVWttzVj6fJwpGFkVLFlhCGd6/7lZWNzTBf6Uvg7zYahM8IBbK2hfXanGJl
D6R0hPXsE5Xaa3bZtfg48mz8Y3RYbslTQh4ZMGIaMWu8/2Ne/iIeCkpOf4LOELEu
WXaZeb6CEq3odTk6uuKiZJ6M53z/DY0369kYYL02bSfmIxqJN3agif2toy5eh8rR
gbGvWKF7MzciriUDEtcCY5h8q2i52Bd7ZM8oswhxVnuCetQO+2s16c20i7K1423X
FFq7oGgbwWBbi1cFTZ27NEq0l6QlF+w9iV8pXs2hgM4moXZZ6uwev2Mkz+lwYk6g
ehQGI4LBxv1d+YA3IOCcXOhsjZJnMsXPRYzwoODrnOoBkd1dATHNwHYvkGDxGMWq
fmejgKp8tXgOClyJn+TSRCqqm+ZMt1A8M7G0QZbpb1GYqifQ7LRgRiTm89z3HvSW
2JHplRXThGlzsmV/gkbJIB7aKO483hAe5Xfz05VlAYWSzyju8j617f2KS2GTcneQ
1DRGBwTbLUd7c+Smq8YkmX9PJIKIA09lBkoLnP3gf2bbEvRuzaigOa9s74WuC50w
SeNy2rU6YoOrDWrhfMxFII9XFGZ2rdPQcAh4QsExr2ZAy0ds9K6adjq94tmpARLE
eJLNrJQLd4LAK2MR1J/EzMrmldNzajQ9O/j1ckWxSz98ELtxBqS/GcHJF2RxIDVy
J1Sa+Y8PF/cfBiVpSNhRMrP7VhnKBMlhaQeUUDGsniRNms5BXhAtuCL0kSemvaL8
y0qdKvNuUd9Q/ES3xWKde8gDCVnJLIRafLCoyJHb8N1jKrP+vOoLJDfUKovGWkea
WLQeIMQnj6j0w3kWyBRvTLp/NDOB5Q6BjbmOlJgjAoGOZTHM6FHcUrLZmtJ/lOwg
OWmlYTJrfYv+s7ROoojIv+bBbc3/G+6DltCmUpe4D0LjPtsorj3Sca5y491m2JAf
WzXUBgibyDyb8ZKdgInq+FtsPCziUReNYQhzVYKnEnVHezb1+EYDGKARAFjwcqoJ
FyuQ208jWbxKbUCH3tQilLOegZp1z2Hn1HvhSV50MciaeVCi68gb6No+Rp4EPtbh
LYsI06u0KzcL8sQYFcN8+kU5d7vJvBU9vx/Glxn03GguGpD1WoOUQHq4t/4u3WBw
Bql/WnBhHjey2jhx5Jxu6W2vnMrYVXx/8YKJIaDJ+7cShfB5BJhCODJfbgNXrpvx
tKHBWdJilw0q13z268cFYj+vRU1a54T1OQvRR/reVcrgVUvrjCVK4l8A3IO+5qxT
9SlvnbfnQL4K2y8Fgint6jYiaw6QNdCd2V5e82GMbLFcRTUeFMfuJzeEUBTIMiy3
AVJkD0O/BBC6rFxzhSnaprPh1Y6u2GevSwrZ9nhCGA55XSYlvR3MiDcaRgnmIQ2U
DQGx4i2Sx+Eiz7WDtdSPu6C4tSb8Bh7deSC2AGXEZYLgk4/yjsjx7DiJF+6UX9dH
5u99vjJgctPSQm0qvKXd0/7qW9jCXL+R82x1jWu4QWKasg1aqrfmrdpxQqCFy3k1
GQpYyP3WFzTL+Co8CJVtEKjvRtxXNEDOUSOVweUJSOj2oqKjyeDKYdrO2ZSy/SUJ
Fy/de4f6/GxwtcdqQ0f/xaVwT0+6W4TBCOGRYEHlWEp0D8jTLsFSFRDLl0NEPjzA
6i7nbF+I7qA5qImGXlmDqnKlzTOkb08k1smc1Ex/HGLGvOjsYu+sgi/0x9bbnMzM
Jb1KQlqhQglghhX7hLvg7Cop0urtwslXyU3Fyn95RSKsMSLcg6C+XWZNlJ8YrcAd
CuZ1q52L3g/0Ali6NKhLVt7yLA4NFyO1dtedWSdkKBPOg+Jdu9cnJWZnokAM+MuW
ikrpw6jZu0VcjnPaibpUmfvz04pYLDmgnmoBPg1sbN9uTC43X/REUwjv0ZDEmvzZ
pYZA5kJbx9FvDvqFSKx0sjaFdd++xB3+SuEtmjrdnELsyq4u1uYTvZHI9BtZsseH
MFsfwE+tc1RL8pROQ+jDYuJQxrieKyTKOGKq49N9hx0i0YyAosOz1nvo1M8RSfJM
aZZfGbL28lrQ+wuyESIEg/dbFKdHO21AbW5T2Om8mvUpfYUb8UgMSlBBTFXe5iVv
/3hsBQfP1hx8AQ0Ac+ix/mPw1i9OvSLz9klt9tpzjIBz+PrJpbvPr/kR3HOjS7VR
q5hS+J85x0TGENPcdtuC0boQ2n60yzZ5bc/0tpS2Srg5AoNfBwkcMquRd3SSXjlB
L73fC1vYjU3MeEog7eY5U3fdnTRicrKupoib1E0folIu8QBVTt4slb3etFJeNg8f
JsIQ+TQdRPpFoPS86gFRDqrqnoszsNwpHZ8ovvY6LWefu0pdBrdEeDeWdlDPangA
C+luFJGVfxgj4a1086isVTuRRYOZURt0+kSAzcmX2Ps/UTBdgKnxNwpcLEbz8Abd
aWkIwefVdqiNGOPbA9odM1weLrpYfUD41V+2rkVlI18RzH3X5kfrqYi5Fw2b7iVG
+1tN4l+Q/DHHasVqXmlzfitBCDBC8jTayLkXr2gwM5CB7EUNvCrlLl7oscCQ8+DM
tPoVAej7fzjazAD4bJWV5SQYvKCgmff+EbmVjOO8WTGlkyMK7i/qxIGuIqO65m8u
uSzxQhXTrlZcSZL68Dvxbwnrxfg8fhY58pTu132xxCHhG9QR/1ocXgEhpeAQenJ8
yemyYX50VC4z/cMrefeC8w80gWlqZrT35/UexTJPC0n0cQOoOfX0TdHpDXloDMAM
2G9FnytpGGWwLOOwTqauzC3SxBQKC1Bm9H405MmNkkThe30nl9dSAVWbKYxRMaAg
XEX5s42joEMHxUPV1OHbuzNPyAjWuVtG8+NO2FrkmuB0c2XJ/eTL2SWlVy+VWMGZ
D9g+tnHepjHg+5eLx/EjNA3lVkNsWwdo/Da4pGmhTArwoxFcSPiBOcjmQYt7Rbul
SwCeRsRD2zrBeOYHjKEcxOwgV7lCx1QCps7cB08M2bKuCvfQIgN2ELSQrMyJdQUW
ZhKysfzNdNhRkmLxYSA4aayRLUqXL4qd/SayNPrmrjsbroa8L3QEiS+Gr6TIKMPT
nMT5ze5iojcL5N7imA4AptBGIqrWd1gQ2/AaIekCSpOBpIHZjf4SOHgTbizVVSWG
FZJdq+wOQpUQsCnQGvFKnI0e/HhXQeDrfmSzLZmVx2H8vKtjfsILNMd/GIRFEbPX
GavqXVmmEhuFgB/BDY+JJ8GW3c27rMEo1Cpjwom0yfJDFxZMuF5k7tE2b0zIwKiW
HIdHFrOJV6n6tqCt8Ahn0jGb39oP05Qz7MzIa5tJUDZS5+rpTN9o9IuGIm0VFmo0
CA8MphwRS2JZ7Ic5RZyydWr/Uu9peKxkIpE9gjf2lrSlNpIiwUQCYQV4BaJx/XXu
J6fHA6EczZirBt5tF+J7cFID+elucteqR6N/vaEasabo3GnFuXoOaVcmGVgvN/ws
fn2754jKcIznesFdjwIBxw3tINhjCF59s2Qyuyf4FzyCE36sZ6fgd8h+sRsIZpiP
Hgx8wTJ7H9M7AwB9uZq0CTqVMf4Y0fGd9fxIT7+uEuWA4ThojLYOj4PDDvPqwZ9W
SUUZjYOoLigetfj0Tk2UEibC1vYIwUPufEIUKkB53fXp4LE5JRw85snubOzZe0Ls
V/Z4qTF4pc8Xmo+70gAxpsZZ9itm/Hc0tvcoP2qIHUG1Y+bVMTHz22YkcvffD9BG
8/PeYrE7WanSYwjNQbPwce8slEmy+zywubvIqDKJ/9YL9rCQ5QfkJzawHBQS0pjN
GaToFmVAFqbol0GycrHTB8fjCTt0KcrTEs+yjal+4dgZDUXUHJK9X6qjpOlsEMZS
dB/CY3xU1siEbYIoqyhOtEkQhPddPHGXUL29+5P9ppgmDYyu4t4BFneSU6GFeeMc
mN2hN3JIflREeuxZ4x/jveEav+GVtnHPSFPbiNRu13RJHiBs4ScAykgEuKFuTOhW
XU/6dHDekOAzt1B0PkEecuKMMdGlssuBaNaYgO2Ujm/nYwV4xJqKkTdGUb6Qx5nh
ujf9IHQrQy2YLIjalabkpTTFinjkBH9lUlxsksG3VhLLhZbM00xdgPKmcLRTzwQj
FmTSKdj1MqMuer1DcFETLib21uZqb9ED6xKybVVdW9VYpZcFryWJ2xaf2LPuqbQk
blrxqtSfzmvviiNal0tylD31sehqQH31XCFe1sB8a1uDOVM0/VFQN/s8XEvFaOfp
UwMvDgtg5dMv/kZKzyFj7hBrIn6i1Ipm+AAMr4aTejeb128uZoqMZ2lIEFS/QiO4
YD+2ZerAd9MJELg6nNr1Xqc+jWvbtAvNVHJtpg+mtM2SGCeYU7VxfzIhhjb8X+1G
K6W6m7h5Zr2Pomkz2g9bT6H2QN49ohD7VLh0aDnuSd/++y5K5lDxL+L8qj46eET5
i5+uBACKE5PfXWHnWm3BxRf0D69N9A9Z7+FChy93BrysRQZUwq8ccnEtt26wyZL4
Ch1MHzJrP37VjTkKyTBQZFJ54sExpTqCVQwuqf1BhPsIJHQuKs2iUhwEQfifjtru
ay8dVZGHl6ezkgxiohktf2CRZ45s/2H8NUW5Mb5ikET7QHQCHR6C3xccxeOs3Bc3
c0Dd1A6X6rFxhVx8NW1gERTgNunCRZqbCdHcyMEngd1qhxpUAda1TCww5LHzG00O
W7ieDWsM2DUPkpM/yxgmsXERTuMa44NRdVB+3SQ82Mx2GYe8PIe2dJ9mcRlBoOyP
aJxXQo3JbnWWVn3GGkAxdQruoGhr7HLXDTklNYP5d2I1Skpzv5H37C/B1LTSFQ3+
Um2hs4YA/z+DpEUXjOrJHM3rPCYwCzc2+Kqz+W6F2jm7RL06HqgZa0S/J3e+c+kV
/As6FlbyIrqtmt4YaVmBHlRnP/rMFv2ZJvA1bjG1lfoH1ZfZo+Ti6Asf6z3J9sBD
3wabsNCjnGT3aBPiQf+CYNT/TBQFHLsoig4Z8jmNrdjLhkQPW7AaJepAtXV1Sr4Z
ka5at62XApdeFJGDK7rp6J7we6BLoHRr5fslk+eAY3uCuDCuNmT8ICr9ewoMy1kq
6jUSBu45BVuCIh0r/Sgc+R17k5/QHfSuZeBVQMyzTbVq0FUMRWpC46xIW4TYDwz5
H95mVGwWvLO7Y1CfZ5Ul3TbpmQdBaw9iZbqORSo6OFY+LiHikrU8AMAf1q/W3i+q
t5OLMjsPfQUlVYFQ7ESeztbcZrDZUxm95RDa2PDUbv3soSyxtXCs+PfrjaebGVHZ
7YWLPFNjqgTcdAEXcZt65I1553+3TcifBk4nvHxTZ3lgPqGCKKX+K4Qxv76hGQvZ
4ySyMO5LHQsOBBUm4s91TJcBlK2EbYSFY2+xFsjtKKao2zRkvHZSbG3xs7l7nRLV
fGoZ1JIuk5afpInx1nPf01R+WeVVi+fwkfv3zAk4XKFgS5fMUkulWbZUY3BgLG4U
+6EMKVd7FHB3QahOX+3odkABeajlsl8bqvMzwmEXQ8Mn4jTCYQ9Vvm2TF39uM4+l
yUlU1VdAc9DDRTIaUMKwP7u1u6qQIvart14ymyjHT/+cyFusa6GYIW+K4tW8UTh+
3l+I/AQeCpyV6DhN4Qb+03J9K5g1cqSO7kuElLLTJr8vbCG+FjM+ACIqDmkopXzg
x5R99rOzGDs4BT9j3s5xHLtxFW5cNxnxqKxrARzmTHXFev3Ty8OFCN/94Z4Q/YlW
sSZVk9ybr2txLzw2oKQYA/UxzVhFwSbDTFZykFGjolu9mXQeM5jbyznOGaIgrlSl
z9f1nTisJwWVrZQLkWB28FKYyjVvrJsCMJHEW1ICQp6SSa4uOky6l2wOArfYxFxe
P65ldMFV1vKTM2qDcRapl/OxwYBKS4N7LPXT9HkwHPXgMoU6dXoxK6CKZoQtH7j/
G8BX86VYdCfx9eITh3pC3GvRn7nn39/l5LKzlR9E57gvo0qBhV3IY1lJYYfndKcA
o81QYHWzROJw596bMOmlXN0VqrK9st+5b1n1m8LYA0d3+o7F+MWo/EA+j8nHdwLV
6pn5Wk/7rQQfnfpdHNJyDZOv6mmc0RIYUVHEvX0yorh1QYL11djk7Fv62GRBVK3q
83fd7zg0MKt3vQBsdkjoc7/kpoGf7lbdCcFyvfzoZ7UDorx4ZMuQW7YvatyG0TxG
oWoFA+4U6t4nApLmDRwKwzlZvwuSjgUVvSBjJeuDaPQjIeSW4qr/FMv7+kFLi94q
jzQDfIjhWg8N2uFCfFFtJKC/8C8FFWCpBOGjielklqyZr8RSxiEsUbvCMA0qvPI1
TfTptK6juzHlVxvjeTvpCDT/5lqLuf1dArLaqZQ2wH4fYfW0cX3+JBUTrWppnAmV
SqZ9nWbCBcM+kzsVopZpTZoUbXylt/u5HdEV6NfNyHxj/eX7O9FkJMxXh+BZhqSQ
I/6+5/xbbUYFx+hOghuLNmcj45ExvdcvjEhloA7cc+4yl9hWWLa2NQT/vjPAkVTr
oGaiuIFB1HoGFjgIFiQFMMbEgI48wN5i3Hfj4S6Gkku1G4zkmbwFBflYUB48C7CI
IQUKXZia+Moss55fi7Yzwx9jHPF9PEFKv5WdnVJe9MOYLIHc8s0JTnY6MBynUqcK
76YRpaCXto6sVGB5ugxBWOc3KTynenhSeWItWb24AhyZ7eJNFwr5LOi1aSTF8O8q
6VNWRGA3ACo/X2z4nJ3YK96VsKTHgPoDoU6+FPwSbN+HZYNt46dADx0UlH8QCM/1
rDXTo+h/EL6QY7Qf5nEGoTLslVPIBYJ9qznJoP9DwPYtE/os/g3zZfNpFcOH3Ga8
9885DBzwsU3qeCHTiSyDgbGdz1UwUAEze6/uHpkwZdTXDfTzxuc6gvlg34PKQiEU
dUC+D1GleP3KsK6vSIHrmYNXk+XBqmcSwm9tQIt+hde/dzQFhcQVoFQ3g3WLrOjq
O9q/ptL8guC0GKSBwbUAOQ3++aWrdNGPboq+RDEH0NhLXeIf18VUr00TN2HEuRRE
oPxifkpwQCvOhmwMIG4a8SafOsauJm4yQSvTBI7rnH7Ou37AOsA+k3+p3cUMknmH
Eh6pEcadRUkWWEzJW8rc/ZBm4rHT4QsWKnTSj6fG6vYTf9pWwBvOn4r7BeePMnGJ
M05b5XUkYFwhGfa2DrJCDl8oVRT5C1jbvtn9GUDyrfhKsHnQWe52ItMjbFjhmNLD
9Gj74FB9lWIuIY1qe/KMoraSa/pOIwZJqfOReS392Mfhxw1b35rOELsceUD47Etl
JTvrhpetSTlfR4fk37hQdzZqReKtFiTXa4Ce2SOHlw7slQfz0pyjr9pPdnj+9xL5
3ZGM+6F+d3sq3vzdklrYfGcSnTSifhCJG2szLjzl1ShDXxQqugO0h9cMkgDkUDL1
Oy82PhKxHy+Bv36XA3g/UXCa1e9AxGcqKHqZg+oOaZe4jgv4N/jSFwQgTkrC7F3J
A5eocWRoOMsHol/LsmmfUr8723H+IjXh3csnYHPbamLS4BdePDi1QmVePCd5iovW
NCcz6bObaDdH4Ghsc1tb1dlesKzLL75HRgYaJ2kjBVezo2Hz4qrr8JiLjECdEkN/
5TTTl+vDMCnZnT/SQAr7Yi+Vvdr8LK9mj8GlFhw1NjUIT2ZcH0asVOq8c0JaHX4Z
hUYs8l0TbPOaULYr7ncKD74N4SstyzLH4APtQhsm2nRxEzOaIAWM0unDLfEwdSI+
Jw1TLdQbUWZ87zCaXKejA+4sUvScYxKCRqp0s2xpiAPtJcCvswpdP60bZJWYZpIs
7mikMPWrvabCG8FgxnJKkvDdS2c8gWmk4NiC2WVl9vhl5S8zwUYheUvnw12hLOYc
M4nPJLmJ44XTsjBR7Yh+8Rv3Y3A5ytPAy1R806nske53POVvO0z6mCN/6wgKVJNh
NuTIe70Js8oY1+NsPdS5v6G1XSVFLU4bo5mFlie21dcdiZdtyT5NbhfO3/MC90N1
Ryak7rSnbfnFQ+lR+GU0DPomN4hMX+pgJ7D5ZNUzeKnBajoTI3xqmK63k+HkBqPq
JhGL7QAvQC2P/KQOa6VMvRuNRvrBdq8jWv9qKGvLfXE39QypalYw+p2qdJuOHxWV
OgFqDUoGRKQyEbMdlZF6J6PxrfAzCx4XCJbN2b9sbvmp3tTU2rOA0/cEP2CLcXek
igV5gwdOG+9z7QT2TxlaSABocy7vP7Bt067OaMB3/KwMLIXM1jWvW6NBHm7DOEmR
mnFA87TPLnTlkyJklmyQFsIA4vxHDd/ar5v4xuWzKssUV9kHcyzP4pDs0fZwI3mc
C9WRmNdQmM3EK3cjrGBqrGCpBDrBqdTNTC+jqZXeX77622H+q+4zBT85HH+3XEeK
tdf6EBKSRMbo+yNWT+xVmEhwobubZfa2SrddrqZ0DMwAwlRfHq7+dOgicKe9cd6W
KVajFPP+L55vSIYqcmRfQ/kfq2OMcDI0jSgcSoZIeBSztrT5c1/TFkUnN3tLNTb1
BeaKxJkgiAgkitTPq6bLEWxWzOFxfr3Hjq+9efiaro0nuqriZX73BcchAE5wxcsR
aRGxRptjIMHMouOCzBbMiHiREgP0ewzyfhYS9iKHIoaoGCeBDGGlL6iptsiUmgcH
gdKRdB7a0k2Z8ViZsrvCNtgdNVAPhyPYkhIlJxskhOEop/iU41lb6qUprXTs4b3c
0BK+6eMdpmo4thpOacuol9ASdQtANH4hH8OIiInPpqUxvXjlvvLN8gwpRe5FVprl
HPS2yhO3hrnaLVXFTz0SxeJg/y0F+cdloy0+lVCz26/MtL95YvcgdZhVlnieWHJ0
HQ2rGW15U2dV8BV26ZZwpWPm8WLuZ1LTyvuk9ROBWOzhoKNu9a4gZDk0AFrRcsga
s2ZBzB/QxpMgdQ9+lBvQSCxgfRQGjj0R5MAf/NetLjilMe8h/dIslXuIRsze9ROD
gepfsfxP9IDWOTc3NErIYXhU/j5dKg3EOiqgkW7zlljx8pLJdinC6Ssyb+8K19M4
CEjfnrMgKomVlINMbFYIPnPTffack1aUJAArYmv+ZIPrsJJB1/jCUX9081cS5vky
3ZPwckSiSzSL7FkUx+j7pRpHsC2f+s1V9uqPJGNBRbBQeGeDGMDS+wMvXXnCvfAi
hAILwI7+a0wJfwr+Teedj9G67CIymJdrKWKxrG684C9a1wa2BdWYAifhCi7Dn+lf
m/mJBSiRJICGcG84CuYitpU0o5VUlkNCwolq3MAQ+/nFj1MYZKRWEmf0KGq2UeGF
txo7alMEzSrLXquOzsWO2WCwG0qBIbWG5dqysR/AFPgqLJOPreYzFG+WhaV0nfZx
NP/ZTdB0tna0iUjqhQXLvgXcuRt7GHfc5orLjp32Yi9ndFkFnvs791XoPnBEdSRx
rL7XnzuWjO6ZpnXDqK8K2AOi8srIaokYRyUaVl2ANf/sI+/ntMpb+BdNPtzY3nI2
Aht3c3pvcfS/sJBQuayEusKlFw1HSqsiXN3s+lJp8yNEQfbp9gH+L3hlQucywXz9
xI35icRy10kpyarYLhcxKpNqtYk2t+CGdNqYgcOnd0IG9RvYqCQPb8KT6nx1crva
W1tEwBXNTh2ggfxmP/mUjAd9Gf7jKMidsMei77XPQC8cE27lErBkzZ9LHs5v1auB
miTHedZHUOgrH5UjCYtVhcYS43rJY2b0ja/BFWdMigUascAVcwzcf28EU+dVXXUH
ZD2lZVD0W2bPuiVZmf3PFZyepurJLoTCyr0FDCfHbF7qVY3O3vf7aO8b/QpSoeS3
zqHekXJLWEF6SqswPgfyGrMoeJTZxn9dQrZYOtDBZjh4JcLwtuAtBsM3rlrvXFLt
tMhsfuMMs3WoY1ar1BaVVD9jBLUTWOxZKTpBFnpwPrQ8L9/ncvUIiEhsP64E9tFv
+LrM7CZLOw/kd82wHJ4s163oHgFgiz1cVIu+zdYW+7cqWMLUA4iRca6X5Jn0CNfh
+WY1qtm+4WRVWaNvBAvdZWE7frJMa3R0z7195/sI23S8uUWGtrvCZ+SaPpdB4gMC
c8BVITOFVHiIk2eFOn4tSoFPrLlt2uMa/zHhIqeu3KzGq61RkpTs0n+9aDx/jySy
+L0MoaGnhBtMLTmrDQN+7JrdMARVoysqNUkYI1c8RCdD20BB3sB28VFw59VPyULW
159wlLxym+cgYJPomSEjsygRjYJdz/qaMgpyJFnG74jSuDsPMjpDvshCVbW9EG9b
fQxtxqCf0DJT3rPNzeMQ9kJK6ApGO4IsEHoGts4st/4XiziNlPSA6Wu4glld79t/
uH473M2csj0mePQIEmARvfvNDmxa+N7LuWdRHH+WjdJISgNb52gdkQPeDNxGUcwM
4LLkDnvggPO5RpJjWn1KHjYV/cQOfayR+QdDK8HNYxI87UyKN9gY8+wwHmbhKm6l
QkRwkTtkaO5T3Nq22WM49Nn04lpBw6cQ6l31TNkW5/kpkesPz/fDXQhrOGKShvfW
I3KVSp7/wYniedmO+7C5QoPRSQoDcbYo3AP6ms3974tA3RgDEZJIPEmjsHhVkjWn
hjPz6VscZJOD/K4bAFaswMF4BXqFi2P8uxO7hyR99278LPnLAsfOALocrnGRV+xu
BM0vuN+xT2PLMV/e5BfWKcOWB3o+P1R9/6mTHrVHQNQFKTfvhLMXrmygl1RtccAr
n6uHTR6qMmJ4r3yHqhmJFajYRogEEA/e6YG/DgmW6c9f7vjxfwNW+DfH+0FPACUD
QO3+jDouRTBs1Zgq75jg4EYSMbUSj4zXbl9Eo/XmqcBH/+Gzg3mzaaNWHZazgRqq
6guCdWVy9cSQiBC6wOzVbVPQg+3J3jC68luPfMH3fiji0Y4sp/p19IChXE/vNTNL
A/Oa9t2Aa0Hs5/S53nsAQ04q6cvmNWYuWsbP0FbrzXhOHtjRUJ1tPYnwIMJX7dF4
WhHhjMqceR6K9ADW45yCjGklu9qH5sA1UEL5gAX39Un4nFNQR6NSNUVaR4qpMDwg
mgaZrPARTyTJ9boOF4dn2+k/BY30FFVCB5p0jabRPzZZK/GMRYSRh6dUt+oYilGC
91dyG7vztGPrvYGTRVL/YDgmtbHTOy2npCFVmjT+Ol6I56QEmR+2yNyOXlop289R
md9npX0a942zGKnx9xylu4ktTbXLGts3EqJyVTD+v28kllemoXGZAKa0O317AVP4
Q/YFPzDP6x7VIygdjlgx430xgAQgk3z4/OymZ4YC9fHJv9RQtWmtlZejjqwQ9xaj
HcqVQtmmRUvOFsXRS5qIgQg8qHnW2+wo51LoqQ5ItTx5Ed2hrs+1eyw/cUERg45M
+NU9m8HCVdwyJlyGHAtkT+s/lLIO/m24yMMnXrwSKcuaD9EOrvsI1yKBnanwYooX
roiLDs261+LketBMs66aaHgqPTNMmExGZbcLKeVx3nkVW7lWOuT4zJUfNZn/GCIM
TG+1efyyd5LZNTzFw+MEw2Zfm6Krvvc0jHtM1TDE/92rlMJWayixbunWO9d+mic0
6jheHAkLOeJ6t7Yx19pbSxTtR8QVEEQ+gEFJUy9Tfdq2hINFGKT+fRNVgrsZHqIh
j+q7E7EAnUS6WLlpjz8/Lf9shFhf8wFY2wqOgmQvvog7FfBvAs3OxDXbo9XY5y5B
KnrF4nWySyUPWy66U0sr3heQo73LNeBH2q9Y9ZykYdnSU5r2PPuFo1r9VUHHWYck
iDEuEsI3CihYZDvYGfPW8969tKcgic5/fJeLdO7Lnyd6lSYxMeYurq0koB05FVEN
bMcfuo9SNNi33m0QENWIMHBaf4q07waX9UhiYvsns2BvH/h0BV6ATWGV1y2FKuDn
+BYs5kGb4rEB0MS2NdMy0nnxOK3iImtjMGWUpAJKsUTHf4XqZWqUzltdGwsozkXc
Diliu0kyIXhq0Y9CT8DrYmhGUC/PYgB9Qy71fUT0oSiB6o08L2B3WWp5yqNxGm0n
7/VgWJyR5bJ/XnM30VR3fgwdqvHpGo+pK9fXS0ER96h9ol5VO+GuHji0Tij4zpGY
0l5cnuN9k8sT71jCU35M5eT6G7ZCAOH5UbMGZzZIP/eJl8sqpgUqBbj7u7iziZza
uuHueP27UXZEqrPeMrH6+pBQMrS1eenuEq9KisCp1qi1LRQHP6O+DphdUJtNdkkq
Y5pHVphWe338JVM20ybH6ZbLQPWPugVfXUueU0DKOCnQgjS9T8BXjjEnfTXtI2Fb
tDRchSHqEq6HhLZw+pzDGDXJWouqsP4k5OMxEWgOtjwnGeSZ7KEwMFufVLhjz1nY
h5sCIFQXSqysEs6bO0Y4VoBjy+QPifKTjHXe81jVyzhKY/QE29/boWpy6RI1rFTC
OnhVFKO7dDoyIIioDrEEjnGs7/T1ZVKXC5vMhW1vwISNWVDkgaW/O9KE6cAAhryl
WUsroawIz4lJD5nr4TOdWr9oVvrS5ayaD+NjBkG8kyia4jKhUgH7nF0vzNfVeIO9
ZFoF97u8JW0eg2JGF/DuwoSJKk/yWb6YrcvwE5/LGJfBhUraetOSfmsAQYwzH5nV
KZVQHggaF69RxN11143IdAobSp/koWjhP4O1MxNNY1DoPJGu4WDmfwneCRQeIDPs
PXMv25bfmb0md7PCAMh7LvAOyBTwvl395fsyfv3tgsEs6gZjjJUuKx3LUhP/1o2y
AB19tQq7gZ/H0tYmTnwDvXX8BzUQ1odbFBSdbSmFQfpSfnicFA7cyXY5h/VdvpDe
R4ZPu40ySvPhnqw93REh6GfbxGZkeg5w0ZTr5g5ZQK3fzsz2JUhdgzIyCpee34P4
0JyBRfAFTuPBu6UxlcnSZTepYsDxJ4M4l7IeU11mWTen04/vrIOWrv5u2Ef8nkd/
lBFh3eMbDOkX+nvREHKJgcgyM9WXdR6K+eF1eDmOrc9Hd2qWuJ9Sl7pdvzgSe448
tRNRgBIdkTmgRplBccnuhjdSAdFWSTGIbvaNZ4OcyC8VkQ5fnHrGrCXzldgVCEmv
djf7zFQs64bdM71Q8BxEZ/IcXgoueBU6SojRMofvvhZLGrwNmHWQLQU27wrzDG4F
/Kkt+1DK9Ci+o5v9quo9wTo9hfkrjThfWSU3MrbmFUyB4V7Ay2uAOJItCTXckr3W
f9BLDBDHDUw8xNG4ygqTbdELzAogqW/BTcrsvA0XkUGdiDVJ8Baikhw/gmpn9orm
uv9xbCMSi/bVyF7BX21zqF2EMdPZ5nW/sGjpg6LqIK7GAZ+RWr7NJowgv5cdIyKs
1KGb9nVmyKWuxdL2eXxteQAQ99stn1c0j4nSG54BBQGR/OiFWeNTK8DH9jdVTGCR
llftj1I19zOx5PXQMuQvghQXi19ehdLMSIPmmKmhojpa9uQlVf48Uv3idxg2Hi8l
k7rQ3HZ0xfckb/dF0By07BoJ1rK9oEZlO2FVTpt3TzXsz9fL2pw4TwjrmDIIdxiN
tMZ1Jwd3PNujLeoCDQ1JPuInNUDhuIimxdXzmNYFVnokFxIRZItjmCND1O8FIPBN
XEPe/yuMh6bs+jxPnDhdnUcgzZkMqJDpE0o4D+4h6EardwZ0AVFsC/H/wmG1xvbZ
N7R8oRMv6dpgYi4PySMMbUjyIWjNkjQtP2umNnsW1dzdjaqhKGj/sN9FD693M+lq
eeB9/7mSS5FI8o/RGxrKKQ28/iRyI6LeJDWrPBG/UZ0Nuqe6U5XOnEOOILYgh/DI
GTA5PcNfXtWMZB6XiBPFAG273TZp/IwIXRkyAsY7yegYM8nnX1V9Vw2pbEo6hI8E
Ab3YcLUHv2SSm9J+vOCtOOVE5QA/Tf+BY9uVSUKR5UCUggtpZTi+jMHxO2XdP4hp
pB+j5KfTgd24e7NNpnlaBdcbolEILu0qb6sHISZxnXmSyMfreZUD3DNtdxzH5nJC
8cNxUhJckG0UJ9WAY9GEDAFNrO8GcrwvfwpnR78nG3cDjUmXachX0+xNLRfzsa7E
xktDu5I463Zvs0PC6Om9y6zghG84RRQfziF7wHJHGq/2TeeBhz41rRjEsYKRcRnU
g3D11C0sLTBXkuGkjAaehA4BrFJyUVRsmA93e9P7FIPHixJLTw7bc72nYFtkVyu9
mftZCTMCLMF2h8kzMMWjIBQQmJEaedNr0dvCCmsMty1gx0q/i55/CzBWHj7/FFwq
rCeW9A4559/u7rOkMHQxhXxCGSI2cMFaj4Dw8pcd3BDaA+YRb811NYkxIWnUSBl1
koRmIJV7qJ3p4j+VIdZ/byUN4ioApFBjMgTZHa0nrmxKEDdMz/J8SC+es8FQ9F25
J09nxnHvNzfpKWOKNnJv55sZXGBxpEj/gS2icG6/+iHMs77OaryaoLp3onAG1TIx
gZ6NywboEa+JKmQhEUSFAs9oM+GewikoWZnjyWudpYuSuzpJV5w4Azm4ceOj1rRK
zV2pxBcXFlsKVmwmvjf6uzXI6UoTVP9DVQAB2QFjjFHhF/u+SzNQYQfYoq9Ibxss
GCqzaneHHzZ70EdL26K/0WI7v5cVeswC2c4f4rfIhdEP57nQbcTv2biUPLilsQlN
O7nSb1c4v9IpkvwGl4P3W+T4wCnR8LUPPtjAJGbFqKfuixbJBEiiN2BinBoDPg3S
+xbEIiq/9Umae5KwE6KZpEb18of3X0uBV7ZmA+a28d4rMw/HX+BPT/9AS9ewXuPK
tDTwKy+dYfMGLcXyCAWwI81CrKKR5vv0bgUhnFyxCP0pGyt9FocXTCryBVhF/v+M
YqzckUbT0YKBOI4IsuyzpocqrcC5oMmiyhkABEySPlPzqXUX0A3K0uZsnUAMbA5d
Dah6/JcNXLvnt86WVG/NsDYoErJVuH9gRXPeX/KrFjHzHxgHA8XpzhIOy81Dt63y
GJYRJoMLEEGC1HL6XjutnsbYdjXMh1+ufS5mcZlV7VNz6I7NILyFYBKDX1JaE+57
nuvDCelYdHD9iF/EOxZZsqwYKzh7wWV1OXIZEwk12GldmiQ8rwPoLR2Q6AAEvWLo
RQIVXYUCJHI094AUagy2i/Ua7rG3HhMeInYgOGqqZ8+Cw2NEzkTgl0DctaoKDJ9s
MKEeis757baS4rrCuM7eM+MUoRHRg7EIPUWOm4nEha7kxylpHMYryd4TMViwhA+o
1Ic22DWaaHDNkc3PDwvo+2xYGjfoOWqqZzNnZ+OjVtQ4ODblac5kdsr1zzQyypSX
rXZNocDmHA/IwZNqhyFBX2bSXHmdEknPZ5Z+Ne/z6+2M4b8X/+swveWVbUZjghKj
KZ5YlDnKtD+N3Rxi0+ZkPP1JYBS7pqKXPEdYAUp1aaXbUJL2//jP7OINdRZsnPce
onLxRnS5Byn0S3Mp3FrThI1bqXmlhyuckFWu5iHaVruoujUZSN012RsUOSgDYsGY
56E9nD9BWv6l49duD5Ws9gsn8v4vTOxNU7HOVgXEP7mvLu5kHjclidX93ofND6zX
u/974ZESPHEJbNxuG29KNJPr3JakT0Y1UFuzFUSaJ12OnWR3uBIfUSQ0paUK4dhf
XSiQNSq+6HfEUXQC+JgTFCKf66/dOLFAMvYUlai6VIfSEYDQ8tmGhQxPyudxytYM
OPlqs3I57Qo7zH02XgzJ8EGPVAdLpsPVOFONd7b4swjmqRvb1rqBpxEyjGjxMUth
ApPztBNmoOW9dXB3esId29dFeaEP/YNGeNR2BqpUHNd9g6JvRG2McBhgQoP6jZDZ
sX3SjyloSHLgwLw/SYmdKJmQh3Ajb372GQSPzEgo6nvQhgZjZFsE9kN4B5grIROG
B5A0qIJ/zgwJ30EtdSs2GmCIO7zenqt7IXwvgtWJ81yflhQPuqbgjTbnviPT/bC3
SZqdoPl6MylPe2kdSWM013L9CtxG27+tCL9BbtR7+dDnaEVoMeJjyaCEnCLGQNGo
wgX3MRTwOnXP+Gs1ysjDPCR3JZFFW1ljNnDxXte9MezkJgdxO2rvcDFexnlXS7OF
ajfroHd5Sjk64pZzReUEi9X2NGve8eqbmfwr3gNohdhHXYY8mvvNjsPRBTelBDw1
wq42HAuW3j68g4RKhb0b9raKog7/0EvvdgkXRyT6Vqf4yB5NKT56PbWSQSoh3nuj
Xy0QFPjtDrBGUXeboGPlQasVRDE5nm8pqac6tlMXsTdY7RBRlNvT4PAE6UExIoIh
26/+neTEWXTSDQET8QCgwZNcdrI5kSSnpFLRiRHHjVUmu+f2XgsUDn5cpSEF5x4g
hWBX0Ocex+cef3if7sjvV4xG7hnFP1Le4aqEVc5w368vg0qIKv54MQf4+J3zxk0C
U9pvSb2X9zdNQhlOJmWJxTXMHZc4qLgFGeEVMBWeveHv4e0t6iD4GVOwdz0Jxa1Z
BVGJgVx246+fKgVjv3e1mVwQ4kvA7K1Oym3pvFTbYt00Xjbu47Hqu2ZJksAwBxz7
et6z8LjGxO7KIm5h9c6aICm8ugOWq6UmIuZNKdKU7Yo2TyewHbqG3sYhB+o8yk+i
Rfd6B2+hnDoAnnMx5vLnGCp5XCWthof49R0MHkHltKXDk75IQFPlZR96ipGKlg6E
ALAH1sbX+rOt0W1G3hqbEQs+AyRpT41XI4/Ai6EscDy9PowXuvYhxFNIxeS9Q7Rg
VCqipkVuIbluAJJBiFRe/2mb2PiGN2Y9ixK8+XnLovtHdMyzFUloVNgUnmDfSGzM
pL3rwUTzsuQqqHgdTwaWR4qiF/8Vg7KvfyJ5vmdEuz8exphKM0W8niRgWGkc/cdS
LwU/pCuuf2jizNQ0CbtkqnIo7zlcXBA/uzH9gOoc21cYEbZdIXxkSNWkPKoYYg6P
CZPIYD48ipxqqRWi+K0ArHFJmYaEKe2hFy+BrItneqk5HsFVilsMkIHujOcMPM3n
6mTqGnAXS1wHGDArXouyioQYzSRgEEtvOZZ1KeRYtmrcEyQbDXWQxc2twoyGniLN
oT63lL/K9SSdNYCFnYJLPwGbpQmvV9OgROaaOOAitsp73uxP5uVMiKCr1yx9P9if
vsE48ivRD/0NpspvMaFi384tA+fwGMJjCEFBk84jFIlwdpFDlrbQXb15I7h4/o/K
Ledi3Y4arcj6EAbc+fxwmQTgAUF6DuHH52kfusStaTeZB7+AqIz/wLfWarNmlo2N
YflKzYmdnA+F8W8rPR7X+m1u1s+BSDKM9meyRtj0ihpCIVxAvBEnDGs3haMJRtKS
/9hE+Pgs3u49VQZEUeKtsWgxy9AJJFALBldbKxdlgiRijAybd4oFBe4EFnyEbCjU
bLTfEgOZpdfjhNEEHbMe5dujQ0Gx4ro9i3HDpPG7S6izttlm9ZCXlPXso0J5SkzQ
1SeEa1/EpzO5nAI5prdcX7rcGthqvbpziptRZPJjqiWaQ4LlrE0/J+hkpFzYXhn4
ktlSB/sU7ka3OmgaluRwuzEllKC790QvQdj4gSZ5Fml5y2WS3d1VjxDzZi7bIxn/
N5IJRObGxQe57uXWtnFqkorXQUPJkRLz7kk5rzxrDKOcLvyOg2gP4KSUqLXSxmmy
CXlY2e3rK+qWWS2xsfO13bg8R8gi2b1zGwWZR8qyqQSmpJ+3p+ns7pF/AxtZDKdA
3cuV5ZgJcT9f60GSveXvtOllwABtsb50EVpVIdn+fNwG+7/CkwNOgVA/VYKORNAe
okRuqgqoWVGaCWMEcNEsDbFk6yie+FZM2IPwyuCPt352igvFiLxZ3U+62HiaDH1M
290mI/G4L0k+XRvxoYtEujbw0G93OiLkF/6F7oX2yf9ySJgHEF9zW6ZB9w6R660u
nEWcRw+nvPtMO8afSb7pHCLaxLsVXyA7ZHwbxUI5Tkc91s2yOQ/4EUa0fQK2pQvG
l5wbtdQCQf2WHcJdv1EcUW7/YgAtFsvkCJSuj2pYJ6/TXYAXVigrny7gK48/uVLZ
AFlTmdyKEkkx7U9fzQ1cHBDlOwkPgPF4PEf890daVTQXm1yCIyGm0IMY9/TUL/Sb
PDYNa/ivWtW7TLajM3to8HOgRRJP2eYxtyfoZfr0cQObbyFakOVANTw/fyjCrwTK
ZpjmzAZ6B6mOXqCTmlH+r2HvIe9YBciAMCD4COcGWHkvhXw8o9643LGV9lTlZr1O
fo9sPsuG8YnnVmp5Id4tXmbMf6Wb2rKBmGrNSOBUP7A6kzLd7a4pnjg++H8zeUV/
1R0F0tc4nWXiBTYPxSPmH6Yffu9FivOY8dmtfbtzhwVowkeGful+C4hB+gVMM1lC
h3YzYKtuCSBwZr3Bzk8kOGwTKBY+OvbvL3P3M5oGABjGJrmuB+NyNnrg+cSbkavd
uRGsiUUJRi7JlU/M7R7kiX26uftwjtXJ2vWCIQRk1TUH2HmHXHyWhnZESKCiw++N
qb3f+IvFZqEI1y4tnK6aW/oqLiXZvY56C5MozfpfgEqMkRs1Sk37Jw2Epk6QS89f
j+cwGptUdrEShS/F7cc2RJXrS9pLgyML+Hgq7UuzG8xrgjGhfiJQTmd4b2DK7J8O
hBDA8ZuFP7/IMm0iluN5otVjqT6bKzTQHRtTVuJFRgka/31iXmuyamZA/jY3iVKj
YD3tQsfWtFMcvsXmjGtV+c3VU8QTDyfCYuPEGT49BFuXyfLDF/TMDxTO85mrLUSD
QNnMADGcuincMubHfIrZQbt/cbRJfsgDu2IZcNQ6Ogawwzb1xdEppayTyGy7RQR0
1ZtvIKTGmHLH+8Wejx91uqmS/WZSVJaX0grNWQ1HF3QCFX2zlPuyqYFZ/cteUae+
DLvIisAAyWli6VEO2n48TOl6G0/Lr4oe2hlFoDBr2my4pFrF3yOc7sqJSxtJe3IW
lWRGS4OrmGBSkfh5LW5LXl6p1pRv6MMcyPFSxsSQVtNWlLlIEa31o4q1zeLTGXPo
x4s6ykXTwg7IZXfEZ5B32S05riqmTgbTHA7+MyfjPFuydAsL/0HpyCvUrGlbx05p
udWD/lmZNetUcaiSc1pAgN1XxBmk43huYwApueySa4UcgqrxOwhs71OkS4FWzCzo
97eqazDQiCLBbcPx1rVcDRrtfBKKgn8gNzJUNV9KeSQp+CghzXxlsgMpPWhgLYAy
QaF6wcvTi+pXsgHi5KoD4nkIjQXx12fzAKp77ElxJ1U7Pn6kJZPBXtkJJy/KBnTO
HsnWOq1EFbNwna8wOP52cz7IsKVE96RC1GR/on7K1nvygjNt833IQBYYz8tLgI42
OWEJBdTRZublSMqXpdc7SEBBDiK6pioqliXP7FLnxx9qOv0YisRn6gR7gYUulm7/
fXombGP0xG5OAN8S1h4s61Va43iSyEedbepPxymFkaHPxP8bxw6xBKDiP8fYUvPP
Jb/JwBcBRXK7YqgiRVog+5Se5K9Hmiz7uHevO3cuZUpE/5mK2U5grzdyRBKgZAxt
BtnWDFeoENz2U9AfyG7MZ/RhnVhyXnQUFzv76dQWJer6mvNuKfyuIMrsHOMKKaQH
bh8p5Nll6WkaFHqugGMsTm/blJoLXOpMaz92Sp8fZkrrZl2RRxGRdwVhViMLcrrX
Zv5fOPeMJ0HLu9BXeLjczaxzzVTaIs1Z3UfWnFovjkyrXx/9Fr6YxK573KLKl8S2
wmhGx6R7gJKmCrPjxYlW21HtBx/f35Ianlzps8DP5n0Iss3bCIIZ0iOrjQthztNB
UwiGi03bfIXpBc8IFzv2cKK3G+6hFNvyl7aD7QyNTsYXlbocdnl8pFw5Cbsamcpv
BJDrQH97d4mUDgz72m/GkA8pXh7duxtOdI3O6zq6j2JTXJRGcz1e1q6LDNtaE4hn
RbCIWBF3fdznL5itE3GuYTTzUkhSl3BQrCj4A8s0pBw6kiXAFm670JK13lWFr3ge
MLK1AQhyZW6qmh8uvhsbUpvrjE5tmjTOHEVYCylJb2C/hrsGKay2DON+Kby7OFMa
HBKfuU2PP7XH9SfGrxOXDiH0xXrbzYxY0hwn9RQEeHQ8F1F+aToIsxZVFyX9i4cd
VkRR5VNPPHRcIDk6855q+hQZZXU4KgIiHYjFr9CueM/1re3mDhs1CsmON9TklUcB
aL7SOuS9iEt7fBbgt8UgZ+F3GfVrGXniLlgAA/k11HQuj02Vhimk4xZtXrgBPo3W
TYdTGQkK9JgWOKH3tE4g/wrlrrmEcQJ+wPXGlfdM1HbJspzpirghrv3bvRruiPEp
2UacyVwKjoUHwW03NHMtA4EizVuStzVB9GcZnp5Qpzz7GSwTbf8J4bAoHMkMLlZd
CMcQoZ8LgJmxu2ncJUo9rcSJxVW1qGJrxK3Yi2VODmzP1tHgvdZF46cUTu4UPTSA
nHEbiO45sh3ZcboKoilBgQ5ajbadvcCUB2jQhsTHJ2NzaLSN4/3p7JcpH8lwyh+e
3Z2CowiLxIszmqtTrZ5sJxTr61KTlhCCemVDafnSKOh7y/KbF5shBqu0jKl+/KBu
Uon0RKqfj+prlzHYSi0Grc5FGoo7alvYNi/pzujQl/CFl8Htwbv1TG229RWgQW7/
wKSCJPvbrNAuHOCeyynqrrojkQlfi1sR2hhOjGePYVfMGfV6SS1L5oh0Z3nskJBl
qssJ/XlTuKQAyI7ftACVHMOaKVVeurdrd7LhGDLPUo0IymW6HKaI9b+y98mEr4us
p5tj/WeOzcmQbD1j/hmcCgfYNgHZlC/FOxGSG7FyExJKMnX5axnoBtUXmRV42J2k
Vwt9YurT85AkYV4wl0eeKC17F7bMW6MAYEihTTPwZPL8RdZD2R3rSXymPHiZZiHw
+l6lGJ19RU5/rzwOblllQ8NRSGLL/OJy8hBOJnPP9uI4hYsaSL/Ch0yn0Mxh4gJK
b8GBuRMMDtHAJwDgu5IUtd/k+xcUoBGboFKjIcnCu0k8TzA6jtwePPpfdBhF/JSq
SJvK7YMyBXFo0HedkdYWDqyZJZkAYm/yOA8OSDwNGqQgF/SsE6pf1ubmLSe0O3sR
N3sd2jFFsEyCKWJ0lUsKc9NqfLLEoBpikHk0+ZbsdoHATER9xvef55ysF2vxT0uv
n1W4IbN8kMOfaoyjBpLakVcqJ47742Xp+WCl2hco4tAW8+XJY3c2YqALg19ttCLE
PzsCOtxzVnMgDcXzbkqLquViImaBK/YQo+7NRMB5SAHkgBPoAcr60L8LKpgrPkc3
qT3yvOVAAhOoT2lAba782sK0mzsa8N/aqmR35nl4TW/uBTNbz5IUTPkT7t5d28Eb
uCEeRf5cd7vyPKAmyl3uh4NocTJFqjB+W14bvlvARC8hDBsiJMljhybyknBexyVb
UsPw3WQM/FJ+FcFFlkTplsBidXrtbkmVLL464P7Tl5zZgtEJhnE5T4+AOoBvyt2G
cc3u59VQKyUqaZyQNieLgsO6GWjbXYtkBYgOtuWaBORfZregzfwszl8Ooji6l04y
Bge0JIwk3ZduDzjzMwa8ANqNNkIGqVh9CG9aNNz6iqDa2DtxmX4/SAni388mii6K
8GNDx8IKL7uBh0tLQfAYZrV0yVEvYcVWUta6KxrIimkDsYyX1OYdR2aSyNLGGeEn
rTwba+lD86BK4DZIH4jkWMHc3XeYk4sSDQAcX7RB8NHQfqzzkaWaHsHoW8TMmFZl
KICuvHFGpVtXJPUlA7hfJtshVzJQ6bXwr6550gmXbbrXbfIbtfbgn/NOZDEI0D/8
rUi4hLgci6IIJMCQpdGl03icy0PZU3byQT+SANONRxWml8N6Xq2v5NzScWO3DUA2
rKgPQu7AbTx12Kl3t4p5OHixBVUoT+yjlVD85uRt/eO0u0Z5yBkWYjUQx9IKZBeZ
wEup0zFDc7aWwXRLQ3HPs55VQn6uyggVHUndqTBwj6o5d4Z7Uie1n7UeXsbGGd6u
jMRzuCx/Vq8MDolFRy5mbacvJcLB8Caj2/TNZVl1AKgutYbOoz8fscWUjUx+TBSu
QjrL6yn/baQIe7l1ZSD6+kiiIGY/a97cIh7vwf0XfZ6lmYaEbaeRoq1qUyxRFgbN
l13XPlk8+oKMks8tXar/g4kj4zuv71U5a6ylr5nR2fIs4rZU5hfSXTudqm5wPIFe
XA5wQ1cfqpMpKzQXO8iWQ+heLdsd8mVMfQgNzdp5QVnDGJF+kKlWpghSWLf/1BVg
NUsOcFSAqWKG7K3Pf5xq6j86mYqsxhXp6HuxfYN68OOVieSGYrnVzgUkpm78EWZe
Q13LcIA/B3ZDSFtzs5ypWoZ0JzeIlo0HtcVbknLM6I20hG2K0+odrZ+njJtkh1F5
CjHUiksSqqLpOYf3pugoZSH1UM288ryFecVvjEuPSJ8BgzQyQahEpWc188Fi5zC2
ApVJvDapUKF6/oHEdDFNTepRJHol5maW4SqQeVuKOUR19resBY94CocsyGDgEDjG
7J5ERMDfwcF2WV363CUAp1HHkFcQ3ON8oKLC6kG62y4k0YFQ0PUhCMbzWf54Oiyp
0uGBBn6HnOISmJwjk3Y1KAPx6p7Qn/B5foDZivCYoAu90xib0ABQ/AjrldkG+K3M
mkQIdyMucAZT7Ko2Vb3kPTHGEfSkyQbX7WYugBNWY7g273SnYvIYOFZ7mqKJ8ihr
2BOoPjJfA/NMFcxKhGSWy7ZhwId2aKOGO1D9OznFa2TfDNZ4S5eMepO4t1ceCRo3
CuFmyrF4USOkPjuSNedi2JLkUzXnJo8PCF5HgmTPajuk1APSD0P7lS5A4HGKtPbB
BcQmGBE65S/g5DIh34KF0AgSmYvaV+sQP2xvioevKpePnUBtyWx7IO9ZV1iqME6h
yd2I56Fq8RA3g/c6D9Mrfo1gMruTnA5nLIXknSrigjYQyy0KNZZorCB90EYjnYwi
Emw3acFuj2hYRWV2Uq1OKk4YH+EH+l/UogE2I3nju1xLCn5AYD943QGmEHyKl57N
JrSObKlCop6XjQFhfjGczX643+yI8neqq2GaSkBQoR1Dzv29Bh7bf6iUlPGRk3kE
2fEJj5WSvTrDcE+dGnyfG3mCnhW8FyjW5/ejLSBz+DVhLH6lk8sUNn2QUHXEFCEI
Natv/KNFMkd2EdMOiVlarZjsp14G0H4oNXheJuu4BX4MHRWBBmmPAuAWRwP+iBGU
Gpj/ItAC+H2PEwnTcIaRKJvvUuhPggj8bBEt6puplSXbcnXzC5u+tHQPAZt8Azn5
hlAm0UgnC5cHwP42vJ0lBYCHluenADJNe07Djr318hoxkG7r/fjLcmXh3/nwPwts
pePP6c/ndSCBoqTy3hce2dj8Q2hCaE/QR+Ps/vubSyS1qUO9ZdqLsOys4VOsrbUW
hC13wnh8BcC35esTptqPcPG3qCcfkcnkvyLeXGC0DKm9VEu1R2gPoUS8U1QTV1SJ
HKOGMRwI7qbsxK6B+zhK+DdRygvvduMJbI2Cw8reZ5SHcw0qytmZU2N37e4DukQQ
p8+TGMVXT3G0OEmZHx7pjBYSthXXBqsRfIYBzyJLky5N19at53PlzDbMTkCApBKS
5PLK4JfhGGLe48HwjGOj5g+YBwHy5C/ebPQkK+yP4/YJnIh67o+PLBmRTwMNqKrE
Avv9as3jEPuFZUscIS8Oqx2lILFt3P99EogL9zr1fODTaE6oio+ed+rtmf67hAB9
YlA5DZm/3/YE/U8U7LN9LBRdQK/GhpjYFHpi+MAf437duxVMxOcxrIcNDHFu2u2E
vcUKK+r+C2+3aGX7KWuoZW6fBpyNGOkuEjeltWZFN/NcnFBPMIGUZuyiNNxowdQ0
sfkgCOjK7O4hE4IEUMS51f2i44/zqMwi3JmwrTzCbB6kTj6oEE6zZ5U1pSPN+v9Y
G7xINUwFtaRaSrKIr7jf75o8uqazj7NzhQKxBmY2Osq9HzxohSQCHOLe6xEpur6P
XkU6R8fEKekZmoMftLGvswWSn0P9wIkXvcNT0+38Z6/Vf3FsaYoglwSKt2u4X2pG
+zSAVXgH8ufsZOX0jxXTLkVStBCRPIwxX3RGzlCX1LzlJIM37+o4D1EwHhwC+t0H
GO8H9xHk1NFtRgxqE5BkendnDAPc+2LfGQIOdiik6ar316ThHK8KKYrwy0rERC0s
wYg9fNgvvw7ifu5H+wDMqa4a9tiG2DEnNvbytJtWPCXp88xQ/J7WwNhKpVqmZyr9
fokMLSYbYeJjywEVrj46IXuXd4jPLC7tdKU4g4jr3jg3XdqIstgiAaO7W2rv3LBt
tFF2kSyFEMZYd5LKeaQe9a5G3fhC8bJto47XmxQsjpqlFGnHKVdLjGLSv333MXaU
IMOAfGHxMBWGeVbESGJyI4S5cxZaZ2mJeQG+W1vXwLZZbiEqtyVHgkPQo6UZxucK
TpnZg2iMgqW4qYaBfJ8ofMwVj9hkNS4POD4dbzIFM5c+BrT+d/HT/EY5ux+IvDRZ
qK+vUfWM3haW9DNWV+leAj+T7034wwyGYXjlW0XRS7wrvT3ETn/wdzyy9A8BFXdu
L238mFGW3KOv1BE9mI7GhSUiJeA4cgxSX1RTXrAd1LyfquP7z8pcpNBWth7DxCJH
dPzX6qv8ed7nfr50e7cbl0Tgx8TXbCoV+nvJx4ilizZ3Rs9iO10wUkU/sKNsPqhC
E37+9mKPe6UXTR0fkTCc3cth652lz628MXoS7lSGk2BvhpGUxC/yw5QEQhDhzt2H
lmXX31+ofm8xWebkAT9CDF3IQ6ESydc7spXtM9fwMpuh8Xda3+Jv7ccEjB6xN0wj
X0Kqb24ZY1gbpcHJEgUSfkqqafeYtEgFCtAEQZYVZ2g9lMTru/we59jn3O3RTuh3
2guMU0/7JxYrhTYR2o4jPDHoc5Ywzknoe2LyLty31vbPcVQ7s5cjI6sL2JflDZSO
O5i3lck5/Xe7fUAka99D9ncvDHflv3Uhnqbq+BKDLkFBsbL2Ca83Seqs0qssbf0A
SJQSS6BiHXckOG3vhlPr7JaH87auAuyiRB6eO8dRFATbVO+PNwyQgY3oPBrP1wEo
uiaBgzn1GdoP9+U0pzYg2sV8HRQ8mkqEzGPsabx5JnElmvns1BF2KPVMcP6MUW+2
WrtPMdLmMpCpG/DY/aBto9DnNMbh5wadUzL4Chbw3ysbXOTkRcDj/X3kj90HF7vy
mqwo8QCdsBXC/w+nufT00m2tPN8/8M2ynaBObnN+2Cm3nMANr/yhC6O+9oVgkbNd
RuNigmt5bdyZNVYhPlSuTFv4gAHgZgE/GbWHBaWH5Of/04yiW9EK79QeXqfnx/ef
Ygf8DzmT1i8o0Zu9ljbwZW4XHuHH27vqmr3RpNG2270YvjmVMP2g8qUSYskZWJmo
RW2cJ2VbpL09lzN7ZtipyfBxD2Nkh81Ay8UiqjDk5jW4w/IAY1/nr925w7NR/YD1
xNpHco9i5tGRqRMtIZQu40suuSfTwVXRzYOMplu2siP97jqg7XQaT7eBlI8kMj7D
HtaoFRWQtUFEvjLU+57/kxpJk2yy4RAipvbPKpEDDdpPGchY0FgMiUXGyG7aganm
OmTx90VbVkkqL3XokRyRjhOZFunYnsQPGe7AK+FZ0PImfVO3Yt6GPzPos1RHPNBi
HfHHNYzPrbFiWXdejHYPRvjkF8uG5NW0E4HTsjbbtCs4JeGhcXy8J00X6UKJisHk
KsRjFHmzfS+jM2YApTg58/5NN7KRdvRDSOEt8MstNwfOO8VV+E6wTn+X3G8hd4Jl
8afjz87llQUeO0VI3N6wgrFijRrItlsr6g3MH1DSDDHMEq0BLk5tkiHasQhwdPX5
exdupIhb67i71YpCgiXaVX5YniXmJKJfIez3shGqame8mwMzL5mK04lMVOLaC0kI
6dlj5iWd42OUjUehOwS459oZqEKAnOsC5DgmHcBbCiNlKbamY1dQ40NAjHKSJUIC
6tkGI+zSgV2deFzgWVZA1KqQkXeufgz62DkWPvMl3CP4s2pyvcO8iNqpMZJWMwuD
l8mwC0aB2XYoDlyPLTTiX90WvHhJBBf8la0Rv9AdcGZKTbfdxkVBnWTsQA52Q43L
+Tilc0pEj9/Jw8MxlVN5Taf7GuEYF9Xsz9koHXJWV1qCQVp3/HZt9zF76sZdoBzc
maz+VJHB1YGvL7Z3lHBudFYTEAYu/jnorOfp0b8n60ZbK2GNwJJIvwhaGvfEk3Kd
Ednsd81ZrKSe7DrJr3VfE08hex4T2Cu18L14Fr+qqc3+5mpVtL4c67Pl2JvY0gIK
MjK5j1K/xX/9WYA6ID0ub1i8irndI4OqBtU47nMqnWnuakFzVuUrzhGpqcTBv+yo
n14W/WlTeaRm2UhWLO/89PSqEfZl7x1yEr/y+SFqHXWjRrZdQ6Xuu2s55TAryl3k
eAhwK9bfh9hOMgkE6OrcIPEaBI1SE5zN+etVLsERCE1yR0flO26zUKxorBAqCGPu
JW0BvPCIMCSH0PpjBRfgprclXfdCnxdxTGqgLpxshJj02zPjmg+NwB7JRt+w8t9w
/NdXXM1n03aOEjHMORMBQZYQmSvGJmUvIRehZRw04ZycIUOwN0WLSVShtp8vmT8v
6QVCDBqCAUZVTE8a9E2oDdOIDzE4tb38t1J7aqY58zP4RQULj3YTAJpKLChvyD1y
6uhMrSSz3hc6tgnroq4XgLUX3HwKkmXOTfjm1kJdEoJbEIorD4iUzw7LwPal1sj9
q74etW0YamkOlmMt6Jh8yp/ZdoV63eLIXokzbhCTxkL5TmMY5Q0NnWPskS7yhFXE
w5t1D1UaVuKYbNNxd8/OIq44XEp8EtvrgH+/AgPi+/gXM7wyi6XhlmdozZiRaRAi
zErMZWZ41S16g9PeW98FLPDQPRt6TP4VhjT/0GguZ8JZ7vfx71x/24Q2p0796ogA
0CLe/a8oqmhaVZ0z1n7lVfHrCHi1kC13TCSCmt4nYgeyYh4KIXwmlqSdMsnjYXMt
PweiKtLxrrjoqh2NMadVrvNjQVDwlfADAUjWZUgbATVQtIQGRR88YM8MCeVe4zG8
YshoIZJMiZ3mJtGiLmr68sVpkjUQbu4HjNbdHlf27/r1lkdvXtRpJJ/K8Ok+rSwO
sERoHUffqIZp5kU88MT36GiBo4uhB1BeX7b+Sq3kX6RJ25bo1ENVDQn0O1Qmca1Q
9t/eurutMkb4pq2jqxxtepWQHjZFd+OV02JpFFkx5LcxPFJhrhTxUGuOovVY45r9
u3mjqhOWpH/FYqw5vyjEEoIaLNEj6mTHTOBDewVpG56n9lXl82chn2BsxP3almtN
YhrsP4m2ElO+MSlz+eMXsIQyu+Gko8MN5zrgwaaA6YuqoawSExIqQ1ykI63eaJac
ZAP3XpnpS+RtZUxYD6n+dIYtDMCs2rlxd+2J0MKSmRk0EwKEkIUMtYZIFHIccFqK
u4/cUNom5tfXT2Ksitf0XjUr63maqui05CT9J4ctVXwyTBBn96pLxoXaULTeVz3w
M1xVQVKQ6ViICfrEAdLMGR+JUdd7H/53f04Ljd/VBoIYj4mOkKh9NNWuSSXsMo43
aw+iVnzKsT7ch4e6Ch+LJhQ6WT0++kJYNa7BivqFCFerR1TsXJ6obcHro3IM9AKj
JJd4VqgNoH/t3trhHwgrEF0xAAWY0OLfGP643CTychCyoiaLDZma/COr+bon8Z8/
dbmbQDrzr3Zj2jG+Q1rAQLwbmbD1btWGZB9wrHK1hqJm/nHnWe4BX/Gs6d0yaVVL
iOSO4urV44N46VFewuYPp+yG5XoMNFQWZTEdMeTzfOj2559HyeRlCM/Jd+176MMc
om7kuL/9fp0gkFD4lzG+ClSAXPdnTglcvk3uKzVELJDeNyqu2UuqmH7eNOYUy0h7
wyjKS91Pwxlh1f6AUyhEoWBYPaa0fMTJl7d2gqiaqvnAzpNz7aKhYPSKBZXUUbC7
AWadNA9Uk6UO+KHjf7af7l1lLHmAWzb0s49VZNoMTgxKwc/uYd4EGFi4WHjG9K+a
Jhj1/nvtgjM0SaoBJIcH0vChGubblLM+HqbnmyVWCliJMVbC2eHix3ATKGCfpDuJ
FJ3QQTalK8Cu86DbXFoeQsLTQQ2EtC7eSNduPpDro69z8Wda6b7eFEEc1eAAxUIO
Lksg8uJmuXeFJdUeIr6T7oTyNg3nOySbAiXpfkyJ9KEOJvraWf75ODiqPK1rn5LK
4nxN95GuCjwert+dMr5zQDLeUQscYuwpmmOHvMBPKV4SkwQ5x08FnDv2/rKzKRTD
7HP2nN0R5UCD9pqe2W0WnESCeN4KM5vDq9soGTg2NXwcZlPkpomx518wdfrTuSyM
MhmmP5uXCohO9MLsICiadZthpV2Ung4okqBHnMgepkA/2o3ZJ1yku6VXAvO/XBm6
CP+8ch9HPUkTVIUUFFHqqW6KXXbvJAgvMgx8rrupSr1YSU6Rupu8ir8hQaC7STTZ
GUDmWjhFNGGdDbT9sfDiIQQ5fNUbDKcF55mK+Y0swtCsuJfDlj4FUBkzMi0yYO7m
3lmC4Wqbf/GqeKnDkj9Pr/0oFddkKIHVvprvfDJLj+lsjlv5ArbcPqxx3Qx94xIO
9U5upqq2qpiqDtgWONmmazWaZLoETSWFSyiiX4uTrK3kxI7nX7McmRDOUJkAHrcw
nOBiivp/F/wlx8YNqJCuJuD9QEa6ykwRhZruILB2Li7G1YNrEaqRZD1SfDVwkZTD
CbM3CGoVWgnkulxx5OS/vNFHLvU/Ibi9ZnISmOKWJWJDwMS8a/oExsv95lUFyMsE
5OQkDH0SKPmQd5pg2E4q5T4kKd8ZdqqD0UDWi3BktDgayaIf3yQOaWNLlTQN/z0h
6DfZiVoReIIVY3gzzVSbj17SIJTZ+/njErjhbv7ncHZ38gNaHtfiPm/z0DT/SEXQ
zYm/wP83eMgcclod5rQ1VcdNNJwYIDr+T79o1+Vqw9ETlJW9aU9xMqPkMHlubUTs
84SS/14E41NdONQKhTJdrp0UiZUYfA9dM8lqmRHslzl0X9FoZboWmtIHtMvVoPZN
R13PBIsDlr7Swj81sd3fILpaz+dB8r/JgmPDijOVPx3Rx8uKm/ve9TSnDi+ezsJP
+jAOBBvW1WNUtHzzXQxDMm1HM9VCbgFYc1ENM50oq0+9TWjLRTvaM7SBB6Sehjv5
BONIO41/C1DphqmeipuF0smJjWgsyZsRcLN7jp+YeLTUcpnJ7/lX18jW4mUoBdfW
WqiU3qfF7u4jQMEB9lFvk8nfaZqACuxHyJu1XE5HgBMTtpGXjKU9slGftiiGaqaR
wqf+jYr3o63NvniII2IH41zkYPhszCIC3CnWg8v4nqOpZxIeazIpaWyZHQ5h9NLq
ugEEdRY47hMBPP3f6T1xErdEsxWN9GTtIx8VxD0W+UlSJ/Cy2tynplUVPKm4fmJP
F9rX5iBrI6eGQW+066CCntYPOPCev2TVXGOFH08pv7J5ZsZrWp/8JiseFdOS+PzN
jxADpH47gtALdAKib0yy7oKMVL/LAeHvEvlwxkTEEi7mvSLdylcyZFc+CvrB9JKX
vxuZXNU6Jl6oJW/36k61KaMsYdJUqARZTSPsT53zk+1mmQ9nGf1U0jAS10htDLp4
hJqu2Vl2CxKL2S4XUA8r7fqHiq6W4x2LDxNgtpV5XeA1Io44kxJPgQjxHjLrMORx
RVtFVx3xirZ6FGOLTa5wpZrz+fDmcQBLhtGh24si/kzHXEpMtl0rJaAzxOuKhb22
DtC0dGrARzmIe527yhsvCbSi82QUGxjlbME0bgbTPBNEZqsKqUnD6eYdaNmOpS3k
v/cNDb+nq+Z9ywyTtMllfctW+nQnukowtOLprge4GTiAJDsiix20kaha7TKvUNDQ
Ntr2cAw32oyK4+tIUi9ojHtWqVrMJm02hcewwUB71PCEqVczG1r8XDPUKc2ETkUW
X9O9lvidNI9+Z90TnCfecEbwk4sk5psYvvboGMGSgnwss447AC2JvfMX3QH12uBM
eNn8Dqj7l9TaV5IsdpiJI9GC/Ll/duVQexDA74sz2mHRxSQz6Z9DYLTOtohGKtfR
scUeyi7sCzUvjHu5q9G1VY0nK84kVUkyOOat3xDjUlbQSTVbsf1gFTp6jNqLlU88
hdbUajFWRRW19PAzrxWVxZUBBqlVEWKZBqMw6hTS2YtAWYqk7K8vd1Rvxn/qvP6E
t7RZRYdrUoyx5mBoYlalVwg6qUCnEDcnFxBOh4t7iHomo2k2Nnk4VXmSYLGCZbzU
QwsLvU2bJLPAvVz0lEDkpacVR367MeHWGgfiHoGBPBAT3Gk0O9eXV2F4KXow2f59
sdqRFZyXp+xUKAREb56ig+eoD0HfWcU4WYrLmGId772Jz2EIfkd7jq0Q+zXgbxrp
P5FWpn8bYHNo86XAeRmi35uwpCHZfWRIBRXnWD3+TfZrSQcxQkrIBlXT8bNE3qQB
GITo3JVqrYovWg0779rXbST4j8+yHGLybyOi6c+mPoDS89ucdfI4NAry/DJGjL7b
6DB8lijQj8OeMlHEiKHV5ZnmSDY+QoJkTJbP8/utUL1TEs+UzDricOFbmmJ48gb4
nvTm+xKXAP6FwUia5nqwxFTxysVV8+JvUOKYslcH0s6zJRFPMbnzxOnWRn3KuVj8
5GqezVUeDntal2VC7XdT0QG+49TCd8vFFZ0clWw/EyCvU+DXDiaib4S6e/LJjs8k
DcDJGv+cneuNGB+X04EfVRPXkkwf/5rZxEnq6bhl/RlnQKBYpQxNrEc5Kce3ksZs
4uSvpJfFVO4vj1mQPGJ89w6uZClSlZko2+C704mnO1AZRWOxQ5AmaLHBJGlFkHH5
wHqqFxb99Fq0G7qiL1vl3xDyhEhDjv5SfARSfX4KQpworez0UCBWAzPCvEJBZZ0+
mIlrSwzkac7bUUSIJlRWP8fMYQgqbQgGQaelfq8Zy8TOieByYh1wttq9r6no+UGr
vmnZteqTIm5UOFQGOB+SW3aUEH90vmAmj7rokDmvjK6ORtNEpWnTvKXxAy1fMW/G
NU1/0EklqpCKn4nx02dTk/xIzB9R7YcQW/ip7mUevtGQWniwqxUI+lZUIEVu1rjB
arpTe0n67TyD4M9FEBArin3aq4c0fl57jL9fQ1DI3agA0tte9UyCKE18K+yPwY6U
XH4YY5gAf1wN51ngx68lxFmAbF1WRXDPsaENw3O1y9jjhnHPyJr3GqbMmpxnjxNu
TsgaYDwEy7+AckicjiIg25YM06wiUOQNAjrF7uPmd/04J2NfdlQQTTo0kkuF/DOz
9vlrNBlqM6whUQhaBybpIf5MBGQe7OqJTY2nmKoR8ABB8p5iRy1yjWoMFcRZpIRv
LbATJNhXz1eOXbQP2h0k9NpkXcAXSe7DYmwom4m5ZeTp50qtUUz1sknhgzcX7Rwv
D3iEz1cokejAU+d7mgA1hglQFF+AzvF6Og5gT6EMaI6cYdCM5aBzgX0kAxyogwy1
1mNc7umzjsg738SAViPMhnF0S4x1hYTIwWjxvFBqIAnouXcksM61ERN6oAkHkKKC
TD0cIxhR4DL5H8yixOdYpGOgFH3KYTJDZVnr3nNU27d74FCeMPrAmKESqXioyoe5
KH6FUR7sYqF3PxB1IkdZtxYmCc3n8PEjkYbO2c86eszA5V63wM1SUxGPHo51vHzd
IlVwjLBLirqwYhG2OWpaNMAmDidC/Mx45NXDxWZlICexvn7uAG3mQtbQb/2dmZwL
XtkLcM8HS5rWZlSOHHexib42P4wapN3cP5r5OC2nwTzX4Sv4tO1h4TOa59Pcc3lU
Dj9c5c+vm4YDO21qO+tYi+XA7ZHptxQm2tZ+Hsp/Z22Y5FOBQ9AIethGJRg77DPG
XmjY7khZX+JDW3AfFAxDsRilCymW3fWi3hFO0XDFHHOXOFaHo2+4GbiYXQQdnB99
McPCz4tYMopyKW6gUVelJfx9xIox9XvAkjfG4SGzAcA008SB0Ztha3S3jvcLOByd
HCuYnVcJx3KYZmHie8wK/N7/qalLgH8MBuTCPFxDCMPMj6SmiCduVGz2yfrUmCcC
S54GH05TwK1uV575qdSSB9dGMmNlAOTkF7HL17SR6mRa+J53JTaFsjNfbAL6mP9o
16bo1ehi3LMaanJUpHj78GUs8sMehwxxSVIcpOVJoLQeYb9d1pGIbqrOZ/jLnNH0
XXARUMO3MLiYlCagG4pE4pk8+LXrkWYdFU/dyNpAZw7jciHgKW0kPoPwASQ8lZtr
BLP2MfJIMnxqbzqHzdGXzTsckPkghunhZHOoOPwj9CeP42FbnwKTvFp6N7QspxCh
g3ccw5IGXe8TIW4v0n6OULAwxv5txaqPSqIgTdiclMXDgaO8TGvBta7LwuPxrZjH
a4SjkulU0r5L5CIqwpMc59CjDxRwIT9r07l09nz0ejzJUN3vloskq5FIfFfdbUOE
TcLpRI2SA9yZRv/VCYPsdHUEl6PFDsXIpKKZ4bO3kbJUczk64IAJMNb9CJ1WYZ9e
6mtsk4ABKgT1GhZtLcD6mlwyH3pDhzN+qJEYSXovsRombfFLaIzVdU48fOoQv7vk
ErfvFEpLeHLhk2VV/SLzxCdqpz6HEdiUz6c2P2l12GBAlX9BAOozRvr0nZYsCYhD
5/YiMZ3Pi1lz4g13zpX/A+NmV+rNLMbBTzf4w+kYvKTSAgyUqMOM34sDeAQjDVoM
DlJTCMpZy+ZgmSovBTmaLIagNjBKDH8DqgLRpOZQEo984g+d/T5x3umKaT36CGp5
ljo8qmWoRPhdc2tCkd+phvHWoa3BBBNeI/o53MnSPOiqDTTZXC2msecFrUzJx2Rd
/Vs8VXJC6Omc1UPKfB+qS29m4yir63HCZcTlsAPDAT0k932rEqTj//ycHIBI5nxl
2bWOBe1HS79CtuNgdrNx0bDNs+Q9Z5cDwwfaA4FO82/OBemkHY5dacfhC9KqTouz
uPNvOdUIZueR0zxN3h9WclORCujnrq+3dQlfpWclu36xebJ2UHjnzSpE45tabxmK
oPwoT/kFq6QLglpPd5BX+8oTTfj6JhDMVXW/y+/SxrrJFxWq6hOxRby8MxAuWW/L
X7fcUj3wtdaUV3qsbEDvzvUtMVVFJDK5nZFsCDLe3M/FdnxWylElYI2H+ohtYQwp
F5Z65nKrT76xSpWMGlEjcXCUmslL8IeDXDRmA2rBYIqZZbcfA8cIMLVujBrIhq15
tlCbuv+m+kvyyV493PPpXyCUFNQMzC3QoDs7AhMZhKQadNvT40JEJUHjiBCfDxPr
sAzqj4bgVdfpp/VSfcNNiCgmJFXs6BUNjn4XbfTOVTidZgpSS4UvfEUdaggx4PxO
DE2OR1IR3ImfnQrDub2LAMS5wYm1vn62dtsJllbF7myddA8UoRNPoyaT0kMtj2kj
yzoXD7AIdCBBiWbl8YNmrqnSulGzZWbvCcewS70Dq11NhFNa8CUbmh+TPDlaxfoX
nvlGT32G2ErHeak8LUL5tGidq5NV4jCUCwuSvxHId+1rjtvnk/HuzYwZ2UYYEj+k
3W1M5iIG+gBUEfnqLTDlOZ0dfc8qG/dbOeV1GhgXnqKTW1//vyxGvWmx9YvBC2WD
TXBrxZSgkehv9QoVc8VF/bKNsqBq5w8/4YRAQtvIRQY6U6yzeGjjU0EJO2whCyRi
fOmU/YjjFs6qEZZm1NwJh8z/IwF987ptX8EOFX3Tlk7atO5Vxt4siI2uWtaqEkZn
PF5Qj1oVIBohtNfKaE5BH8vIY+megg88Yv6NaeZU9yBljVa75TtjgDhTO0SIR8XU
zRrF18qQV8luK0DZNDwnALxhW5cl+rY7F1Xotbhr+MsdHiQEebSiGF63F2fvFNat
uowAlPL111drOcvJVIG5upqMelJNKmUJphliEQSMFlLXqssWdEZRToTHHSzzkJpG
YTpBx4vshdFqC4qAjiOxKCbgF2wTVsq11I1DcsArVkjIZmHte6hH3cF1sku3luPU
QLGmEVmSY40qpDZBPWjFVvNJyr8Ih/9wbYMo3yPqO/yikC+x7/sPPa5RKysTDkDh
fazw6waOGK0n5ktqLgbVkUtvQsVsw5fZ0ACMZYR/za2fY64CM2INiJOF5rszA/Iu
gox0CCkqb+J3zqrTTcXeZqKT/EiTOvFGUaw/Dg4KbKlXuc0JI0r7ny+GN1cxyf3l
Yy/O+du7yzQMOQQS/gxbEhI1ZNbcjTVW11nVLaF4b0Okpy6+j46Zkeq8najv4Njl
2Bq5Yic2betlfmdxVu6FEVCpEO2x6GWolnHvKeuvo/OUTm8kN5qwPCJsw29at4Kn
bWovJewYOpksKh/PU9WrRyyFGds59oBmqeBNs9H/cs2Eq5UNtlo7Kd9BFh5Ye1Ds
l7dwWloHggx5ZGTWc58h1bIQ7LSWEr2EQxSr6lM/n+ctxrtN8qk4xzukxC4T8bCA
rrP8Qg+8/UK2HXs8KDVJ6IeC8TL69zx0ACgWnnN4PaBB68y2d2b7d6Sw7X4ehDuf
j3mwsGA8FTZPRK4C4GVWR4cQ39TXhPIT4Qi3dWs4l5YNsdsMtU1srYeI7i4vln9m
3ubcOxULV1n4fm73aLTZb4JnzSpftA//F3hAKvNyaoKLxG6Fs/mLJPk7pk6zpqSA
qK4RCIPIo8L4NmfOUqmgX1YgSKNDliVKDT+5ParIkFe5I15LsuylP2KB/II+SYoL
N5+V9GyTFR29kK7ocqJxl1kDTvoPtrfnl1lZNNK9lL60VHVnNTy2elW78TDeOTA9
swEv/FjKA1IUNv2pe+cvMQgMZLpqYamsD4UxMd6sSHeJD/mjlttERNt6n2D8Pv3b
6Hk5esjyI6aTB/SQqNFBtOQyqfqD9wxEDbWjjpr/NEqkQ6PFTECvTXJde2B0lKxw
BI3c+fXLYiWBA8kj72iQ0JcoqWcgh77otLzjmBUD+D52PJs8iJ9N+5IfJqMMn6U4
QlLUskWUMjL8Ky16xC3foyVVQ+qqPCY/l50t5FNwmbgS9/E1YpEvmKi1OrEocEyI
aPcaP/eohjQDgnuwppXv/qcsD1MZCINAFpafc4Rkbkj8kl6MMg7rHRKMM8Aj/ZOW
E8O7vlk5RabLoMlG4zSbH5WOqK9/jAa7CX+g9A8YVK2I0N80A/bwD/zkb9uQ1SFh
tQyC51jiJZEm4KtE+zdUVF4hCKuT/+6yroBqEnD2dcuozmouZKxr3UTe21IsARuY
lgNW0Og/JbqTm3of4goe9JP5Ii7JGXcJKJGIJswSwFEuMpPYeX1bAE7ApcBO95z/
8Gyl0n86+NJq8wPCXjmzjyfgxtyLKDZKXYK6IIKtSn3Bo99xSHD+Ujwe5xr+bmNZ
vMf1J64D5JvnlEHT6BN0EjPBwrDRd/YikVyOcY+fTBlfKpnnjZEf5ZM1+UlZf5Rq
kwNURf5dKY6cwogfpg4d8bCcTYu95HgiNCURoy3c/9iKkfEjNzjVfJafqKKciOvV
a5RU3MNtB2t4oHPlM0G9NiojFoads2qW0K4ir/47S61PkwDn8pzhjV9Y0we2SGDc
w796p1V7O2Uf5Nkd2cTZlayLdZgkt/17T5fwlu9Jw6i2FzuJ6fSCJyMcpTXKt00g
NiDb++d0++zlcolkY0KZpWO0Z1NJtuWY5voJDr8UQQ9T5m/qBTZn5iM/UPD8KBdn
2yL/ySJ1mc8RO5KY7H52Fc9BFrW3LHIyY2pxGiDEwGksQRenGpHIvv/hOGHTXYYO
jjIZgyJCaaVsIDG/qSJc3uhvH1kWAiUkiZrRpjDcE5s1RxiWxjdUijcbjUB5+qo/
9xxspA8lUXfLP3BHFsb0zXsxOSU2cWlK2Ba1VdG0iBrUlGE4uveCGntBgvycJfUr
5KCeSyEhjByHMZGaTG9vIpUUwvEZXcbTTPn/f4kaHny/K56+bIh9TX88eA0DoPZh
7FfbLgPtYjrBvSZeha5PYLn2enbGU1a5RkkWb4CWGsT8bYVc4leQ9dk+m1FIxeXI
n/GRX6RXe4DC1DmCMx6qhJRK9007XtD4I8uy0s0EsNK9rfHMg3IiSfuXkyWkbIOp
hh1W6s+UgsXLdzamc++JOgIwxWig0JcycGigDX2UWikUzsFLWDwVpBsPuEz+7UsP
NeZQxvxUEbU7PLpxp/53eO+kEFoz2EiGJo9XgRjOf1d8RenZeSM6Ffnerb84xmz/
+MvFs1ZqcifTXgE/NPZrh1N1sybUTmdMQXcIcIdKHEJz6aZMwjUjrH1YZHYV2e6X
AuFQyLVJ5Qt9sbgy8WpaLhzUXJ+u6OAVnATA6nDc31Bz6gekJPy+ph8N+TSupPp7
3cu8RyD12HtEoG5Z5RsIFccMkRFR7MvYNhvfMO4fJ3pO+vRHclkjfS9L0PRs64ZE
Fl3iHE2i+KgoTgcMRaDUo3c4TDdoSXGb0/aibVa0V+MEtmLLu4G6o1pSCslM5aX/
mr6plZgODX+FwK0Bn19Rgs7ii8eNfoevyqq+2Q0l3Ekvm9k3pBZpX8/hCTmoStdF
eMyBmFNJ0SAv0NZtwa6XcFR3Bm2cxsczzlpM6zxzo5ZSLXvDVLJ27NPSzxw2jOZ6
UiPIsS8ZmQ+b7mDG7mf+llen5LAsHXHOrQtc+8oI8SESMxVUmDdYny3bE89rWg/3
/w2aJmS6G0fJN51nuA/YC+faPcJK/VFu8CnP7+Gj2oMG3gboessXLWGnuUKHXdsY
qFJbWj20Hx7RtXe1uJtZrJi0+wvbqI+nNsTMCKXzacwfpQDO7bhg+5lbpA7MOdZe
1FxpSgGDGVXgzlQdG8OtYjYxK5HKuDYzSSTuB+P/Nq5YHopAOmUJrY+0tWgyOkqY
Kdcr2jMJ93+Y64pa2J+JdyIs2k8CkVcp7uBDXpZCrC9GlLQqcnvXSGJc2AQgCzb0
VIbWEESNzAL7JnpT6gMhXXjHfypyQCmKmumjfNZeKfdN8of7FtlLyVmOuxL76vvx
+aA0mcEYGpt2KaOH1wT+9+/1LsBrl19WyaWWnTVW5Ye/IpxsTEPRFTO+j4ivr/Eh
OJk15PIdKRoq7/7JXhMiQCrhQ4wIxoS1RyVVY1OTVxQxjLVj5snq+e5LTnfJVGxt
TRXfjhPvv589uCvD3HBkiWw/2/A5tWL9V0rHfRiZHr2/TkKiccEtStPJjmPQttHa
N2EHDNhEshNcJAusle0Y7vaKg5c5JFqt1CjvxRchT+1aLctVCdE8fb4hNZNXJkUN
dSzcdPx7UD3VYGPuHcHNCMKqRBfaaMpIdExY7uXSPXBf0tAmmwz2YFUJApgtkQ/5
md+2CSPCwR5nLD/3ZEGJVP3cFCIm72xgPC332U+rguOXvwW+5RmAaIf4eEk69vwp
Y3aqcuLzWCRtkj6Wavla0TsKxaVeGFZ83ymWaFFFzQSJa+ArjgJZKDbPupcy6Pse
YGK6KA6e9LDh0OjKKO4XKfPumpzaW+TC4Oe+7U+Qs+THA5nWo7keZYlHpWC8GT8u
SY4tmReD60Ntvw9RSGtxqCDskwdII8IGcVQheb1TlqOpPznqIkEi0Bs2fIE5fEui
TFeUiFqhCvMIFwdLzWg70W9LtQN1df0vuktxDTTJIfhzd5zN5huW8PAAXHUDIb9X
R9gNXK4hPwUo3knmGo8MtZaXvdi4c+Jx1Q5b+Q+xKYhpY+wLp8FZ/B1HQl9+lXUs
UooVzP5wkuSuwMIa1HkaGOoBGdTC6PTaFRqzGGmAvmnQoc+3COiQJPTk0pNJEY1o
fTRqVPQ4IYNGht8LUBGR0/1rXUCRe/smeAMBPh4Npiq/2CqncXIfMcQzY4KPH6q9
DGCaagE3n13ML4Hti+AXQScGgL1btagpiFMNjQyHw+2RY4vLXxoG8JVG+uHk+LMh
NNjZVuqppXd/h80TX2fHBuedRzPCxECpc5BHsnhBfQTlapEO+YQfQVBk4ubADNTt
1dBFwNEtPf02X0a0FmDg8FTy/D0aJM5fF2z4xT7YQLulW7oyKi1xXKZ31fjq0RZT
AlrOZQbUN5bcU0ySH4nOvjdzKIBAnz6tYbeFeu0mhvp8X+oXWDJBUYRkNtVywg8H
AF2q5DdoicH+bJ7jRFGy9GPkHfcAqF3jd9VsSvecOk0Q/lncfDSEoxuoUOb+qMaj
TGo3+pfNLkcFVmyo2XRQ3S9T+xRiYDPuXbjdHQfhZgub61RqwH7hHAEIj2bw4aru
dg8QBulD/5bH3+5T0loJYeEO5gMh/V6B9S03vDnh598sgSPUbUdF0zGjTdcr86QY
DdjJ25xyrNLfXBtjBok238tGtFCnTD6gTfLc7SopLUfy/jF4zxpxwiTWV+8YTrGx
T3GCq9XzJ8T9pDG1sYbB+2B7HTjFaGfOXK+BxJ8V6HKxSMESXCRG1YsEj8nP1G+d
DG99Af0+fe33MzJwTYhTnWQA8DlLqVaCwDSMlF+czR5MiyKN5cTGiBE0+eAcwgaC
NeKM5f8gQvk2MQkN/LCjtkj4he9J61FCvK1S0DkDARX7DEJIdusQVNKn6BePMK4Q
YL7ltWkhhkouLwYoFTzziqGglDq+R0GaOsQUHPlVhZe94QM/81ujGhzhxTr1GivC
Ei5o6T/SFNwNnkdms97DgDufEieh0xbboHREi0Vwv3EZG3aYdZ7PGB2bSK0r8hFF
TlXpQsBB7+1llEQfEcFHIPSy47PdTgoTnzv6yEXaDHxMBFInU78608j3k03W9FTI
ABlLlJx5S1KZHsE+K4qc7iKmAyYHboHRM1w2NqRIXbqn+IdE6mEEQ2eoMX4cC30k
cFA5dLC7hCQSJZzVbdNFvl3dChv1+l+r5V6meOelOIwmAxGS2BX9Y7FUBQqKhvvS
zAH+2ZMF3P7XIk59V7DNHBCEfCyGZKY+HUKHn+zJA/kxs8prGiWll7/cEDyGh8zi
GF2royFXQjL8WRfuGPzrSxKXerN5F0UKz5pes5izZO8faVQhItaGpynQjqNgD53n
X471gS0XjtAGPG5tlUCWuSo4y4XX9yFFCyT01xuuuZnt1UL7dF3yMts86gpRSysz
/EdKfBrqq/YqqhSsgBeByKgsbg8n5cSTaKeDCepLSVogwa2J+3lgIspXUHJUI0zO
YQYtbTBp9rsXKiU5MuildQnczFbP1/+FH/xmwzbldpBT+/hFTfh3uLPWv+o8derK
4Oll8MYYVtFcxKzCvgddTBG4HA1Ri55otlTNJeRZu64xQIYI0kTnBJsbjYVQV7i5
WmRMXpkBSLbGf7OL+h05UQnBV3bGmNkhc7j8xaee98rITtob0lnUAu6KmrrJpJHM
0AGjQGeEhuh4MogL0ITVUbypS2UUxwB/4lK3BlPd7y4JcoLl6oP0JqdYp3ZR8PMc
CVOmErGNSJLK951aQ9R0Fs6yCCnDBMOw8cpra0FpHu+7YIX7WU+FFBrtS5CSHY3N
M9Lr7PLUxIBtgIuk7zBo41YDJ4L7ziElohrfSlxKzQmauvtAHrL4kl088FJlIKfc
ymqteiZal0Ycfve3UzfbBY+rAxDey7bzSv1V/v5ZvHDnW5Io873+ddRL0J7nwd8U
zZz4YmYsS3THcQwle/EoQlmqW+4F7/2Wa9GmjsTYnywixifG5aDdmHH5f0LN2poV
/3Gr9YPV8zbzWEao/5IHTYIBJCjgcKopx/OHUC+8KcQfVW9sj/YV+O5Cw9jCGr75
EOwLOZhM7cg0vvyydbhesqixUAdV9liroYCLLiKqINi4t9CouTLUEQtS96J6WC+V
ukCa/SQIgIcd/ZwAs+KgHqRQC/vyVlFr4SEYZX16vOns/ZKDiHblPi/XdoS0Mm4D
/QHl0rfrMcl4a4ZqXCVsOkmEDFd6ysU7CjA5gc2q/j/uz54LC68+iEytV9NTSleY
GqX72y/sLOynSOvnnvq7gG8XXbMtG6BZNAOmJ27h0OW4XjcOQxIt2iDndRTzgsTV
PMEQwmxvKxyaIjIuJUJ2iTjreBAd0ZENaWWWeVEbdrRavO9jxCI+8fbIrp2wanYK
5h3jSaP6bwU1W7NgtAyLI8LdFNxzCwJiFIVS+D8breCzGchzcIIn2SY1HOgMJ60/
wuTQ5cFb49w28ym1W2llkxBlQXKNcyNKYEaxM0c1/0uWRx9fSyfuF2iYP5Ai6Rfq
jse5Q58sK7a4/NWhUwuGQbl+RyckuBbqVPhS6bXPbbD4qZGtMS4hPAHYdxEF3af8
w88JraoE52Q4PF5mHkDLkbtsik0ODXY7W/x0m4HYPOiqCy8NEKM03/qAfoHhE4TR
G8wwh93BqLVmbiWr/xxkzmLheMVA0RKLz7ebHWu6/gTYVnfdApgO5clzboma2RBt
Nu5KyRSkDp91k62w2UCy3GYKYbPoiP1Nd0Ze6sYD2QVQO230H+sr0b16fH/iGbqi
Q3C1ofezOEZ65Bhgv4Lqc2SU8sWy7Etb1ElhzuEMKT0IztUM83TJfEvD6NhViJsN
JjbtrCrqYHG5bJOUoTWnAz1avdQbp83vCBeZ+Exo6OxCEI8HiyubSLL00Vk3d1R/
GLXBlfKHZ1YfDCG3Cg6mC6B8ejiM4+sAJIbznE3hxiy3l1eu6ZFeXteMddOEMpaB
UI5ef0r4HBLXeaoyGYzRX0J6GhTmYFb4dK3s8Qc+wkijTccMe8wihirRlpA8Ug4q
uyOxW10DbPxSyluuN9ULy01KLuZTIyo/b0EXOHO8dFd1mEoVBsmDZr2/N/u48uUp
P4OSjj6wjHpl3cAbgTnzY0gtRqndLvehdyqpBJglMMvx2Hib06xa0TEHcQOEMxP2
Vj13YW3kRoUvKkaBbWF2xRLysfiHtlvz9xtOcgsaGLCQ0aWgor5ai5h2b9Z0BTOI
xR4Bg5LBGZtHrz183kXlSapfduCk3v14vhMC3NDY/4JAllRqfUhjWlV+ENMlvE3a
vjge/iBCuYARuPJ6GQ4aReylQNRLBhUIWt/QE++SmIKWCwGx8XbimoBV9MGSt3Mn
ue2QsI1LWSGsyFxR7BpOsoQMDwGRSxH+XU/sZcV8z5euqveK5xmJO4WHgAzcyVYa
OnZ87yY5JdMg510Oqgku3CtIGV8TIoBt1xZ7sxUY5OuoB2F9OQIHxEZkOiD3GNPE
uT9VzeCsdoSHtewh39HGdp+QeXaQU0FYqiM9/0WeTNsOr7Cdw0pQ+BaBFfSdrgx7
4zZFj4EjTtbbRNO5hUtJ0z64tEcG6u2cUsQpU3tVGIVr+Ek5FbUXTGpLhAmj0rDV
+w4tmHoFZnAK+GwfLdeCdCXfXxewp7Zwyc6XQUMtADJEApfh/ESiUz1222BmsmiQ
+V6vuJ/YmfJH7rGXKMwejHsNo+m5vnF560shqjPRrMn8Xp2hD9xWje5a2iw/nl0H
wUAXL3JalGHdSgxdHWZwAIcTkHv/ND+H9pPHESop5Pvm/Z5qo5gO4liP1NSLeh6r
LjLoRLh5fu8w8G7iJls/wb5XloB5Y6L1TQwAYZhLvXJhyUSEox2aNzXmaIWMT7VE
76HwtJ/6UhcDQEqYtvpIGwpEITUzyfX4RXbP9KnmYIyCZlEovfLE7yv8StjEyxDY
Gd7gw9/YfELBFBI8Fn/NlKQVsc6hBW3yiC0BwxFl3rx6Z/B848uV8D+zK0/5fPEw
U0NQC8UaeOtPG85R47eRhrWW5rAvbSdVlxk1P1q4yw2lASBnxnwNhOkInXU3s0bL
GvIllJQd2EfX0F8OqdnQJXV0Pr0U7DL27wjP8yuyMVUozZRh4vBg2OsV/o5O/e/2
BDuwH+12NhPKvg4+0D/XWYxOeuFfhzuKwxV/M85oJUace9gmQ626uW+eTrst5r4z
vH277N5ZZJJLbH0Fgxncx5GNHKhxnnqPy4K6j1ONqofW2mvPrbB1U2imLaNfgwE1
/dCPB/vGLv3fPFXcS/Ar1am5gkcbbgDZrYj+AUigNy+2i206ZTuoe3QIH5qHpAtZ
FsXzITldNgKO9OO1+xW5nLC/9YgFO4w3yb4DcSEsdOXUyuzW6UvPF/W9N0TxYvAp
xWmVRUIQyxdXQ61gmiurod4nlH8iNw1m/9vFjnNDICC4nRVLmxBe2imf/vEXXwbN
RuR8sdf5B4M4QHUYudA4QaOp1wjhxfjv7QahQ89VJdxsaq4HCUrqQI0STgcslUOJ
37NxjCcWHHhocKi3Rji33UB11uqhaSf8m+sxzpkyAj1C1WzNeibSRZAs9zZbSp0M
HPslPxvdVJId8LUEYz3ph0wv0XNmvNz3NAJvif06PAPY1xPi6f5E7Hqfsw+A5PAC
Niv+mmXr9PC4HQAbrMNIzU95sGZlGQ8ehqlorAd2c9etZeQFXzb2gagN+WiKZSGX
4Q+9O1MHp8qi779QazDU7J64PYTSmhG9Fh/glP9hs/eKp61jfnzr07sZOcUgNb7l
pglrJRlM8r/b0QikxVNwsQ2aH5DwscDCvDMUde5W8sSrPlfYbJ2kHelTTZfYfAgx
jKkM22N64zfU2U68BVT+YU5ADhXe58pdp7iG2ib8yiiYxtcy5+aXc+AGSfrZ0Prd
tOFRFM2AA80IfGr+jmvhSe0WOWjGqoYU4WWkxtjfq/cWSFu/j94yqscDYeH5hI7t
aBitOK5wtHFHpKmWod98H53Wd/6kSzJbpg5CcdYeGV64bhcmWFL0hdhTECNfads6
X/DG8Y+M4l1ZnYmYNH0dt/WhmXj4pB338K99jSHGJakW3NXyCzjh+hQ6hZ3h0M06
GhPncVtm9jbNF6PaLQadr1/3SLE7FR/m3kgRWnkEbK16KbMIWEUIWd6vm1I4Y6z9
NJ88efan8T7APBWKwMehU1NRuLhSNd4r23VjP6nEdW4lXLf2lSnyKDjnI/mKXPjS
ir2Q7QO4dmZx8a4m0DguCZfEZMnfSWm+A+RpAG5WT107TZHxT0snoGoBtvjCGTcH
hXsZNfie7YMDumstpm7jJOMlvKoOXpRAxp1T80ADGOqeiYkCvWp/Hk0EkmSd7aVx
njtDUIj9vsORho7nRJHroVbG0lRPs0I908uzyFigKBxLEkcidL4vapEQ5waDJsi9
TkQRA8KJfH01RnX9gg8+/90Iv42E5svyXrh2y73lU/EnWmwZ4HmMiIXi66Z4YNu9
n34erLJzNQqrVJZZrK25WhqGiRqvB2ORilJMEDhEc+pYX6kioUBTsH/FE5zrGmlt
zZI8L0Lc+RG7WEdAUOw0TWFyM/NQnXy4sUDDUw4otHT+lSS73fCmxiEcVe8WCLSW
SfGw6Ay8pECb9kUV889JOn8M1M+zZAO7fyJvyas0zIz6pv4QrTI5qxwIzNo+P7Ld
Bxx5JEmpfLzadaYwThLGCy5milLbFQWHyBj3SzYRojy6lijhyHGW24wyH2FQQhKr
ERUgerB3LkEyMw9G1ccualQD0Jz4SNiFoHE6Uqir/YZPBhxwz6NlcndWFdO36NMW
ktNgsfvmn6/eVi3a/NQrFCm1b0KuntEYhc442H9IpJqkdefwslSwDklaSIGnvIDx
QjwEInGghuRZUHbC4lxfK+i1ZX6CTLJNnuZ9eWYxrLyS6TRttONx1eriwwlWlRYT
bse9RtVVFxpVsEsPek2D1vbtDX6FMyjZSDPPLq2qQEvytsPVljiDH09kc286hv8t
arSwpU0M10Pu6mo6eEnKLFFE1o5d06LMvHrGa7bkddEgOzMPKqXDbNLRq6d1sLD9
rPZM1G1iyKJOvRR4cUz3tST1ZNXhzX+QdxVbbtXI5jtvPs7N90Q1ay0M98Li2Oo3
M0lTqAS56AaF3UJSgpgsLODSRBwHwAGeS0qrko96l41I8glRczBV3JyH167kUkTP
PmRrO6YsTtnHMZ3f+Pv0IVmzlSSJz1T/qGpJ18kK3hO1eP4LnO5FnyfEVUh+ru/9
0vl0bDxae6+6Nb1zerd1iGPWub1D83pvY58+8aRsAbF8PR4qkrwMfaOXC0RBL1No
67T2XfCWRP5YLxK9BNIOdUHx6ToXOaE1eZilGqFCYjQxTaxrVSrztCUNp7G7H1mQ
dxvlILfqWWnun5BbhryL3T/S9IXVWpk0eGAX8DYSHOTgDnwrv9V3YAtcI/OgjXaH
y+CAtsqWVoOQcI4e0TtuyS17e+o58xIb0AOot4bwf15TzniufTCXxT/wFuMbgYhp
ph+TWgaZ4PhvP+IhhRoRoKcIytbNHxug5EW5UoPjRunvBUjkbNQqlecqiQlv1eD9
nhu3IEACc4QfsUqfHstNDcnarW5vr5Qlh4XvpuU/ieOi20wmgti49x5qgbDTs3E+
NB/pjnCSIezkZZQwVMzGoXa2XgENNHOmSTAFlgepVgt29oi6Ag7gf/L+MHpBpVaT
3r4ih9jNcdFZZVpI5Lvasf0eAzIcXAYDLe/jdMzWgVBddOKfVy8hMCulQa+tSIa6
dZ7l+4sBT0Te7FhDII3qf7K+U6Z1lcld3azel26Prcca4EpTyFOa5T6QTEumLBTY
azmVGO6O52NNEHaRA4e+GRpU27TQGzCi9I1TgQEro23FKREGQNXPVxVRTqbX7gAA
LkESrG0VCGWmRnhKBmrFOGmlPogKO59/Mb8FwdnGmgkGg7fl1hdJwtkcs/xfJd1W
FY4+CHDi2JjZS412fY4qCoUF6c5HvOtF9H3G2mbUx82Oo3sOuxX+cS6KDIf8VSbe
S6rEYHVCV77gRxQOrbLbsh6I/DthR/kJn/tnZoWJWlwwp8+Bw/Li3GM9u1Tb07Xn
vDWdHAnaW8CCnivVzThbOGU4B9JiGgrzp7/Pz01fIl9XCvZpgr0k+ti4cvBEg/wt
93zd57GmrGdCiGvKK78WDgdiJp/qg8akOBEVORHLAApSA0GrjC7AVQPwAJtkvbAX
VKlG4BUawcqfbI2nkacbSW4+HFbor5g3fv8TDiqWRj4ztqP6Wrxt5QVcWk4hm1Ja
y8Vn856ylbuQBhwMd7oNNHDx+wqnTbPNztDKy6gkLIV51FoS1FA/Uz1dor2zrbWR
7GPgIUOtHrUpsqlylDlnVWLBa7BzpNCexmEtc2lB6cBqXlXkgjSWcejhGxKkZbU/
68Bs6Nl2pJZxLuLrvpTACggejisPUc2A86e1gNKbdtWSYSNWzH6Pw/jEsVsffs+p
X2doSYtj5AN/9Mi3+unOuw/nThVAKjQYAsMAngcjLrNcv6GmzAMQD3ff74cFmp4C
PDOY6y+TRez0DFrNQ4Du4Duna6fRIDJvqqWB1AtJForRuDBnLCI3oVR8i299Ny5j
fsTQmMI2/fUOVzw7BJEj4XAGjc/Ty/wDFw4P9L58fx9FxWGfmAALuAIM1c/itcnY
a2TVPjeDDo9VdxCxN/344QGPDsajK5cEqprqLaVk8ON+m1mzWXE0LOR5JnXAdvaZ
YQUCL4qBud/cHNd/CSrHElGSJZbBcUxqxG2fOk7aHoCXodqQjksFZK7FP91m4Ojt
iLqMEiBothwIdQAB5RMbpk2j2q1OUWyo1+xJmlT+iQJZ7EvjlfFFXsDdHcWsFVq1
tZOF2KKaTjge1DjSigVk0gvoI4c7URl/2ksYi5Yu93Mlan5lYRjD9S88PwcWfIZh
MzW9f1h3jBmIo+fNVgicIS02Kx3R+cMclD/m/zeqzMfzJKzjjof5/Q1n2FkIAVSh
WCyjJzNN3IJrlaf+2s1Q97syoowmeTh4fBGcsEkCLpMwqKy8aTd0ktz6HIrKkSj4
IO7XqeE4szCS1wacrR9TlD2GSUVGWPvoY7PXFIWnktc897SDlCee83twHFtEOZZc
NrMG2Nc/L1jDNdPQXgI9OPEY2L1dfVj9DWBT96H+Lpt2hAKqaWpUWEBOHDyMwXQc
4cM/2xAZDLnl8fW3wCUZ48rn0ycQAgQHmMh/OmGvgSbVhfuFj8+KoGSh3YFc2e04
87EkVPoZYs7JTbFCrrUs7zY/TqDLyJtMJ5WjwU8sp2BBzCFGBZUEdUhYIMJIEI1s
HQBo3mJ5nIK4Ha3xc1aH+3EOBe8NeeGLuURBFjheQAhdxhigwuFuYPxRpsH5bx59
hdwrbdeiPWGRI/h0i7cUZcbTXs7sEJFaH0dbsBlXmlZSufjX/IJnDQKtGAL27xGV
R3umQ7QnnHt1OMWab7jkN1Kj7C3IxDp2tAWvzW2kBzvvmn23SRd2SOhUrQfwJoFt
fHEx78N4md75i5Tzb2711jV2KLJU0Gbo0K70uLOPwtfNPoDYEg7nBDopzucJIb5J
GfxjAKImaWBumZYKuf7L2eQ+TLo5/0f6aw5N69Uuj2wUrJD3fgP+sTXNM0PiNJSq
1jgWpUc5K5s9eXJiudyoP/qeNNOgNAAS1qOCNhKmlcrpOLzWPXWafiGpTKuOuwJs
cIYellrTSc6mWtCGNP1UEm3mkvwYCSMIbF8b2mnoYvgVxoOhbx/6g+pIFgbP9TD5
Ia62QmUnc3PvObXoQ+5J7QgUqVmlwhDwpqHATL3JHgMR3ilp7fWQ4yHNQc0x9f+W
qg6U20XhdFIlLQhEwYE8XmYhkRQ3nhbeZd23bzBg5GZzOp/IFfgIfzEo4zrWt3sl
poaVV5/uAOGQ9KBN3b6P95NiyLB0T4ogW82byA9dCITNw4SJGpA9UMZMn9GgDTTF
/4OOg7jKCeQkJ9Ust1CFEfFSAtLZ+Z7XcKZO/xOG8dbh5MJoyWlRRxMDuJUQI8GF
QJwULKcjjFeCeWCEYJeim6q9v8QWOSh1mT56IIxZZfqryaD+gtNATIQhWXLE018k
2hnvSrreiOnXIY4NA/bKv/4R1eI101sqMThuXDn7JGpI+UdfxT1b4qg66TpCNkUl
vHaTp4h35MJp+ZBtJTiJ0NEmTNvii/z/UVU5jzQPQ3tP37dOELwcK8ayVo8RtBp6
TUh3UCl78sSwZfrIyhAercx/fZmBgDKSDOAkqTV84Ki0lqbfHnMjCC7Pp+oC6qKY
thTuBnqZBResRLDNwJKAfFPuZeZlyF3htWg7za1iAHxV2fARAGlm+6mhOunf1Kk1
gH3mTN4NCzcthVglBhXfld0j7cwAVN4QtO7odPXxc8eAiRbC+q6+CG+mE+ZKSqt6
9wFeVOfxTgN9BPOKId8UMsLgNSIseKQMw2OLQGQBFUHlCyqsJn7k/7QmwohtImC0
OOMcUa1pk3uXqUMLT9QhELgQ0aXxlVDSVgvY8JyhXZMf5iAZ3YItuSBt+62du2Qg
dqF5MG/4QyEZyeKAHTosphsxfXVSB0JdrNZwm7PEuM5ouBjLedyAKdsnnczf0+Pq
hiLRHdJGZN4t1lg7vfNElG6AuoSq/Mfw5xdKwkYtgqx8F0D927l6Jx1R/bFc6ICz
Kwtwi83NyESWXixdyyhq1jcOvx7pDyO1TxHcsExkC6WPh5DQ2IQxLdCnedqTgo9c
Fugr61hgYcvT3neXtEnVk70fhtdQnRIV+Is8XMR/dI2AoP5DDmxW8pwERu0NpfhD
brHVRBLIsQTsBt/MdQGR1ZrTET6h0DHyQzeKwt1vibssABN3Ydm6gM369QAA5kvS
GyAOeEcBcXNP4ddjSo+ZCyGqQ2TOnus9M3kDPDji6WcgVCXNfzS5bWJB3dKnVWIP
sO8v1vpwUVNeeIgAekJNKP4VHdW8TwJtoMK/XRbva7Q2Hyup8y33VdtOpKjYobye
izkAVEtCcrT/sNA6W//EsQsYYA2Cckl0NRqJTsh/nphL3IfDcGPsJhpQb2ojc9Kg
/8My1JxW/lvN2YwPQSzq3AiiDpL8uGnPJZXd2R+zZBWdGDxJCuwH4RBShxaZ6HrV
scsdSahdzqGKjL0cIzf9QY9hXRnCrZ4zo79gdkgtMwXYgMSMLyHj0KuVbwnExbIj
uQj0J0zpZ2fbnvWvxC4nu7dsoLZIfjgtJI4TfS6Em8APJLpnVnpVrGqhaw81dJVn
Hazq1PAdcGjShk/7b0f7ttZFJuOPcn9mD7LCL6b9HZMmvHO4Qy4LdTlRBHgdD4x1
m9BD0SyrcT2CJziWdf1KfjajZ67w54+Pn6g6sng6aSKu0PqM+5Vfp7ZaicCbuQRc
ybbvuWLaYerz2N4yEmVfEf4s6yqSxIi69HlZf38vnpJ3GIsSGwtYVkK5XsPpQKST
VkV9aOOvHUNf6mlpdgHBF2gEa/6LoEpB0ol8bjyV3YwhMuGGS8V9wZI//LYJI46c
9KXKzePgBQbtZBhRiexOsc/bmaTmN2kjg9Tr9eK+BPQtP6Do5UvX4VtR7iPqlSmh
SgbMt/72SzLRydLePAKSuWCcMnImHQ9nQ/D9cWmqdjA2nsvJPQUm3M7oWwBWSU7B
U830kf7htw8ux9eAKcRnQLUDMAJyDK9ezN4Jj7XZxw4SWqKzzjFr38kAoqaPF2Xk
Xj0NgNIZcDm3GiA1saQ+AQ2N2yPPJBS9hkXVC3g4OX43mfQ+0tL4fI9KIywC+B4u
+OdrE9ol+gXKQjO6WuEHH9GEd+9Cs09kxO9uBJjSzB/1xg4FRuNbjENfm/b02vDN
ZQX3FHNwJV/7sBUZAEVP899uZbj9nVKzlwtmCPMrAwD2HzWuvYsKKHx9w6Wj14/6
KBiFinfnYkyJvfk87EmvV5Ehfzmj6TQrI4cTabjGjZuIkFXAk1OI9IiK59F9tJ1v
7CeUYrksZhz/s7BrpGISoEbxqP+BdH0z4KbeiqRYuKgsEUqjVCCgcQM5ugcPwMit
A5LveploZsWfPnYqmGP+fAfE3XImHHIx8DHs8BaTOB2ZNBvzrT8vGBeYpPUvHKFs
wru57abJWxegJ3PIa4rZqSIIZzEKrxCb8rDeHHilIma9Hk4qVc6SBFx/YX1Q5U99
mECP3ihK0YOfHReE+LTfRk17swAzawOXP+5z5Vk4KKsAk6Z3Z5BHjBaShecYWn4m
g8iUd9pU3ugRk1JcBN1DqAGWDVMv8FlcPLjl+Mf/LEU+KucW9SRfmaccAnjePmD2
/BudyV1wGh16HdeMcboCIAIqcSl6Cf8zJ2aSYuNWSEkwslIkRuB+l3x7wRQTrzS8
x/fIXRLg49SJebqpxAJcy9sWWCDrHdC/uwXmQ5pkI+lpjEiy2wWWE4dpb1orZj4A
fW5JsZv/Y/CSqS/mZUHNvC5V80SgFhbX+i5W6/KlBffM8a5ui4rd4yGANG3kCtT9
y5LuEe+3CoTofhulRVyezZTRWLC0Rs60tkNcYN4TGlI6vjAwTyjtoEazebwrZK1Q
by2PeOo6SGzVs7GkurLLa1alaDMJt5lTzu3NX2eWciXEx/nN9rlH9tb6QAvhsq8x
F4PglnFPtDQoBPxa7uEnRm0yriESPxyQHMd2AoawHGvIQaSk1eeixRcRoHNGulzo
h4sdcghgE2cy/l8fVAsw2/0L7a62tE0STs1sNqkXk1+wcXhavzBG87p2/FlHioU4
3IemsTdSHZIYriVyxqwjjspm1IlS1Bu2anyB/PHI3GxKN3P6HZr+4+89Uwg/km7X
llKvtmg0bdPgRLoLGC4FSkh/uM6QiMyZeltKiWlqA0+cjiY/U50QQ19UippoXJM6
EK9xBdQ6rMbLk9O5m6y1pbOXJ8guCv3IkjGs9KYBvdiYKtLDmlqtH3vmxwvB6Ijk
w/I+CbqZCoHWeFTEs/B85+X9UDZr54v4plSFrINK6skSi8yrmcorjuS5kiNa4sVk
+iAlClwK3SG1dQDybgzWFJjz6qMSqJi8N13o29PqHaxp3fhDyxuzWcrWjAvD+yRf
KM24owkwJ+87gXwWGUElP7UdlOqhtSaedhvPlXZW3U/iz2RTgFKKAY9h59YJSJBV
nK+OA13ERqS2ZKFSYFuTYaopOwzY2OWe6/7MX3FwSVzK7FLdy4WwH8IJbChymOQk
bO9JlQtjZvARzEWn3aKxHOW0EiIKtSQ3HmNTukTRmpoiCqzdRqei011jM610QnZj
izuWGs9sGQbS243kPBFbVAfx2IRHx+hqbZD4hCD3uqBJRaTw3AP6gf/eBwib6xvo
e8jN0BYUK4uErtJpybQeqUw9c3Re2r+dGN6kDMNds4ISIjbUkwVLsvubg+PclisT
NNk3ehe7Qd3Wi2D7UH+2t7GHi1AYzRhMLLjw0gRYQ3jyPHB+it8/AD5vgyMN1jFO
xShfby71aR2v6nyIWI9DPryHRetu6IYCP4WfX43o7IC5QZj7i3opxrqavvq5HDq5
2E1PUiZaswsMBkcI/lu16AbSsteY6ctEA2Q2ZvB0L8uJpAMWbDidmaaQwlI2PCQA
wV/yDlnDUJUIb5EOdY/DYI8crjZkU/miN2cvSQ/qJHWGyGnLbBBz7l+MTJQ6tYCj
oIqJNvbcRKmAcMCxQr3975VxY9oPB/o7J/oWCqX+d2VOeiDhaYvFbBAAF9NLGT7Q
WMUlNrR1DEJlxxp1DgqajrwsBcar1c3L2U42lZ2Wvx0cvnizb2Q8SC6nwRo/vwc4
gWoJaNnuxZN7fKjd/3+px6UP7Gt8WaV9yDnn0oVrRgNg32PQzx5p/8ut2QWNO4h1
adJK2ItEw7DsZjRxJMpkilFf1acZrxoDzuVyojDht1qxJSRNOwy+18+M6aOM3cEv
/FJf2ooFj2+spPXuyQOsGT/TjGhqcJoSg6HEQkaPo6PBpc3ujsj7Z9HJgech7/LV
9taVfQZLco3AhXHWfHofQjQ34TfpPNlKZArhCKMTYKhhcoMs3M7jHvq4Mg0LkA12
WvIznRw7unJ740afhGkoUpdoVdgbV5dbTQp458y98GXlk7qzFoIBAuyVCkEpTQ50
qmwvzlc66zKDE0fe0eH6Q47gSzs2Dcwj8hp03lRTLb3vnSAfeiTkl1bKowiKgirB
D8RbKkZ08lxUH/Zl1bmlmdgplKHP4YzFJopmv5jrYUp4oMZmoR2wFyI7D0hPEaXd
gi6l1mi32pqsVnFGxpSU9AkPM9BPrxyqi42M0BG9dxYuQ7Qm/T8LzVYsqn9ezeHT
O9FW0G44mjySrx2O6WLS+mzwptfhKvSeyJgrzmQ+Uw8q4QdOUMbggqLY8H/mVmS0
2DLXrshVaERzw2gP9LBkDuFte1zv4MSjtyGECG873epZRTE/6ck6FJqKsUxh9ocp
pyAMt7K0BeLTBqMSX8P8wSpg6UkJ55CaBDLMnydll6DRlYbzAZrCURew43yRTYSA
JlDY8kAJwDNTJKE2mgMarOk1FM5h7hnTptuyQ6xkc2/8CNYtI/fRwpU3YiLXO+zi
XWJu3MqRywi3YPVeFOq2TG936pFms7zNoyqccHWnxkmNh7VZh+CibphbqdqExrAf
bqeja8fsiTQlhn1QGIXlnLuS28I0P1RFwlzSQkLu+rKjQk3KoalrML2ljpMxsZ6N
ZfG+XuMceWhH/eJ5qQWdFkb1Jjv4QIuZxlGhazFJVyfg9FxeOE5ElcrT9g2XYvcU
ic4JK6wLXKoTOjF/Wd02WKSE3VYvbea1X4BKSo7o8/ziVKUSm8VeeSK7qc0akG0f
E0VgYMV513Fc5Zt78tq8zZo2R0psnTsIGTp7TrxhuhhKHFzv5dl5bgISRTGkoVn3
TQ3Z+j/Yz61raoqfNMc1vPogZM1Ug5SDlGQdI+5OBka8UgoWpdYpmMgZAGMc6LrD
kOqV05mlcoguWmaIi50aHHwIqXB4D89VqiXGBq/7o4Ke92DbgHZ3/tN6fxDumUr1
Pf7jNvPwEPDNCHiEf1p1nETS2J39tU8bnwpmtGNAqp+yonBcOqgljSJdVcVqRdO+
4BjYts9OUPHGZAtMv1lj2EiHABiWK49elKYwpUzUdHU+eDywWmwwVWm6tigTwzIb
CxgIjBGsIB474fDapn4TY7eC5lzr9koNCFZavWhFjNc8E2qZwD3r0KgJRTMUqJO6
VEe7WBnFQUc9X8hPk61JD3XwO88n/UQTD7HBQs6mbcnLP04ydKBeyFNst6F7gFvc
2zPmuXdp7xy7oJtF2cM++Qar2yC2uICt1Bzi4PD2UyKpuMg+zNm5ZvQdO2bmesw+
uUqABa3MgwiP7EH7KoG8GMbPzUyxgSV4QZp0mbmUv7irZPLNKuA8sywq1GkuWN24
+T/UFhqA2Cl+jtxG8fOwTzSUHAehuPLmas/9SQG5+tkzVmYBiKU45CGBf3pJl+qo
/3gcS9RLcnhae9IpPJPIF6u7gYIVDjftRNV2kWQ3MJNigphC495kbdlJ3m8a/c8e
NFpcaRf+WxkexRFsvP2Aq7ds3aLCjkIrWqjYCRoDPMOIOtyX61+smq7BU7dCMKnZ
iKbq9yYihaT04oxpyT0iuGTPNscwNlKvNyEzzOmkOf9wt2nGSdbToZ8fuT4YYA7J
AZJAiBg8zfCa2X1Tw6mZx/jSSzZ+caElztsRFXhKT81GbsJU0f6PTC3AY462ewiO
LZOSGUYkJngp1IplmKkAK4smVhNJhGom4ZjH4Cy+vWkEAo3aspEi47lCysViPoCP
OBEOwf8lJF5njggOyrEbt5Ci7Yi4hmy8jxVmt4QC56LIjVH+tfSRESAzyVYNZNaC
QYYjqYf4ybF+yncsjKfTQNO7DdOnfAzm6yLKSGOQMHlGj9O7ZD1OVWCYCllruINw
4wS32UguatNmjWv8ELTjccYfTr8yrWiraVY9omuDfzF1UNi8BzIkG1EiOw8hzMvE
EXJfBXYtIH7PE56koxXdYXC5K+hSPh4W3R7rW5KK6T17AadYStcHuo3JH1p/HPAm
PrKaLR3SQxnfYGmuFB/AWi/lsLSGXr9G7LudycTjyFieZ7YRdgVBQYCIeBlfhIZd
z9ISMEtW0uOlojgX71ZB5PDlmxstrF+Y5JIy8kxGIFGLWIYOQ6pgI1sM5Mqy397D
DmRiTvBHQ8O4Kcy90mpFnUE/fWZldIEUQl9qdFfb1oi7xSAScQuGkDwDdl/8YAmZ
OnX3Mqvh+47EA9NvaxxJgPDOCNyOkuizd9fq8V9csvgYAMFs+i65g7gzG9nJ1wFm
mmsMfkv9zU47qU9RwRllos8+2AQroKtSFKA/q3F8Vx07aDm+7uc5HJfR7OnZvHKm
5E1J8ZHdLa1IJyqg/1swCXo44uUsxOqE7njunyxMEquB2MSWo4B0+ViJpqtJh75b
CxnaGkqNmgoSp3T70KvkqvtH4AGVEFzOvFeEXyLIiN81JsWw41hdQf8VibwkNJkE
WQjDkfvHHHGx5yOcJwn0qxdpL+EQVn52ZbD7cB5bY37WZodOS5YcYSLnDY4ULwwO
c4d7/jmCVcFayneiP/eYnqFOdDoVUxAQztp9An7CjGMbsDjeUsiD97f2kSfmO6I9
wmY4LaMsgxkcvbE4HGqiegSURqNznHYxXN5hpWVsLYI15PfJbcR6u2efQvukR0Tr
Fn298Hwx4cPM4fxJQH0Wqy6GwY0R9PHfv8iLsVZZuOZ8wAn1IHBw4528bKhobbmt
/Vi1ARyCvf2ely9ywmcQzd2bpWol1kFfmeL5ifMxDE0JDrYg3lPr726LMtaB1zSv
rfh/lfE7uAEIUQTJs3kDAOhyGOjCFhN5xytrHRGwOZqvkV51Mh/YblmPMHAoJneR
skULDv1UdAYe6AuwnXEkYm36Zh1mY3+VQKmnYFNeX4ljDjnyNVT+dcQB4TaSg/nS
mW8uULVZlbrbbr8KcaaAr9twhu2IQWGJkwaoP0fJSYuoRHNH7vq9fdCcolWCmXxB
I2hi21SvIfr2T5S9e3MAxA5cmGx8dbDYORNzglpCj2sbqKf2mXA/i9+NAid0rXZs
7nTn9WynzFr3NYc7eVLcHzFwraojM5+ahTHHGLOgANPymkx1b+APjCwxpLYziKKn
JRximo7o25jmCqT/1UKXgTY0f9FwizNS0wK9djDild+7fIwtD6rtwMq6BUW3/CIh
0aBIjAt/HegSeQdzkS+Ukzsp8K7/gQv6aqje/hkCQNoEa86pYpAfs9EiahMd6i1P
eFy8ToTDquey8v5TPb2vfmqZXiduyY96Sb+YFJYxLaIVI2A7h7/2T0KxxOAJzL9K
8ExNNgsE5ANS8jl7HFKMq1AZ1Eq8U7an8ABbCzzgXfXiv25gIYiKcPg3raYFHKsp
GrAjAwSVglsaS/3V+y1wPVcu/NCbc9yjp2Uiy7wBx5kIVrL/3uOPYVCnx3uFJq7H
BOYMV6GJVh2rfW6qPU+N/9CI4NPCB5Z1/6SKsHRmw1LAl1YwhTkI7LjxMzwL4xBN
/K94T7Fe/0f8KMeldyYjb1M0jm0YHjhyVJHeVvXnXHjHaKtf9P0j0TnXHXK5jtn+
XpLWjr+g4SoVRbO/3hoBfn7VP1eOY3q5t3kMP7GVMu+eArJj17O4qfzPoRRmzLtZ
r2Jv7oBlM+weSRyfKNV88Un28SOqET8cXKuIn7uKuYoxCMe6oHcDrPqp8IQVTxsC
RtYT8I1MIUw87uM4VBMGONtrqroKn1eiHtTbZLGxwtceli4LvEs/vU9JOFrdGJGF
22ydYeXRMTyiJaoze1vkpnA673uJ97fcX/I9zooAW/BW05te7w/OKX1fQxp7MUrZ
baTyOhvF/yJjxH5S9gXVinATl9ywfC8aL4QfizQ1jVJnMNAf6RpJ4SQDX/TEQH1G
QWPsCHSQRXf/VUfhUdEWmwbGZe1XhuJ9Q0d9V0QErO1nvJOH2QyhxlOcSM2q9xjs
NYi8DibczkTVc5U4mKWUXVUA4WylcdUBFzl7kY6z1qfm1awaHsQ7Jh1OFDwW8Rec
R8UpiM06NW7fz83Vhsuzq1MmkkDxcK0mOfje2XRAlyTdyqwVJb6TobK5N4TVty9N
w5XX7osSw9NhD55uszuGFaMhGpI40R9n7Cy/Q9+ECp+f/zXBWJXQdwgipJd8ymvG
NSL/l6rLEl4/Xmj3a+KbH21uU19GSYlhqjQ5LBmstWoKHaW9FKxNjCD3LP91gw9E
jSDfQ7ordoNSeGXWs16tPHsUIM4efy6+jwbQKT5Fuv70vzYzlTYNBLX6EP0CNruM
Eo9sfDI+JsYrLXDXufFqfjPWJHGMsHjTJLwKQeuytwFwFDmyVh088gvwthrQuWDp
RgpLU+5ftgZLX/BGxMRIYEdsqeXypvjtocsZAs1RvlyX5446LgkWpsrfVW2Um/Qw
KDjaYGZfeTrj44XBardoFshhdsoHfE3Sj+pAHUZJ1vRMP4cs7nspLJpHz9ctU3Eb
fPksvBdR+A1WvJc0UavxPHOIgYxIoFRh/ORgMDadIy4wdhGW/ju76Nl6nx4+hVFv
dCARFOG9vkIBpNLEPJ5JUkpIX1BA8DDpHjKC6O5yTjFxaOURB1LIXA6QTsDrF1hx
7gO+N2S3bT1GKxzkE7MycK+lMo9JZDMOHn5ZllTRbBY1QW/tnu+ZRYCeHVFTygO9
+h9lFhonWEAHvOTekaWWD+o90LBBwfk/DE7mMAgQO+VYlRQHutqSFquJzJrKQjwF
QptHLhHOIULE4UZCUGDQ2Ow7lMXvmyqdoyp8YNJL/08MC3eiQjpwGAFg2ffzGZ/D
daUimnGvJ+DR+5kuJOXtu7/LlcjaGvUjik87ie6Z835Hw3CRBH4lLRfMbjmnWgHv
96JbLhSgEHI+DVbfZFvzvL+5PXvzRovUmHw1x0uIPeDjluFhM2jXlX16vdl/gCLj
v3rQCn2hsx+JeerlPRLWmUN6E2bob/ppfHMVX2e23E8X0DZYsD+qRPsDdtpASQqJ
UQztvcC120Wk8fZWkY2npSalhILWQwW/239K/4AmHY6VSYGdca+3DXrlbNKEETMv
cVuv90zEemivPCaV0Ges+uOViH1alj5rqRc8nPlJ9BAzmvTsrm0kb5LGm4GRe25/
+RQX+ZoysOgYj3X7WiEWLh+k7J/i5glGCMM90b2469jM2D43aHY5lYstTicOTvoY
fdZ5S1s0SmSaJ9qx7YHUp480e3zNWE0pMD6No1ePF7qgSwjHSiHXB5h2GXD+TvTw
PUWLGgMwhhoS3NMOzkpIVE2/m6gO0Rm+ofzRSUzea2dK3Y7p3HWu9gtZIJwhR7+L
r6Ke/fBdE1fFoyC56S0NxmOkXAySYfkNhcpYSybSYg5E3zGg+sb+wmpv+3s0nv03
ax/3bqXmb4plc4Tl2WfrzbVcUjZN8CFQBOHOwHP57WPrDJizkvL1diHhpVrUNEiS
aJgW9SEwbwYHv7FyUmV8HssvFVI5OTcLotk6H07tg2/Q7nPowTKLbLXkh7Jnekxn
EHWwetMZl03AhFwQZEOxS50HoV3AKkyOP9UwLemC/a41yieCoJA+KBP0Sl6M/wOq
01nPwg8Ikb7LsK0/BFSl1zxGlEjOSXd3xcEZrj/tvwzka3NdRf0FCYbisYSqnGib
FLvb+hd/pK74mUeaLNwsIbxCreQeGBniEc4yCWQfaihlIEJklT0uJYrsew+CZJbv
vXMv/ESgPzm8jBbnNzhC0s/z9wofr3AHB8XCCgizk0SOF8KMMo+W0iSObQ69syqT
iXf7plY9zSvBkSdYPVZCahQIs/NpL77TfpSufLJRQ2vQlRn7cMIT8w0/Osqb7jli
xqzNR27nPlckxrW5YhWjjPt25o5GNpDnUHPGt/N+xepSFSi8jixAImjQfnUIdK4E
D8FOFIe438xlBO0aNrBab8A3LQce7kQmHSdW3w1u9/a3yxf18IvuNekdX7zLRsHz
5jRCdwpKYsp/kACeCLZB29wVWTLbF2yR9gAumG+nju9pSEOFSdKewUrIpurgnUiI
efeRONI4wIIybTPb0roZRTgF5XBa2pKv1tq45IFOTQ091TSI0KLpXpA7i1fmlil6
I3QfBYDBtGS8CqPEZ3mtxwkmsobmLhbM1UwvRV31O2BMqEo5Is/vbQ5QUPP27oro
SuQ4Zww5Pxyxzt5M8GmlIEeRZtnFQ1NgLsQ18Czo/wRyRQ/0YLcYO3ORynMEerAJ
HHgMCODu9FqDYey5G/xvieF7cZUlUhaW+uG6yCeYSB/nWFctfIE+UdUTIM2Clpzt
A8vWaLsL2bvCN6gjq2hXrMvXQuSpQI0wznSSJmh0ptXqmgjSZck/rI/oN5sbQ+Cq
/4ezvZZ5ahtEuqgWhagQfFhe8P2vT+oGcvLZiE+7scL7OIlS3bGml0er86wa3sYh
+pKyhao+U8+roYx4gZLCCsCCFgEe+Hs/AcQ9QkJYRgMf4JbTBEOIa6xVuNtcV+fI
n/1/Im5NnjbKnh4zqQqeKEoQExwYfnQy/juB5FkMapFK+moLz48nn5xenIEbaWJc
gbx6BLdI+mgHmPNpPIpCxbjULfaRA4UsTRhSVZaX8JwbHNWySH9THan6CN0n1Vvj
eLOUTzgcocdQKH+FC4RKWn8zaWjLxyYlrG4/S2YRxLOh0UI5mT1JQHy1XNj8ibsY
Onw57Uj3Kz8i7KyA1ArxZV2BWBVt07HIVaP3HFgczUG7jvEPkjpHRz7AkF428hWj
FEHPXzDs+4jy8nevxQO0Sl3hWX0dKflfdDOSYjO9ZrnfFATDAjEUUQYz8QzmibpE
4DGOT1I4mtsrS1PKRXJ5ejV+ip3TNqOJJ0Di+3c4IRDYeeGpcPPGhnGDJ5E0OEYS
IhmZgbwKdUL2IZSZ16J+JKTP36YNgAoof7uigKUsTisvk0a9ckij3jxmGORgZAIn
zBr6e8VIKOSQJ60oMYBU0EYTcVhQRrk3w1nlQ6aCrHQ9ZIHBbZISBQssWjuRiWDE
QFC5eNQwoOQ7DPAeO8TsOROrwELtFQRec5WaycMYUv/BJtJ3PXS6fQLmUM1+vJ/j
nARj6+28Eb3rYFTtRBcAPGVCjK31IsF1BlZG71wOGGQNpotBKdAZj/LUhaA1tUuO
cLrBDJ5doqeAzhBDNadO4hto5o7nHmLMlNkXUOZLRWc7N/FGkMnk2cbpiZuYa6Or
Ervw/EO0IPV4IHg0TaYcTzdrEGuYSYmiBSQYaLMTEQN7ushHtAmY78na1LwHIVY2
7MlL+VjTp0RvPHRU4busnT6aWz+FYytqygd5wDysBmanSntnybO+wHiZkAacqQUH
9OLBzQ0tql0RWBxsmgetkSiEtXgxGmH2iMc3eanfptsXocARtpPLJt1qfSHK6BI0
4WKW1z//enrWJ6R5AMiXH8/csD5ODvWrnhJ0fKVLLaZsFxlai5ftVAzl1HyUloT/
JPUPpweNMKwQj9LebRGq5f/1oHGzsUVmEuzDcdM23+a8qbvrktUeIPskecK0+x3R
fG/OLD9UVOTFWF+EP9MbiWVg+ROq4miGx8JeY4t4hNxri0GR/osMVWl20ZSv7mC3
lMeVwmp469YDtSGAazjb3zRkO4PMwaDSgAJ8QTqacdLho/oW5TH6Dua+Ql5oqEq4
w8KhlLEFanQHwJVcj3saziHepuqUaLS7dfGuWCNJ695Ds9FlvkDa8PU0duqg1GPO
EpsPiATBTJ2IB4zv7PQt/AofiR0CSoqL4NrUpcCW+pvTKTyjchI4GHSTrefCuEL9
b663qCpqAuAl+rY5XJD1fXEtwiW3WBL9eoGg4EfWPGBG9N4iRFD3kx5YwEB1vvQn
KB3Q1chqW/umekjaaSRdWnetst4hGMPNZ7XBt1S0q680fPRxSQnsIL7xgPM2yJ1Z
kcnWQ0glrF7DTNvkbngVWXhWX7Z/lOb7s3+fwftCBflprjwdnVsc8kmxkGWWGY4/
6+5dfbtnuXMoyq67Jh3lSIAxx5BrvQCYnLCZLL2c4KK2XhlWWfdyrfUrbd1Cr0Ge
NIzupweG6c2m4+YsNA9c6eLnRGMd1WQAwIJudQrQLZlnt3KmkKJiBFpAfucvfvOp
JsCQ5+imM4I+8Ufe24RoEkd30lstsrDiH770NqCSd/0s5IVfm6e5VkeMeaYMg1W8
Il+h2Z9qeEIbnR3PvG+yw+y+uNiIRYTIUBascI8zgLhmpo9r39SKyXc+rCy48eHs
SLcnKWnY8mD6Qz19x0AfH3iNwkBuDiXtIOmhLji4NwWDq1D5eKDtTLapoOQSz+6u
hVmmPt5ppjwtdIFwQQOp6l/isf0pmLKmOT83se5WRES+APqmUCrd0DLZ3mdGAlzG
mNPbffdVL4j9mnkaq5w8E4xvgiCbx6OxOhMp6fnR2biC/W8vlHzSU53nk+RuiUzk
QFanQvQPtXO9+jjYIEb0hAQln3EOkqVp/pCVWhz0PcwXp/YyT0TDhi8x+Wo+90kq
LEeaTofRo3YAEPzbQPBJ+tLMAJ6Xu1fcDLEhBxVEMYyeslgYhbqC6uGRiTPS1fKR
r6loh7iCzH2EJ2YCaXk7mEhrXXzXER33S9dUj0ClBFbfsssJimZE9UhM0Mwq1Jmg
y/eAihyRFxH0rHTLpDj/hOLTFgkGNwtpiEAFKqIwIoy/3cz0QEFt357ErdVGzTU6
cYXq1vNmoSCYVwd4lXkeSCaQK1/EwKII+VW2v8d3862WTewIaUoDhz3oQvJkUF6g
G0+h3ve0bRTusdBbAAYHb9kH3cgx5153pkvrGik+JYqqBReqzznyHptM0KkTSqxZ
oBHdXUIFBA2Bxjj7nnhOockLCu4JFPCnkML7j7T5yLiJHEkosuScgf8zZ8ozlMfv
OyrRwIE+kkq/xbBHYr4G54y2hB+p0TsZOBTcUQJFCik6rojcbTyXmyoFOO7B+H07
tjW452KUwRqyWlsGcGM1j+JFOcJQGH63c32HxTDA8s6vEPBUqZiKZWqhHtM9qa20
D5brWa3HlRmeBy14pDDWRjZQi6iNuap3Evz+GJKqHEHm6lDR9qxkLgsqtlh7CyYE
6KjU99I3WndGUNcH6b8g1/CXNO5V2JxBk9wMLm8fgyB2VoFA88OZpNd2qp9FHUrd
mGD1MpAEqpCnVIZ5ZbbN4LGLrTFPbtQrWPwbjRVMuTumP/7tQjhB8dUgdWCOVnsG
Q9KNb8pcBP8bIvkdD3et2922tbSCH+wV41Qu+nvqVc3MgcXPO/JVR9TiNkGhrUdF
s9wjuDUPlqRRBAJGQhEdwUsFhupqOPCjwGpav/Vr4ZeVHNd4mdMoThbKa/Gr7m/S
RstEgOUJ7kngivQGQWR6VQeaf2QYYGOkhBfA9zgOLCmcKDL9nb3on+wqG38cnrq2
asKM7/c99PGKWuM1XHIIr560vUl4P2WzxWixaWzS1oeUelpOIV9yrMyd4CSlmLBT
sQkFVjEP5D1Tn3tA4/LyS1kQlPptI5DPT2LXd9aGWDhOnuGW0+bNpvMkc7eJVhSt
BPzsRX5FA4PDtt5/HV/zhZEimi6cW237Ap8mZqBXCk6KEp0/gL1EaCLhiCCH1I6R
XGrCG1k+vsdTuglYdNHdYiAn0sAO960iR1S8MfZTKNEsiP3UfPcvtzYY2U8Na4mQ
UzaVrX9JHah5ja4gSbKoyxBNbE4WazXyUBHCIHKVjAFvgtMXx1/crmCXn4KTP1ju
NuWPEf8VZF/jtIlvnjtROTOeJJ1EiGGXaJuYt+vNX5Kw+2aibCzJzdAg3F9Sa2me
e5/Ic+CSou2ob88Mmao0CnM8xoFcnqnPrIu3wemrfp02GS3ik2i04X3iPm4NHIf9
2NuAYdDWE3DLUdEZWbarwt/fYfmqan81Iai7YfAWaz2/jzgnFnYPZXia21CWtAiK
cYDBhXvd8uJq+ZIo7269V7GNLcFaBQZjotJQBbJb8Yl2z0DNm9tEOGtEezYw3evX
nmc1kIB4/8Tm8Ln0EXiXGjgvKLK9E+W6b/YrZfoRsuoQzy+WGXfwRdt9UFzOF0w+
aUhLGLk/ux/z9UKTLRa6APpXHaGJnSVqFwK7zU0yHQq0O0OCXJJnFkQ5G/MC0dAX
hnn30afe/E7yqskwWA2BETc8YJyg3OQyMu4vdsVX7ZcNEDLTKMVWJB+FDpTu1t6C
fxhTKS/JIIaMOXlZUZQwe26SWEBDUXxY9ykpE/37vDhx/EHuv9clxzxbvPLUXI+I
3vOK2RdAGuXUMTtSHllKFhtW/9Auc6rd17Gau/Pet+GEK40IxPcq6wsNi632uBq2
K9qmRqWi8CBaaLU77wJ/p8m6nHTYPlNg4BWH/gEF8LFqPNFS242snuDNdFF0fge1
YMYDGyRYhp4tuZUtuYr0T5g3LzdYOJvniFAItkyRsKiVdzUmBAUro3btgtN0aDkU
YiFq3lB306M0xe1Dj0TTnD5ErcehdzZuNU5Yp1PPlnROFnBHbFskXxHNrH6vnru/
wyG0L/92jGpYxlWcnrbMrkL6HU4v133nElZt9kpVH9CgEDR3TIEfIbMzoIpkv88t
DsbVx+LhrUGaipSBU2voGEKPXHFSS4z08UYTEz9/eDROjVE/qXGsYA4wOvs4n9jm
WzsgNqLM0A1oMWlYvRd4HEOZskCYD3ZJs8o0LdQu8UNiqyPyC7d7hW2ddx02qHzQ
1E+FPb4S2zNptVyEgVRB6GW6KXlyRjl6ZKSIsp8m0OfWVTivr4gecorlOIvq2epY
27B0UzIYNqyPjQLXvxwJxUjp+dUbg9MFolyqHJG3s19peDa1xq8/dgCy1rM3Ekcq
fIlszHDWXJI1PiZMArrICK2+twVDn7ipSORdpeKJhOM0NASCV/s61ZUFhCb4Udbb
LHzmzGmEK32LdEWFNIzKSewUXsEaEtOXFpLG3NICvknvjRR+Ge3Id66tK4A1Zh7w
ib+WuEJoPTdlwSdf7XiXVb0T2fIyxFdM0KIEFMdN7jXBiviwZe2r5Dq85DvvNnaJ
qLmfzKxt9PoPM5EZ18t0C1/Sn6x8Us0K5gnJbVHDMCPzb7BpyY47CTTJf6Rf9N4X
jwJKMcb4s7BH2wnP73oufjoD8SEBjUmxvHBhMDaoF4Jf6Qg7hGa7KAIoDyF/yweR
oFjsLkvPPXlaJYg0UaJ+F33b59MiWe1bFk6Zt1BG4+cG42Gl+r5ENkHa62eCz1ji
XNXqnoYvjwK/aVDDkkbdwfmbhtvs6aL9t/ozXo5Xa4wOSBEZP8eprqUmsD/4maHB
9LgvZzCV+4slKLasc5Vrag/cUJYqrBngg+O6rOBK762ghawWnbjyNiRNr0F1Cuph
b1HkE9oZDbatdHQC3tZyy15kEmJjICXzWZES3jH7CvuNcZh/mvPbqBfFi9wJrhmF
v4kdH0D7E7nV7IUFvrqi2vw34KdHs/QjRXua9NY7ZbmhqgsvoOxqrItlReuPUjKg
kD47QDPC8y+k0PUmgv8WieFaHIu5P2tL+Sfo8iyNaOM5l2htgXM2EHuS0lBrwx02
ksw5ZzYlPlXX/m2/64PD6RWPC4VObRZReW9LGMh39pp3tJ6UfzuyCsoFIQWA//1I
xZX1OkNg1BD0bhLW52Pxfsxq9hx5Rb+1skfUfugxbP3f//bi7RLL7ouT+/7rugDi
mK56GAI9PtTmuOHOpMW4W+sZMu3SXKJgWyDnYIPUColZBJpoHNkwbE2WTM51sqqK
6JtwUTHls4gt05DoNauf3UgODN3NeemHqTPiukBpIU1eGuUxN7WOcLWY1moGqH1h
sj95jsSYjlz0lqVsHSUao/TmF2RAhyHOwHyLFzoFmqiCqJ7xQ6mQRNF5o/ahSAFa
F+/SogqyDWWB+G80ho5viRxmZkPnerQsnEYmT/sbQQlH7fNoUSKqwQ/1/JCfI1gs
IWz8M/L3E8l2XScibjZc8wm5IplCM15mCzhG7J1eRy/QSE/3Z61tCoO0h9hR3KYY
RYW/f83HX3B3+G8DSi2ta+jybelOmIt43jhRxwF+45uOfH0hcRntTPtO72bS6+Sy
PcXOu9gy+0jfb/TFqbItDi9rsTMMJ0ZrkCf1Wo9PROk+k4D8eRebbkW8vx4/IJ4s
7Ik6B+oRPt0ij4cOnL5XHuRuEYssxwd7We59EsENCuPPplpVDuMxCtNwZO7dbzBe
cPy70ZBt6YRvJXXd7yVSTYJ4swcsllhNMLMBKTvztcHK99ye9e96AWY1iIb4kDOC
q4ZIsXe6xaZ2Zn8ygh5O6rMraJrh/H8pIpEb5h6es0zpd8jbIXpoobkp5yx9jqHh
aRMzgyD/SMGHCG6llEe0HrvM7JBq66USRajtgoJzafBDXasYM/2fEFKS9wrFZge/
1ymzbB/eLLhDNG73MXQo/V7Yzc6++8EOL5SE7I8ZeVUNKEWVjwGTOmbgtchKbFdT
ZqjuSwbnP/yYT3Fky8Qz5ZRcgDpi6OtuJiE7JrUD8gz/1sh+tp3dLwGw2axV97wa
dWzyI/rKbaVmhVOdxLyAVFwaP65w0WCE+eSZzHjMH1GWqnsfX7dQSEEaeLE6SMiE
nlkuzRE1DhpOuivTndvZEFUovU5hrh26cTsMawoKCQPQTFJ2IA2oc0n4zMlyxZAZ
SDDcTg1Lrn9Pp7AgJyF3PRM3vZFEJNBIN3ihv52FwWTGqkaTyMUNxuNNPGfEzYPx
a9hI/ZkrYvnE6c1ZN7jJa9AUFSG0OpQWk5jpLEdJ+8PFMWqmmYzZxGjPuac7AsR7
fgo4hBvm0kiD7VOE25EsK6tj9+PS9EsQt4PDZr4idXwiPzJD4gK1pNVRj1cn6+RK
jVY9YsS60rmCPRQifH84eyppnLitILwRdjsxDfSMuZE4LTnY87S898CZOIuYMi/u
1679TplYLtRpheTq0y/q+5Sv5RvxBF6FzM2rzYmBWq3YfKFkCccKLb+26xYOtnfw
x4bFVrOgZZpycvAoPAE1QTeaQMN52xcSdi+8olDJdGSOUDmDdMkhYrk8Ul/DjzP8
UEreiDX830YmszMzJ2wPmRLwcuJhYe7Ve6vp1qNkQ1c7U1qG8G7RYluE6nvlpmhv
Xk4a6N+qttbMyLTyCkQGTqJEIFWMykEj9MgPZBv8GeljHJHQgM+V6S5qFfZS5/Yg
SkgTlVGv9+YmTn13OYiKdSOFU33JJZk1oxVNZkYXzFSMVcVM+3Xriz9BGNI99Fe5
OtJy0lQeCHjDUipRmGfAfE5qrHvPSeBU25L8TbVjwaYy1VdumuobjB3vcnn1FNyJ
SBDQ5I7sZnSE1UF5ikXoR37UYLTbueSTzZGiD7yUkiHnN26ne9UMNVitHhgyqpEE
OFRBEiRbLoXJISBJAIuTMYBqVkDv6jR9PIZXNJa8pRQx0MO8vTEXuLyBE0x+X4Wn
YwDAzduy1Ct8KXXhF6SME49/yug7Xw69lBYP9VcdKna9I0NWpe5O+zbjdicY24oV
Gq4JWkhhhEnIsthQss021q8yFeYZMVMYjLopCX+T0w5yFZXgXGYpdTqUgcRxOvHa
a1CatP9gUQKe5Cmb1JBAZhTVnYMhuh34XpPNr0QjjApVYYlDI15QWz1TMTF0vNCX
sEaYsISo9eSGgXqMwqYzHNN/cJDOfXU+xyB97L4csyNF+wtJuyP4i53RujQ1atW2
eIjSyw92pOM08KjiAexvHqtOa0KRcg0vBTNPkYFnYXmJvpdM1aTfufJ2elLwe2fA
XOcFKWy3DsOaI6f15pYXUi5XRBWou/2PK/yYRZy2v8E4a9yo/E0UFfeERYxEP7D8
PUjLZ947hvm0VsldWTF/YdA6FBw1WWhI0mv82PzBk94TBLrewIYs+YxNT1McQw+N
0c7UvXE1mPW9J51T2kxjCjg+w7+AnJkD6gZIh1QwnsXFoBi55Enl1dQ97TZPeCLE
WG02ooCQiIGbrururQF1k+nA/toZgEeu/8I9AsG1PztU4Up9LRiE0gJABSiwCZUL
JjutPJDUX7+rgyiaJc0hl4MKpJxZbjzi6Cq5QjKA3tlfgqcpmWL1THfB8U0VjXCn
OSrt6nC7Er22kI1HXiUnsqHxb9aXuHrZGTqOECN0rWeZjrlG2BKWxAE12QfFRYLm
hHWgEzNcOxh6H2RxKKdu3W58YxYpYATSvryAecEK3WhX5+mRnFQtfBN9QBv7y9SH
bKyBvrDREQWYpMyuenrBTXDJY9o4o+9hnB1+UdQp/gwC//UMkrYubX8N6mH6mo6R
Nw50dAKPbr9O0nSV4iQVdc+4W2/SMHZ7AGfDLxpU24RsvQd6LHWyGf8cDJ40Uat2
88GrYCIbNKkqRPh3M/pzWfGvLUZbQXpoYO6t6fPWOpZhSCBrEZuQL1gbjVsocBsE
3IXI317J3Ad5k3Fk66siNUui0zDVG3HD59yRm+wGqYQVLT8IldIAEzGwQdlm68w3
4yfLs2ZarhtQ6TUsY0Ra4PF1lpgT3yQ6VJJ2Eky8Ogl8Vznfs+7/Vh9jRO5XqvDf
yJK01UhsIJgC/UP7QcTYEOgiBRXercIxHDf9/8orfgzvf2ZFCA6TTg0E1NMiL6s1
qCYfYmYpxhaqIyxwBeTybTdXc25P1A0wb28ur3kPeSf4Fb0iPEfF3rCd4EE0CBvy
3FjkFmwhtsriAE17hnWL2u+h3WDyXNi2i97MKz5On255J1dA4bah3OSfN5nl2RBN
2hmd66xALdohlKx07zO4Y4P0HK8ZoXOnegrnOwexEh+4P5qTb1lDrEMRJTdy8V38
Wa2cxm/U2O1k4+qMcVOwevoBXXwj2w6/YzWm4CGmvPz/EO76Y9z1s5zhzsPIW2fS
fQF/BActd35n4V4tcnR80H+CK+hKX8XpdFnLHW0Qyu7jHqIFW+EoaO3tBYKXxLAu
eMm/OmHBK/NQjKtZFvggI6xzwY9Pdm/6l+etLh4GVgjW0mlD8JFUwQUXaZW7aHCT
/tfrKG8FoHTrfNPcNYXJzTZqvOey8wPjdtyscudAGdmBinJ29DFF3EuL+hoeGRaG
GGZvMugxZRRlfAz/JRwe2H6CWip2DudmFUoRSFuqilfLmGg400oHQD01eY/ap/qt
w/BYtHgUAdOlwu8wlXhdM0p/B0RT8XAdrvEKaaeD+dQx+/hddYVkh25T/zlC4iRf
WX2FnjxLiAF5YUxJuht7g8rZIFXzcM9f+ue44KiMNJHbczr6q2vA2WIVTHQc6PTF
Z245rUoyCOy3J7uHyUqhfWBRQh34UMENY5rGgxAd34YAu9vSZsBH2UTFF6uvAcNp
7KhNToJRh5p+C9yIlRn8KcDiQsdQfno0NAtSaGghaURNywSEWgzHvmRujGytu+F/
j5jPAY/rhjDRM7BB9mAD6c+Ppz50F3NbsRJMf1jIZzplRVD4Ov57Zww0m8Fukb5H
8a9aBfZUEXR4t4NebaeKdPdEc5AKizvZG/VamD+JQw1KlZEPW/VQbNDB+lCMSZhi
UavMLnzXEj0QGBxTHzTd868fnKRlSM8agvY0bcBbeZHsjiIOk+N1JIqLliB/0j8t
DQiRMMfgSXNiq3xENP0RT/OC0LnK+jR1l0j0yYQOEqMJ2ObJj4fk0S6yK349M7OZ
XLGX37rvEzPZKsCmLVVPDJgt1kCiZedCs+jSGrXQ8NYTFACIypj3hr1qwhBy9Zmg
11ezGpjWSTzE1Ph+ow82AclLZ9R8ZNuYhRuZlF0X6d+050BaoCRKENABh92716wO
utTzZppGZR5msrqSNieNrwULj/GATbNk+5l5+TMiH77aTScvs94c3phHZo3KTquJ
LIVmOJZmj59nbeqzzoFh9sFVVTAJVdrHTOZZ9F48VziifgDwaQrRSfY5L7Qy0LSX
/hX5aBw8l5pKz3ZZCwck1PnSd37zgmYIaJk6yHZ9CCuGwMQ48v2ljR6yeTZJDVFQ
3nFXp2VJgrnQ+v+YQAG1T1ocBV0rUo1mexxizfgJPBpyCBYNpp10JDyApJXTmLcq
fICzeBrzYr1AIF0CY2mRNyhtTsm5zSIvVghB1md1ZO/tqUzFFi3JvhCtMIiDai/x
bk+2KUO7BE8nHo0xCYWHuXFLwKZBHRMGW1aujU33V1tSgFzQ443C5uY9P1XyKkDg
wlOs7RPIkypRhtPIgHfwfYo4mF14W8AAaCNxLCox1aMbiexH0NfA6VBKhIvcrZP8
yhvikA3O3yi0Ay2OEF1fwiGBZ5V16naw5lGYM5yA0uRAwJqq4qIy1Ui34BTfHI9Y
AZZabVAAiPnETtYTwYTH4KY+Vkq3SNIuYFW7zzUpa/eH7daBBK4r3g8bY+KLjzJP
cADNSPdxeCfFFzZ7v3YFMBDJuNmFVpuEENuXI2NNatP8m/fm/ugobcFdQ/ezecGJ
aVCIciHjGnsvHEJMq6xxMeieVmI6hT6ePXmhBZPvJqusT3U2yTQF04yMLrPFLPB8
1dh/d8hrwHei7/Gza7dbjYb1WuBGgvSBqUyOI3nBMY8H/MYR+WrSRpaGJc/5V+eY
nGLiIHGsqS+mkG1x1R7ENOC2FAD8sZVcZQTO04tWAT/oUFs9aghe3S0RxpBsM6tF
asdqhYklvb2PIaeZ0Yn2rn9z6LMfngWOLK+RfgTEU1bVni2WiI0tMqAMscnM4GED
6JKpGrMtSNF656atDajKER7j9ndUFuyA4EEl5zUe7yiKO0xWtlh6PFgxcsW7S54v
VwG6FutXELxZcdlGE6h2sPOZi52V/pf7hTsEfPolr4VreyjZVt7DdqpuCE0nPu3v
q6WYUZXg/wlRpH/v+EZoBZDzOUB7o7iLSN5shNGsSPDVC/h8QEwLTO+ay3PzFaZw
3EsAPGQ0SsewEiEm6ezfAEWo535HmNHyz64gYWkLvOhKYZj0CpYTHv+axNugp4EV
jt09x/HbPDRmW9Ys8LZ2WWVGz+9IczWpA2iacWGfEThJ/kZ5joxMxnhitL0J4WwI
3S1Tarf8VCXQbnIEnK/u6JeMa5vo9guL3x7BmU3B/0qayegtZ0sVt9/wmqat8qcH
3HzZ+TRC4jzrTKp4rFFqkLMAeIE3bTLk/+4cOYmLkScQt+/BL/KmY9vTnB0yUMEB
2atvxOFg/iySzY0HgQ43e12y5hzxf/rgSPySI1kQEtBlPpPewz0dN1x2a0Ks3Cci
6OKTiIvfBz1UfDfAK0bGCmr/3FFY3sfXnEsVHsAlvM61Gp/MTYkIzw5klTCAtL6E
Rt1qQ6S0fgfkwIzfRnA9gQtlYulh6dK2WW5mGy0WJXMLCm55Ll1C/cgmJZWAvq2p
aCxQyfxikIpyS9zmR3qo/5uQK1JvTEuDb19mZeOfDLojL5wWq6xg0BnsBlDstmtE
jzcmvkG3vD5kuoBlxgcpytskKj0c3E3FjoxWeVo8IpqB2AQBFupOkH1/qOoTynrN
AaV2OVy+pP/1dTxLYqrZQ8wuoIcZxjhS2Q8Xx58mdVUPcsLfZAT8F13L09/t7iNj
ufiWnCLz+xcsL1iOKws99GTIh3etmndF1gkPOxnxtB+17/wVNnog/MiBjCtOu8SD
bAr8DeWPxaprfhAF5fPCVxiSkDRmIlBmCRZ9vo4j0fXJ6DVctEYOxKK+oI56hIrB
2QTaH+C2NRkQ5PMhYHUYls33bcExIm0NV7EcxK3Af1/CEP9pbPAO42qlsovW/MP4
t37c7Es0wRSLk+MPlU2/nAhCBi7VHmpvLWAKiPSbaV8GTRR4GKJn6eGK5uPPFYqX
iWL7vgapcJtFz9mZvXxFg2qBq7IamG4KYb76xr33f6QjEjZKL1DqZL4kvsbHf9QG
LPNEkUMOGP85ZSJAMWD1pue3gtMseJaHFde8Z9FYn5tW+FaZA02W6zo1IgSwetw7
3vcg28hU8+A14uYi5innRk9yestfXBYjVCWenOFnJRAli5BwgxzeaKKw4BuOQQRq
3wOVx265CH6TkZHiUtzTImJS44ldej2Xzw8IVqAAXZcS27phP/HDjzJzERm84ch1
5NdVoMJWirrVEs/IPGGLyHIM00x6LaCotvv+ihS3NJGgBmHA6yakyhwI/N3SRBpU
BXVekE/5tC/bB5mV6PclyqkcpSL6nPlqm/vAPvni8KhT8sL0vLXiZ4MvG4onQHwc
am8OznLOM5SdK3/B5x3kfHgZWsOgUREhjg2/6dw+qUFe553ypKiBdIcVUZjgoLWg
ZPatkF1JFlsad7uvzm7nEc8lapLIJCQNx1tZCuHHcV6lsa5uTkq1rT9SMqlGYyr3
oGV/AW/8LU6L1vhswaTO73bIzTGiOvtgjoSOCadmZzEahJfjoz0OBUaSHXQ2UOnX
M3qlLrqh8MRv/jLOTYs2KXPQrzW2jqiI5aDFavXjAUZOhliLnvY0EGpAxgGe3Bo6
apAOlbU+9hs+9Gf7P7V1QpTw9oqz8GwyU6WtokabJrG8soJhvDwIySfeP8Zhr7oh
pzyx3Rgi9fq2hxfKULnFzoab/xDujVYkiA+QtwhgduNPxLUZLSsMxTMCxVd6WrIk
+lp8Hc0IoeU1bGPocDXuLZAxfwvA0bsJSFb+uDtdbR8i94erbBsb5rL4er1E+QKn
JuZ28K7gBUWXFGlV2bOX5GW1dcmbgSSGyCYXWqVNrCr/AzV43MlnB6BZJF/4oqPU
f/jF5MwGQPpoajRPZLj3fv4qLuuv+JDFZMISIOIWnlcX0M0RcKIWA8ZmEWROZ/Re
FKRp/vHjL3kLnE0Sw61QFB4h/WIZlJajIseIMV1kR/fudlygNF2IkP4LKwe9F8+E
SHz8A9P47vCiQbtrqDGNHMLUnH6XMBGyZIvzZ/Jlfo5CjXW/8irSc33IJesF+7YD
R0ougQKkKIs6Jm9ix7zGvCXZlltSFMOIxe5dNDk5z8Wxvxff/d6M8TVKwamMbUsm
j5rCZXGGCqykiSRbCp54cQZ64kSanviY4ebQXyfl93uApVyEjWkloB3MXg8+fXV2
swy4viBCa4+f/Ml2z2jByTH+pgxHH89/2YYGzxU3hGqQa1sOEmVFIrZgh4VzxkvW
Y3GIKAL9wjS9RS5P/J8M9cMJLDBgCdYqISCdtGINbRdMjz7pJmj9gVt04yWQqp1r
eAKvUxL5Pc363CGpejOgQ1cwkrPqU9ejH1j7B1shqnm9vOFu/4YbOG3r0YsB5fqR
oxo56pdPXXj1cr1H4Z+aP7xVRAnjEdV9Cc6gCB2DShNm+Or1ogrNj5/yXq9wtFn/
a/IhSg3Ik9GJG8UpuMd3GPoGFaAtMW/+8TxpPWLmHgGlqqBACDygOo0SFSx8lAR/
scS9DHmlv9QJHfr0BnVcbG3+/Jt16qQi7dnlsC61ypKhMf7J3Sg3WMxhRRJZpmSn
fWZ4u4XGoORb1Qgdk27kcualEb1W1JHJRprNcOx1oDN8SgacepeV+OOubuAQgoTe
u8lJovgN46T7loIcFP40kjMSkkCWu7gn7kcMEb5erYgaCa5XVmJpICr/xlCpspi9
MgKwUAYK3c/hLvdXLvs/ChMBRepqb4inuKTiDx+U4yrRsSGnJinxfd4OhREvCrT6
K+gW1K/EPohTWRKXaC6kktYnTOLLJRniIjJ8I1AFwOjJDg5zIakojV3YReXxeKZR
GY9rpDe8HSzGRzVLAhaSkICbSniNdIMPVEzC4QyZWXBHTqy5f/Xvtx/j3jXNSnqD
sUkCPqmy25aEeTRPOgq19BFbzZvAZ4AkiXFiy0P7N2V3JFLbUnnlQE5yvw40urng
GTsFj6aewrtDqcXFCSlh6uAh79Vi/ssh1n1pvk+WrH1tYjHtbIQ/NUusQ0O+3sCF
G6ufbtOp7J8cR91VtNdH0C05nAq7dzM6gDQ03dbI3H7YsWrxlIbhNmz2FDHU/KWg
bGQIxNgOX0aLJg+ThHJ6KfW31RjRtAPRVnQ3zVkEZa43bdsuEnKvXCDyKecgLwMX
Z3L3VaTJB19vdz1bI5US7f4t+/Bcu8iThs/w5fyG6OgtG8P9xA803v9TlNaY32in
m/u9hOOUnFE7luW1elGdERtWlnTsj2Zkxs27bqSa7B0rp1u+WcnyDnSDbVlHu5gi
3IZWow6qLCQg2RZCdYVADPgXpT8m1DduE6TJaqIDCb7FwMMaqtB9W91uotZyEF4q
bJ7htQm5+T0C0oxaXdzZ6qIfuQpbdcNtojcdV89W0PBsHM0bSaJ/WCAqTPieKcoc
Ke5LqReRRip1XasGtE62+9kWPkYCZQm3NbTfYQXJjhgmXYtHFJCWeaDqlAgRHUUA
66H0Y/MuyASGakwqL62abKZPg56gvHnIPR/OBwYRsK30jhm22zVxutz8MqASPXj8
lzEDl73rIFljV7+BJt90M5Y49bxnoUr151lfANBPyfr1fxhkiyJ4QBe9pfpTYQeK
Eegl0KswzD6jJlaFNRfZvbPf0zKCOt3Nn5b5i2rRl/41ZgXfamXMV4p6c8rW+736
YAGripZRGhgJzsCRHoMWIbbQIcwcpLGHmpoBs0TL6jaVwRXyPFzoh/iw4dLXFyF+
h3oVWjlS9dm63Vr2HjRK3GAyYypVnFBvwJaFFIGsro4rcu9q0j5EBs5px566oONM
qC1MupOnkBEv9VoEVumLKIFXeNTMxzIAStvQjie++m3MfHneQ7etcALCDNP8nHWk
ssWDRDGygItlthVvCbPtYN3llGR48afabkZYMan5WZOwMRGotKfl/3vQFwzUzJ8X
vrDatScHBVbKpZSNw4oPLynZwPHickedB6GdByVMCmbuDqAoQPenXUTos2WgnULR
bTDhTOPvyTKd5cHJgH4mWGpiniYwkpotRoyGHCt3QTQhlixFBwHORFj0/ORufAAG
J+fJyfE8laqBz1i0Pa/jBC88kZTLBMSrYQdGyzlfex1Kp0KhqrkgGLgTzJRPQNNJ
YPTkbZZkFh2Qp1Dl0GlI/mO7EgMIwlomaPFpbWnz925JbQn60wy+P43tuTR/j+cH
/8fpJen7gQle3I5aABcBoqvDJGakZeeinrLQD2WRWrmkHr3skd9H1NF51dH9TsL/
1k1A636qvZZ/5TkdQMxFOjbNALFjYBjmZFpa3Ed2mS697btzqgKgvvusWZBfiDil
AIIvcTEXXZAUlD51ce5qu8fjl2F4rq2WgoCfI/kIpOmZtvu++mcO7jwHjZpdnzNr
B/MjCOXmp11Kc5jh/baSzFzWMwhQy51nqSsp+KhQnDeDAs9ZayCgVMAEIunWf//i
5NYFXJ195ZSD58FHhTqxn+3InVQlbQrwvxSbsNYbg6/NPbfPHmFDFNzWQqnJEy+Q
383aV1BirQ1o1tz5mUug5L1J50X85Car4Y9HBzHKLt+sS0u6/VbdMGcPY3AKwoSW
5qE4Lo77m0HzpGtak/ezK9X1/Sr/vGH4Uaw1uuu24ilwfTrfEIp0rqrPyE2lEogu
0J6qJBtNnpVfpmb/DFFmSVQOuMfMK7911X2WxCjxWXrz3ZyOV1g2P3iwTtm9C0+U
L0NiGUVI5r0k8Qq4Oeh1OiiKiFGOzNcg17b6ay8wYYiFiB8DIKocR9TswZJOiNwI
z+VbkP0Rbq6AaDi5qqDETcOqSkx+DzPwKU4TE/T7/wYMUZGK9XPVS2sB4bmvGllP
hgKsPJLV2SW3p7ANlj2ZH47hpjqXpPOCFALadbKSiJe89V996q4u6AoJZCJqN273
/5pPoqqCzASSeDty0vwKyZt0p59vMUYj+g8GuJwZ8iGR80Wjy0e/cif+swX+lzLL
vouQ+idOOtR65zwF44MJyj27Wzo2LBF4I44sbycu5kvOpWol5ib3p713jYu55REQ
obzeomm6XRKsJqkj1pNOAXTLMfxj0doHeGKeEHrYTCjUomuAknNwvpvPZsYjbD9Z
0Mtj4wYDp837KhiA3/GxqGG4EI0QBCb2o2jD4WyPFJMdDKQOuFT1T50+1d72k0xx
uDryMTojKLv4+Jft0oXd2YeQ8X2WPpKFR6N3TZkXWmi8PBeiQptJCAcPSoFpi7CL
ybof5JXXumIXBMkU5Ol8wIDrDuqVfzZGcSy/MQEzMjmFTUm8oS3UHVJdAqTZ/m8P
MFyThLwNUIH3b2jTCShbt4sXlGFBumjnWP7omevKAKUL2Aoc2F09eEJTYUYVKnz4
W3rrsqK3rfzAC74V7xJsI1klGIGk15G497CEHIejDOAyO46gqLn5sIWiYEpIl2Y2
o40/0TGu+Dmhb8JotBV7QPXcZuPlaKoKNN9TzpyXJR4+c6mMEzlxZtGBEg5HemG2
Ro2rKsAxlftGkAKXQjBrsbu8+60gfNHg/F+UIKgnFU3QRzRBnYJmHwMpoy2zm9kp
qsnfViWo2I/ks2U4AeP52cM7UHkcoICVcXjmOA6/l9RoWPiFZDg7xOz0upxvQycQ
USp4K/TzfQyTxk4HCNRU8NNHIdI+5fYa+Np6Mep3+poGXe3v/q/h3ImtRUO9XZnv
zaJ81hVDqtve9i3v0M0G67JdEcHoJsy2uDYAGMLelm3IyO+m0H65o016g9C1Ta4k
20ssPVbmVXHm/Qx/3EbuGlz48nhN0vGd1DfHu0Izy2+diMVr7zsj6zjh6ers3kMP
/FV38vdTJs/1qKsSMve4WsCjpVHROh66TZCBxNEtesm+7aUHtGiOwOsuyrVpkVsZ
SDPicSNZllMPU0cEyo7qZvdjbv68+E7Ff5U6MGURsBw/6mwxZAPAbgS7zt6wtu6t
u6X7Ijsvrrq8fIlZaBzMDQtC1rUy2MmUCrNc3cUzgiCZryy3NNddZl6HA1ump3Ln
kVY9LJt45IE+NfwgS5w/t8Ze9Q89WzCrC5nga0wV3EP903gyShJwgsCTN7kx094J
1yfLboXkXoRFEdTJa9+UtNCf+FnyK7tp2pu7KNc67GNamadJuXapKqUBkJCcNqtW
pmdrwFVYcn+mf3YN5629ip7XpSkXuCnvoXH0VMxea7AQ9vz9DJy+01/d3vVcjYzk
wp0/NerJNBeDRx0lnYWK0h7Qp1TmsDdFuBlm+jthT/65cu2YwXghY6aHHtxqSL8m
a2vx0FIJLriAyXEf1/YuSni5/uqj7fakYrxnHgnS2apWiK1Gou/6h/K0/4zzk4bU
v9fEGXqgFvb9rhGh8RmRI+UF6rwBELkFLyU7eZ0iL2C9HERb7ITGJ6vGmCAWJv+H
Zz/28Yk3iTLWcwbD4nESXcBB2x92eoLRC9Sw4UdSJRSkOgenzNujSgvRNu5gA78w
s7ki5jmmNspzXxqznyoZGAtIOWm3sHMjelHJoL3wXf35AR7Id6Ob5AolImzvOfzp
5/F0qfqAOx88yfk00eHuitV3dauIRmkPIeaRux26HybsXDy2+WgDJJ0bJzNAnt6n
gaCECMUEhfZjkCI2h4fWMtxU9aieg7bkp42w4q7zWrjFkIHmvjbruUG9rdddWSmM
6BrKZjwWQljS7Xh+VW2yJquME92lzjOP4ApDMKgxuMejIsXEuOAiCGLGoTCOZVpq
j9szrPmGkU7HwswtOkkQKCpQM0J2RYigmFXOVPqG6d9J6wU6TC3N8uPWMh09upq0
9Tlu8CUeK4NH+W8drno0YE5GSJ5nJRFAxjVG2t25KRB/B3BpOcucNiabtHJcFWfT
EuJjAAhJQN+mHE0kFcXl+Lx9j3ek+a2aFXCPlF3Yad0g5K9lb4/HXqCuPY/s/MI0
czBSQntHiecCUngvvD8vOSo7sV+bMnV9xBYUMugRwmXpzeezWQN58AGNrNvewu6y
nvTi6w8nyS0AtjdzDDpGrmk/Bx8Ts3NfbmErbA8ruwQSBsMBC4wU91j3oEfHidcS
wrN2pKVJrN7XOcM1n6VwkagASBTFqlGgypI7I2rorBcxBxvkkxJZDCiTZ54v7JyM
J7hHbhrYK9xMpnCCTmr37YIWL6h1i9fNcTddUKVBMb5WhzZPlD2/Wdde3H/CjjNX
7L4P7srqObXwB7+Ez9lMIo0aV/VNyQFsFnkp+8BaepNMCsnAGcbCCfwUUWeabxTw
+Yn2BnQnvPCMc9f/IY6hpf9abZGGAgkZz6OGCD68U+Fgg5AzuwxdIQgdsfRUPDC7
/AqDQfYRPumfQ65030xeUWdxAdcwZA2U+NEMOzM3yCY6GcH2P3oqdo9JCDWdhQdh
R5hkuKYrf6/TtxFDj8h7uCzs+1VHUL/PF2K48JvStp7SzgvIlcqjNnaZEQ2xq7tm
tPp36suRsMf6V81qgCQCiflP+KaqeK7P4jXWG0azXjB7vWNjMLAf19aZgROb2n0f
caSr/VkMEdgbF/JW2o1/qEyG3R6/eVSCSht06EcT/i7u4xCPhPVv37Ih0saG+sSh
GBjcp1MlNPI69b/jWKh3fvgT/EjXSeTNSWWChE1oWW4n0i7jTQ35Us/ITEH8j+My
mhFE4jnnnPxbOFyuTbzDFLvu+RU7MY1DqnJFb7rGrVsjzH4/2Agut6b2lY72h/jQ
l54d8f7dwtV8Gm20zgbmrgz2xBzyV96XxLdWz8YKV4VMv8Kd07pX+VlHjT9oCmzi
OoO5To2tXAg2QRh5Gxk6eAZv5GV15TaHUlU5sSCZIO8Hetm8Rke2dHlpt7xjwbEg
oLRVvJGuGAbP4VExvS+3gcizapWj2oVYBhAF7nTHomjg1o+lKD9SoD5iilhqvTgT
nb87gjgF966J4tGHpuedIZ5UPR8o1hlHGI/rUCdfplepuHBsc7KTmWrTHqaRYeqj
Iadrh44DFt187W8HMOQAmJcVTOZfNfCK3TqYUpl/ij+RFEHsvLwvhp4wO/lhXCTZ
RR6im92usVD+KF6AXTxRNpnJib+HE98dtnYbxA32If0EFAny04xp6xW0NiMy5vQS
YMv6Pc2/3a8/bSWBZR6ogHFASo3mT2QJk46x/RNL32QuJAoD0CZDnGZuyx1PRU0e
Mmiztf2k0fIMeq3H3yZkGUDZoOh+jnp6VUca4NkAerwujlDpAwK/YZLD1H81gRki
4RZ3jgQRISgg+yH+tUUotRxin+hFBlN4chIIn1tR6AStXcNqLj61TNs6UJQXqJ+2
3mRNTFmHy85aRzYps3L+zPYYfCM2ao0YOebdybqzNoq2e1GSjuYRFVVd/EQcBFrH
KMUhzNXWTykIEHxEUdynAhM3cpZwLmsuEp0N7GuJr8dwio5fweg8iVr4umYeNMnR
pZUAnv2bCF6jbfc7MeTV0i/xPLHIfNgf7sy/dAoA95JEiJZgVcAbtSjx5FAFvBhv
CULUlDncUee05FhxN9Ahzav8A368eEiOsxbPOKdvphWa9OlNBf3SgXEE3hAFHcwi
qNtTCT3frWP0ysOEThKkCAiCi12CbGKDpV45gZYu5lB932xreEbjLDv7zhpwiedf
nR9Db+NasD/1Adh7DPEdmMdomkTdfY/mVSmFjS2Kgt03CvKUAsjAyysaVDWslutw
AoHkYU/VVvpMxFf+2cdJ/NIuEw9qxnaqTLxGCUnmid7qDa2TGKG6pFOU4ypZIM9H
PcCDSJafWMMIK9rAK4TZR3FDK0D1s9xPynqflngwLpKkXAdZDlgA37wgAJlPsn0a
miKNy1yYGWc+0vj0Q0rITU77RtyMaBSmfV9Fu2+30t+8zND+E47Wh/RVyXyauoch
r2Eqte5aTAReoEYHcgQUBNWj0bGKG7RgFCTGAJv/jLzrceSk/ATXF2gzaTc2sLRQ
JXQ1RPXcSauV1iasZFWpvLIlNlkYzm6cpDpGqDoT0h+vyJdMjgLz+n+VK6nYv1NR
M+P8tKsl5JcQzYpY1zUAyROAJxJ+KbSPdHtpCY9Abkl9la56GFMi+HzxBIChqa6h
wrtSeqQSw+vgUXEznP2LoZFMe5TlXBfjybxUSz/x5FgWzU0RQQkfdnl/iV5Eme/B
+7vteLHLp3DVAU6I6AXHkMtsPHqKQJe7Gi2dXYq6pvO9kg7MLzD0Vb/ahN1VfC8j
sf5bkpTCYaKVLSYfE+HIACz7rxDZnPZu1ePB7XMrD4bMYFZ/N6IezHySHAEduuII
KrfWEWt3QyMZlAkbjirvxJDvkcc6UNohAe33EwLuq+eUfuB2CKLTSdgU7VXPM2BW
C35rn4MKWRF40whu4Hy7de3GzYuhSZA6+VlABgcfJMvu/Pvbz2KK/adWkckNQrbL
zIxDERolK8pqJ858UGVi5HV+24QWu1aqOXbkVZKDuttiT5QSIIM2HRf9wf1s84T2
WSwz9UP+kMXrzn+H1tZuvptap6rFgtMUALTSKT0+/Z++rLdf+rAdf6qbPIYXpK+Z
hMBHcS4/t2h9lkDIN58HfCO7j3AjPfJ2sEzuDbx8kt2b5zD7Cr1GPCfDZNERoIl/
+gqQcMPneXw53JB3ta6zana44njCTaFkMnVM341oaPwSWdCSI6n/J261DBZ3+Hxc
37z9HLyuDHNf4Spa327H5pF6HNlrUARJbtL7MMDD39ZaB4q4/twLAGkVobJOk2UD
Kvg/HCA8aNMZeX3/scs7PfGTRyTtDPSvVXvgd0TP3QOHH49rH1QH6mspp3C4jUF5
qFVVpKaduMTHxOAcOqO3gNgeDAKGn9zR4Oft5yqUitwxVZK0cEfzH4sCdGGMxsN3
97IGm54rK/6Hb80bz/CbchPCQsBP8suUUhpTyE9ae/w5rI1750YZEyKShl5lC5Su
OGtDQqp8judjK6XTCQNBz89MSyaqueF0lV1oMOziU14148bMa+oDVHBa9PKd/4IA
k0k5hno4R7MItQvpk7dV+h1NUcIU06/2+pbiT8+p8WHKOEOsyMyWlzv+7+qEJniy
G9R+8+VADpNfC62FM2uUDwDyGPZeNB670eNVjT55kTUAidAHFrD4M/jgf89Z9z/u
tkH5MXxpw8fHJopvZyE8OJ3M3O7XFokVY7JmKVcISy3uIVz10xKzhh6W4B/Rxwxf
99rilFZ9AS9bMHG+k6D8SqQsIDxDm4j3UwX3/MDS8PfLye0iC6+ciEZuYx38D1DI
rAbf+jEoxcrmSiFFe45SCRFOFh0lKnbklIlX68WZi5CIa6+HBrv/hxUvF35Dmwjw
MG1H9bCwjZHCLMmPaG++Rq3erSJL5q05dYCgCCzTjIjBD65zBbKG9cuH7bIKRwg6
OMOG7bPola+L2YHOWn8aZBfUdqdCdJk3R+5XNTvynGbuS4x3nPkynhyiSFAT+OcJ
XT/IJqg3i1FV/WRSPd+SgSs1O5IiODQv+Nr0sKHVDSrm8AZTkK1ALo4dOUT9im5m
06IJmeIfdFNSPg5DmWS6e3+JCsJIZuawgrkKmmiQ39hKPqo4bj3uebAfk0PtZYm8
hq5J2Vv9xmtam0540ZuujqycsGAge+tvQniplsSFSGJEJLYjJ8caKcghgvKMKS4X
ohHg5ybp7tDXX2pYbYi7+StanP1WXvzol81tK1w9/wshEkmpkgaxlcoM+fC3ysNK
gmJPBNqgOmYjWXUG0/BZTxMtUi7YxeZIiRZ0uK30Zpt6qAYrVZ56ctbM8sCetcSo
HbuYgxKOUUkdUtDGcSwuts0ZgBsDunVvMSzOHnHalLG3AuIVO3L8x8rdbWB6qRoN
DQO/HjjXVT2IF18bFHY4suewueyxckv2umQzGnZIPnDzxojD1JWd+MlBtW/32Pkv
r9paxuVAZHYdKh3MQvuyu17mbt1JxV/kFFJ6+IGYRzdW3+4LaRodGBsUDdHTEeTx
aHVYX4FByMaNdu58ZQORGaBTLlv2Vt5qNoQcIFubZRPzJ4snD8a3c3B5WskHFyec
GWRh24h8LMoDyH2NyWOcVxS1/Qq8kQmD34wKC9+jkXuhXbenvteTOrJXr+KJZgjU
kFATqrostG9zUfZ3dG3Fk0IzcKSjs7uHXX64ujT2nJv8QVaLvvfpbRYXRyjiqz09
8QFh5F/m5FwW3yezn2w83gkpABr1NeSKZa6GyQx8LUMC8Euh3YYrfZhxNCEHbXeq
1tXi7Hg4qx8Qau68ev1Ano3LHlLnV0aY/zumCsSzoq1H0P4ZVtN1e/mQ5FdxZG2R
JSDfiyuwAj1ejvcDTN4VTQXXPRX1QgJrwLlOBMgxLrL7CvHHKAQN+nzvKyJRRO4b
7rHJeP3wKsdP+RF0Y2jTlAmyBoXJz2fAlojEut61M2/oDgFZQ1RUMs4ewMlrHVcc
lEO0nWwUUmdoKyNLz8m+zUuHXmhKGZ/WUu4qno0uidKMaw6RfB2CfwWYErg3Z0TS
xeTtpw93Iq1R0pRTIVSu87alXruWuueKesrSquuzx+mmgfIaIqPySk6wgX56lebx
b6AS84cqBn+zBSWujWshGugHsHG0uOlekLsdn4AS93OJ4SZNlDK4Q2KniVtAsb0O
kLfpVc43Mi+M1Ey8IVNj4tniogUlmxYw0/+VzA2NUBPyz+04Wsg3JSERi3NL5uq1
vmlMkDR1aP8PjIu6qX2GKgdVqlpwHPjaGn+nOxzHMq739ld6KfHz4KSFlDfjjO53
smDGORp86DEG8LRnp69m49ECb9Mg1KXLl5Ihkg+fhGGIE8cwzh2Bd2qNLLGUUXL2
NrCKtWyLZntc3tvivFLXJO1naOZRGNOTYYrCC+i7EZwZnyToxabUBKvP868Aif6c
qHBJ626mjepvPcXttYStq2LpP7evVZv8uEQCth1/7goeXvKr4StrOij+ORef2E0i
AOqRQ8PFlA9LVBRD/8ZoDVb0/Qlw8JIX227wbrqErd/msEi2p5eI3aKqPGLdSN1h
u/a9TN9JxCa/Vuy6JmMojMlJ54AiLTVB2mkFdtZUKKfArQuTrRWtZTkHbSJm1gGn
ZbbGFX497p+zvR0xjCGEsLWiCIiMwvWVmQ/HrONghKlJOOSlxue4dJdrT9UmoH78
WQdUbL24z9hUohV2H1UNG+qNq6phH9gM+PxIoAAZdT82bkIXBNAFzUg52A4zPQjg
Ko7e9vHmOb9v73FSA+D5PQD0FouLIC2FdM2IDx7M0LzOaF4bkg+4leddFSNbQmX6
dF9sbeF/R+avbazq09OGdOvg992jp+7/t8nmEHpzab3cw1FDLMcypIyZkOWWFO2z
TKrz7ZnWgI3A9phnvFZfYGZECbmGBp9BecYp30plk6Q5hti4k3zDnCGe4Ovyuvof
NUvxlT9ziJZ2Vuc7qSCsMZIMDPqJWv0G8eGoFWZmCGmLMAq+VEmLqY2SWqAQ1NXs
B81xAYNX+ABmAK0eQ9EYH7cAHd1E9ICeCAP/4p8y5Y8dSFimjr+NYiH8+hsybgH2
X2zyrKPe6c1ynEAmzcHmZd1K91hWGpoMtG9+x7sBcLXtrWS4ObAdDO5bGBHk4bIz
Ppw1WckFqvf655Xm0ThxAeT801ycR0OaO4TfNbi4fXEfWs3vRMqj3S8zH1etz4zy
MyWaRL5lvA8RCXk0xRD80aniw2O1mfcn1ikjfpR9sAFhYzkuW8U6KOXzoV/gnZSz
8czyRk5omW9cBH4bxoMU6pKi9gmtooCwH8Ner7cl5BWmKALCxNO/aneQ9oHjBAzS
+yWujHANElh7xnOQVmhJcADFpo4warvS3QScKC5eX/IyrPCOJFKDkZx6Y9DkMPXX
4MHSfjHdqR5S9WAtYZtt0mO44DQysRdt4l86zy8XkAeGFWDBsv1qeBXJdjVVeEiH
7tzg89QpW6xDRtxxIBjV5oChB6h2BR9A+P2OdL0NHVxC4mOCTo8YLR8JtB3SXvh7
98YOIJeSPL0sm03D+q+3xIE54PimhvAerOy6mri8ozNugLSa2Z1MyD6ArZ8PwOU0
wl0o7mFZv8JiNn7egqi6nHuV0cTpmVvcMxGdYOCPK1YnSO+5HiWabwZ8S9rTTFQf
bwLmoY8fQPA5A8ifmH/nCFWemt0qXUET08Cmb+qIA3N5HnlwZS5WWQ5JBc+DixwD
aMaTI/ndSiKJhIn4Dz5d5RTnWItJWcJuQsC3gTgOvcGmOPjQVEzL0uxfHy3NaiSU
xKIbMTl7VQEFoCKksL+toe2WhsRcF9JDLCALMfg8nfKjIKNYBL3e1r4cAderVfSI
Kn8Swkk5m65KnFezFU75HTV8RtqrFplpCOuN+leKoGDbddnZZTl53RJ6FzK992dz
QUp7u/u/5YlLRVtIcUd+IuCyM0IU5+t7nDxBBF6MULZjWiX19E0yfWjKUMNy+q7B
xaGyOgsMuOTRJUTybRUQFagCQ7Ha0ck9ocN/zDIJdfH4DVnj7D2obgaWfzDSXKCD
Gj4hZtZKhUly0st2q9uOlUEetDxefd5yqqf2/k1EsXFkPOqffmHk88NyKThO6oXC
SX5myPXIQqXNLctHQ41oXcDJgwLYbyLgnWjkhVcF6d70EB6KKEUyBhjxOmKg7V73
lMBotkbtBa+C7kPLQQUPdFPAYMNoLRxAWrbqHmAmEALOVI5jiDJhhWCdI/NeRTkJ
4HRujvxY+SFYsgR4P9jTSCBoB+tigBfzM4aiag2+uOqZK4M6xQs37D9/UGdwQF4J
lp6NRdNeQQK03Rif8GCpDUr2TxDvhsDyolUOHR4RpMdZw1SNhFQiXGtw66bkB9X+
OfPP9QclNzG2eSGwLiCe0eEdYJQGMlVz4PhtgI0arzPYidkuBkJHVzt8f21X2Z0z
ois5htZa+uUewrGuY4Ppt+1PkNVnXV72hqBIpyi72widxZeSlQN2afOktnGZZiRT
f8v4v8pUHT/BN7PyrMHd96er/ELvTd/sS3mEZ1mjfMGfOByvtC2p2eatlYdwjlXT
IOmjIIyqai/B8bJLFfKDce9q2NSr3TjpMZsr1MfyKwcPFCQeHGNxrdAYsBuyj6z9
OBjgPjovNqKsLscMrbVCgzAJYUFskbMfkunmFGd3S2yY757zXD0fTYWwGma5wd1u
iLEpZbYGY9/kTv5rSopft2stDghj9Y4/lbMsuXo2w8+BjDGPVBgwoIA7cGIA1PG+
58CVRtP3zjaTdvCje0UD/j4T5REXpWuO5QY1XRP5KUYQSqC04jxlGVWQd3w2X0l3
b8OCcXd8lCSd0JeVxsNGdLi0e0BWkyzIo6yLXHknfYPbvvMEIyPhtZ49hEEeCYzr
QL+wBxockC8ezTtInpf5XgQtWOO3IWWOXs3CP/B7NjS7wJqt14Nfa5dJYppDPK11
EPoVi4ATl90RFANZjPwuZxF1jpAbu2W3ooBLGSwTmQFUfiPj2EmfPVWk/beHfTFN
0e+0zz9HJoNYWX5swzSUTFt0XRHCXDKVEvg5CdGWnZM97x9m+jKw7btOQ3dOpSDf
Om5GAmAde4bhX8DYVtGaPZ2w5Yfaze38JxBqX24LwB4KxXY2TtI+Xn8WIlLvj6MY
BUbq/5jhfboYGyEFy7BROI99dYN7SeJstA+ueJaw2m2aHJv+df8tvjnsmt2Zgcz8
IWByArDZNEfPoxUlPlvwjuCSpq77rQMUPTVh3jVScUUeqKjv4DajksE6OCTHCli0
OAerGvOtMJ6KQhtXrSBiBZgVbPA60CraKWtpTSszdujRDWeSOnmwmrPTIDfagt/C
CTLPVAjwqbYHSsGOvxq0L8Ca7uPclpMf4dxp3ZWrA2WmyqL4bKRRkY6eDeGcf1an
Rc6peibvu78blB2N2+I83/eXrv5qnb3qGTgRCzCgA2MkMfnkEiIjesaa8q+/oKW8
aJV6BTotTHKn800rp0Z+ZfZBz+LIqEQ/9eKE9JWJTN0hW1SOX01VPVxdtqHjwa7p
xB6iDDehLzMv0vbgEa23lHIG8AljY6ujX1DaxYh3mpahNbjkdow6tIw7YgWjmmhu
FfVp0GcAz5kCcFVlUFKhdcxOfjj9YE/R41epcMt777IbvkNYTtOM5FfayYvnfqd8
m6na47Y9lUcZw4pg2nBlP+I183U1MyNbFni3n86p+mEr0AY54QFhB+NF2t97oimy
zuzpmVV+WF0bxGhvSBdIeqNwk4Rs7v1IDEDnuy+XWny/qKbWIM7YTdLjdwk9tNhx
t01EHKXi8T9l/NVH9mv8ZNrV9hj7K6y6lAr/7U6CbY20ZFFmNfvXxFXX3aupTWlp
adXrBkZHduO6A+7wHkvBNCkqqZ0IsSUa8xO23Hdfu+iyufFoBzays0psjEzt+ms8
jRrXqvhoDAzb8McIc05J0w1pU6GGonSdlaSLcH/CzS4oiR9R9841bCA9m/rLp6T/
q9+7h/UnuM4s0Wd9qsfvl4iOPsggf8cTcYnL7UEDPu9f7gsHIHd38QVcab6w5Luz
ULeXd3WK/LB4YZRpQBOFJXnpp+HmzCZlo/QaVJQOZ59Mw/Ma3VL2wdxW6PzTBAP5
Lo9Kdl1QK/vWyR0CffAUutWWBRag96CWboxZ+6aNcqVsKJaBl3yjWkoTANPjpUeV
DJ1xbYnskRjKXG3Wy062iUU41C4vgpmrtXwCNiJV0+MfO9q9lKUFu91pKs1pUbqW
G+FbsGB86GTQEz75xB0hCJSjkzX+ep4LTgwPEH0Yq4+9WDQLNKBJPB7bofFzNlQi
JP1XrKIdONeAtRQheJi73hgRZwSiApevAC02CcdAcjjyoSHTCJrHBY9RcrC2+40s
q3LB3RxyHxyWgFdQGwq7LDusWr9NMXEAFCCEI5bRM1XFhKKCl9Yr/c7oPhGp0CZq
xDFzdCypg+tz/LlzrfoGfpMSYOvq2ey6EUeDOmDbsWejgl2lTDeZaxkGWTrfiJ/d
lVjPyxz17fcJ+HQKJQxiN79vMlKcpk4LL63Fzhm1vQv3a70JSt/Q5RKePOTR+7Eh
+lOMskXgErI3TyiqUL+TTqddrJquRXgS48SCBSfEf5lNuDVKD5S3d7uDGkRFhdZP
8WrU3IYoLHYNsF2V9nEN4SQhdQdk8KIoCaLYW6Wv0zEAV7287d1wWn2lvJk9200P
oNxfOcHXtKLPLzGgsM6+d6aGQfci0zBd1amB5gUhLLFK2PpG+j0lozYCqOHg7iqE
ryPUMlJY4q5HM3GxuD9LQkqa3mHBxd3dLONJc4b7oJddHfh3uvH7sveomdaMp+sT
Vw2mZpz7N2bm4rMDE8P773t6PfRbnPte64w7QOS4FLYQRN08cH5WtzaVR5ibBAaw
QYl0xHL6GzhCtzNav7FCeubGGL2znPMWXJy2guDCPpfBATLpIxTaAg0Y3K5RAakd
2i1VS+qxfRPzBxy0lZkeEujvR4njMTXjd4zEZao+V4N3R3Y/u26Xy6y1IXtCg0Rf
ERezOwQOzWUCOQlyrfNrRoDSCk103knszM8QBjhEp+6kwh/6+igzJSGp5lwP1jzH
6h3FxJhOJ466yEwG1bREJxQx1C/DrS70D8lfEYNl2VIY7RFqAJu2oyLFmA5Bsbh7
hTnrZLhwXkxLwTEaO2vDEhLuv3hFwA0eiz8jdGQtwCffeounAN32DZ+LzBqQfyhp
Mv10yoP7Q4+/lXVO24q8c5yT6jrWzoVkQnukfSQtaVdW3kuQ2YOPaE0cm9BQE1j9
QrVreluZUoAuNUJuGfojONSYJtsHS0jPG0Xg1A0NMV6OhmhkRlVChMksYSkJBxwu
NBr1KGexah5NKhCnBAN1TLHishRs0rK+09LFOuHGgnh3T2scflCo1JeuKg9J13b3
fdfkpbpQNl+EuSKTr3Y5IfnAgxmSxlMJu+4EwBUZjzC3UApo9uhtn+arTXu2U/Os
qzY9hhrOqlxhaGHkXmjn2gpJaEn2MMOTmbpA+ftZJs4caTeIaFR4+MS3Syep2nkj
t0d2rRWfa7xUHmrWBYAkeol0g+Qh0/ec+RlkOQTyRHmAgEMXDpeRbV/gkyHcI3pF
glvsXD4kUB+XUU0AV6pBdeNsTuomgkly4Fv/bg2Mp1YdthEyi95PWJqRxToPlyMe
IcdlFsxo4vVvx+iF48qv9ZXOx5ndQKRKZymrkGZ9opxLflMnN24VvsW+vD6HDmKp
/dlOkiqTcQbyVXV1HAtrorbPtz6GzC1IH0BFnczPlpWLslU1GyXxnnb5AM/Ao7Q/
bPBPUAyA4sn1/RNMNdFVTO0V7a65Dqy7+YYmcu2/UOp8dz7QpE3yxkfOGef9EEKn
bXyg7ZafbX9yZVTz2gcHlH5WlJmhhF3A643Rew6pLxtA7pr8112Pm4Xet9gZ+Y2W
XNxNyu5RZeQfXmpK5EEnM1r6K8SjEk1bZb02pRW0ayF4hqGXO+3dcNTf6H1ON1DX
ofcS2Sf1u99sM7bck/kaos/iI11eqbg42QYXTi4YRlQ0EHpilnBYkWjVqL0Yj8m3
iFuJVcb0n4CkYPFou8YbF99rVwKel8lnh6eBYP2/FiR9RqEIkqEFmrmCmiXCI1fD
AkEnxfRyCY3oQZiAm6DfZ7B5elCh4D/EUb4TCPYfgZrvyJCaOw2+ym0iL6awT40R
dts3Y8WB+1f7hVd9/QryvGUsdggNdUduFR74WBEidCrEURFxs6crCT5sm4NiSOxf
BjSunUYVSqDGip5SudCylbG/QuQOamVfrRNtq73Z7dZWXPUxy3rvk9F5o9F1tCAq
oj1W9/xAmFyIJNN/h/1Ne2oKnBJOvzfZqaq5G8hcUbUIIKAxuotCdmofRNS+84ng
stnikeBGQesfjlk7kOam7WOlil7vq1vIKSjUy4joBory1GP2Bzzey2iv97CINrTf
cz3zGNgoZGyL1TUMmUYPr0flYUHqfs9qlct1Wd80jl4UYAKFAFWBeMYiA3BpNhnc
xdPCaSQiWZ1kVHwYS/nRGMfzXJgOCpTwZyG0JP3KGm9y8fTPin/ivOIwOYUvieLr
h9HhQYrIQ5BRGrcOvq1mZykfGSshgq6f0KlRnSFlp9wPOaRb2VDzWdC9T1M4H0FV
TFDoymGLJEofO2cNiZT9YBfr1L4ym7sKU77ODRIuC7Sox4K+EheS0ccTALSzo1Du
Jd/YsZbuyT/zEAPT9bBalO1IPDKjtry2IOKGB/BN83Ex9OmtKTS7nxVvdtAGXFlO
GRhmjdxeqq9VSoq84zeGTTtEhG3VesNkWofQXALqRvqr+tBoAgu7KQcWobppIbti
b01skcuBl8HLl8yVSjMNfQTidmOgJI/C9/8EFjNbR69WqzzGJThIT3TRYKfiljr4
VkVktdVbfzWAKlIL3xZlVe3z3elMdROW7a8vGCIoBvQvPw0fEHT6cXzAivFbcoh6
UjuHpivJHfdwQeGSLshcW053BJvvtMnVJmMsBz+04dlWUmn6iVZ6iWAmxdvyO/tZ
0yOwhnLKKJNRhSCvTLv9tkQvuPP7EHKbEz+9pF+gb3AHYm5CWX2FYTqi/WqIuaAP
4TBErHJykWHzH5qRLlEHzUVfQipSiMTqMg1LGycIdrA1P7Zoj4NsV2gChY7vyGvx
H/8t8H0Gnn3kR0nVlu/scIl39YnCFe13WH/SK7d+VgGYs45NjAH6ztMO3aQblYfc
Z9OJZcdVN3NaXiQxKda7eEZpgYJvZ1YrPpWe+avegHZvilissFyRZVypJ6/s6Wer
TcNIDi/sjji8NLevg7krWQrB9CTj0kUYv+MTQdfLd1Sj6SpxF61NwvDe+CDXiOMj
K0tbllEFP9Wtxs1roYObiC7gOL0H+DE+/nygAgbcIFouzBYy+/E6l1v7rOtoI8zS
QtoNxIx/tBuQ5bOwq0YKnWcmQayMoIdgz1QS7ZJkx2hiDkKqoCx8nJ6uELWl4whF
tdqATs1kInFRpjl9GnElzX8W08TbN7Lg3hXaOXOtgBzKWmFF2dxzwo5JAe9CEy+y
Dikhg0WLBIjh67+sgvXziR2XB/uEMFLiNP0VAujiY/QEUS8Xi9gd8Y2LVS0FEh6l
kTzTYNe+EI/s+UmfAKWxWv8LpjApIDq0EvzOgOHJnrfiTmRE15Hn+4ecDeIg/Iey
zNL/qnpJhDz2QnQ4V4KR2rHv+bWSXG71VEjNYu1jpTKijvSIfcYwgXhV2RoviWr4
3IuZj/Wh9trWxhk8zKxfv3jnC4PV6A2V3SJv3BTSN8/XrLTqDtHKd+JUfjuO1xmV
FUUoOffgy3iWQ0e5md5EeEDAuzyLGmbwnA+Vg6Y2LeQ6sz8hoig/HYsRIy84fvpA
acQJ9xi00JduEtr4Z2OBTwgj5SX1XGzJxbHUAKtfboIe1dYp5h8QC6MQmdlJ2vVd
5ZANRGWDQjJ/FfDDYPdm5Zqb58AOTPI+mNMAUT5fc52miqe+NBWZ/cjIPYA7jdw/
S9MyrSoKLQnbu4IB3r0b4ArckVEesm4BF/RkU7r0o96ZB59pSwL3puwoaw18C5Ar
3ODFQL+VJWIxCqS32YWpbTb/kge9pj7A/xQfTK6hIgTHlNTGOaH4PHtmqmkMWsnl
SI0EZ7J5NNQ1kXo7Vlmc0yV18nZZbf8h61hvdxXzofGKLHZCVDtpiP3Kn3vEh8tu
OD9kTKMzsl2m/k7RodvE2XeTBlL3LTWJEp/CrswMIIaRmWjCyg/E9lLTMelVI07l
hIEE1q7APMLeQHi4a8odr/vAsjaNeC+2jwAVBKcyRQZX2d3zEd/N0As5xsdvkIgg
wTk0Di0tu+HL6QUmHAB3AHATWT+LxLvRqFVYy/ifmuIYpNCPUROeeDne4O/o0R8u
t1u+K2vpf8st3hpODEKm+pr3iUTC05qBcuAHWa3sfHM7/jUfNuvdN1MotEcvEEhA
tnh068xDbHuNvT8B2VmcD16tPCwJmXG13IIYyAbCRElkkE/1YCYc2RCVJPzoxcks
pknvtrkVCTClOz7rdSWwc+8wPwG/ovooFJ0ROusGV69Bypez0TZMhTVtZtDboZOF
b2lEEpSFuJq38KjY+vWbyjwUUkhrKDGFToocdQg9iQM0n5ObqUNHbWyRsyOsYrX4
youGczLeWLXPXKEEhi7g7nPbjCTEWaGUjbfz/EV9+CdcOZT9bH+RKKlUZIyb7uWe
eY01YBeEwVJNOwXbjHXQSjObe7/nR43xXTJLhSTQOknTCjEbdF39tu2WviAPv3mM
+cnOxlpGiB2WqX0TCNugYCMd25RnghvxMxhPney9ndrkIOZdFZCNOT/aN91jd6UH
mZNZs4vNPr2r/Bf3lRVhPHWGlyM4/aAPx7y1oEOu0s7vn++ufAW7WyaVraVdDa6N
SJx3flsL3NWk4Sq/RAJKnIjreHIz8XeWbqr/SAvE26t1FA/WV0Dl62I76/osaeNP
BEXa8zDr6m4GDOzNtlZZJUAss9pz6tG+yEOgyR5oHWaipIvKnuhdUBQ9OhPvZMsA
I212p25CZez3TGrexeBfeEO+orSfj6tSrPsKcJwLyWjXoeKEs50FE76/r0r9vp0t
Li3KzDU+mv5aJnewqWuegolfwbX2hHt5dzR6RDo7IquoywX9VNfEkzgLHzhYWVfx
DLFpAWJsT6AMVPoWdfykfqITAR4WqHMZsu/cxQpHBqyfOloxqWalBwXs5LY0DNiu
XlS7UwWpvj0AcB0xVCTVInLbmNuA2ljWjFbt44WRBXl/LPEt9jWGLsEC+YdMVkJ8
qhdZUiAk4u+d1FSil9WIDajojSF0IJqoq6xfZR+tdfIRnByLmscTzOaewN3WeeCj
GthJOoP134+CqjCyo/VEZPmdxSlU2PCd73Dx6l632yDuPZdjhFBmbVi/JpRnk0A7
5n7AD37KwsRZWoA/6v3o2qTmUWRG8l13UDFgZ0uzXfDijivV1ktrU3f58Rd0xf98
tqDRU2iYleDs4PCYaCKXKf1GL9hBCt/FiY04Pr4QCeaajqXRDx3G5uyKD7uw6qGi
jMiDNxJmhx14A4G4WBAR+ecojtcXp4U7E3HT6SW+BZacizHQyCFvw9J+5BtNqzua
OULAMYKUJu8uk9+NEkZm+LNWweNwn5S/4x0/z3vhRrB6p2DYUtwDyG1SdDhNvMEF
uKnf0X725pIDKx5/oxSkMNvsCFWzghaZiYoDt2Zk5fgnk2B7BP460eUyekriab1S
pz7Q+EbLYWGvi1k34hn/5RTKj7tmve5j+uw7L+cK5NEzAasamnse512s/gTBfu2A
uTT/0LMeX7plIq3XGMVR1PT2na5zbpRDYvXByPiWv0+4qwI0a05hXSwx0arZ16V3
x6YxeKgMJSNbFNZG87I/X3QKKv/iYTzHDpmr557kHX0iXm6gEPZfcb4C9nSRvT7N
wFHSbDjWdzhHBo62rRnk29F2SUMFnUsBGQDsNsiEcvtBLE5LrBNRuzUlwXqTlaht
J89JRMrsMbYII2h/oFAB6iiTelvTI5dLSfYGBm5T+lgfij5hyrAR0H6FNdtaLpOH
6qqoZCoI+3E1ziFf+vm/FQc1GR5U2xMK1JfZdDhEnmBHtBl5tksHGwjCQHn9b6yn
n8J/wVSBQenTpO9jb1qzQjmYHwQyzAwIMNuYiv54kwqtNXW6wSCR/KUT7uDC+Zzz
WjaXw5ULgUrznJumgfqGJWozYgZ/AjFBcoBuNUG0MhJJvaBkkq/YHWll3RyDQanv
kKH8oXxPEtSktoYE8BZ127u3S8hbCySKzkuhR75NB8/jfYw2qQhSc7zRHhKHb6Ev
NjHWQzGsT4pkiwmuAimQdJ0QZOKB5ssrLUuwWSfIwafdGEVrMT0pWhBq+F17nGbO
PIKQxb/kij1fRgopHQpuIU3KkGdtY2gBnlyBSq7WXIej4svpTpxQ590Kj3TzxLzT
zKGwWEwtAF0XEXXOz6LtyB5BJ3eFRHfkpNQmdQOPlBzEQSMCTAPZgZElPizlP4yV
/T7F8sZFmaYTikfIOZo2Q72qvD2hrAIptmDjQPSIzwb3kA2D7HW4AuyStF3ZkTrF
3RmummdGVC9EPBnGf/yIDV5vINV9yBxqJqHGC5f7KezuJNXht42IndWCon5AQpsO
2kuAqea3lAYSeBS+YONphsHPhVl9cZA4Jxb0/5mMDpq4gvrubD7euPFl+3wHkbCp
ZAjREf7mc0p2ezx0+loxzip1HKGJzEc1MO74hpOUnBYNwlxB7AjTbbgB5K4xdnq0
KXdtJXiw2yQs2AOSMIt1cmcg7PhB190tH8Ol1Whuj+Z05pmsMcNfXcwmunEEX8MU
n/McLN6a5GMirPpNjARImNiK9OpseQyS3uwJ16fT4mtp0Ys2OdQkxMn4X2waJ8E5
GgIoYPIkt/OiCYHMA+0nYk6FEvYLlzOv/uEFLH8G0PK82167A8/0dI2NmdeOKusY
d5QKQZqeTUE5/IaynahS0m4wBrQdaDb1H+MJpUrxGn374LjjwEcLiWjnpr0gzoZi
QZUbdRVosJucMKz6WY/AS2famaHv5WpBt9JYkh1E3IeMUVtDFSCm0jYs8ZvHXgJS
zi5lIQaWiTZKbBWyZJC4HzmYMv9ZL2L6qgkEEk4aW9umbYjMKms9nL40aLlBLsXp
R9et+xQXcsww4jvPWz/ckqh8tHDDMY7OiwUVXmDUQTWJYBGqAZwFEYKaOoJhyUJI
aetjV8orB5KdXRnvrMkcxOgcs9MrMw+GTdwRZSoWkOD8pnvNS4rrlmrRKhy5PkNi
LKFkRnjXU51GKtIVpWZdLNsN0CNKazUgxk3k7Gx8VRXjfn2RoOJSe49erYSs5Asl
5Es7fZbtsiBoIexcr6+eXxbptGo1Ent9jEbK6QQHipeqnigH7wBScma0xguw8o2m
fvJZFaKQtFD6mjkv0qOKjJuOa6Pj4dfnJtWuDCVLu/jQ4/XQRPPFy51UAMG7igp7
lrJac2yePUDaYJCWcwWoxLzwe3hBva/Guxai7nMshfK7QWGFg7DAPkrJaac7BXG7
2xdEyc6wTWnwAxyEAynKcCfWQAypvkpLSxnQiJt5RP/7nUdoOh+HtC5Hti7Jbm5l
UDO6/3jJYZ3946BNRFbwRJp8HXCKmeLfYXaUrL4rRq848MrFkeA7KkFgaP/mrAgR
TV6zCE0JO/kEJW6Bq9V7msXYPsKhb1+++vsL6R4J19HMsdIrpeVvxisxMzEyM0fw
EkGGtmuyPPQ/fwBP/86cMg/7C2eygACyVva9IVu5iGMQLstiCjgJEZ+Ah6RvL2rP
Hwm438JFq8z8GjXVkc3zapF2XyDqbZ9uWvMIQx5oOGVQc8N1IyZI2Gr+BaK5jCvF
SA3bbSwSS/XWpXJtNlcEN1CCMMXtvKeUvp3BTESJWstt9f8e0suE8dmT7eYmzZGx
tl53hS2X8S+FhuYu+WO8VCSKvGewshaiA2HyV2pe1/CMvabL21eeIbJ8aKp71ltq
ghhPUGNbnO67TwXAh6bIT2nb4vjew8N+MPODWlMsq9HPcPuc0OvAXMlD2Qrbwhsz
nRRthufYwpy1hwEqnmBu8kn9iSk/z2XLi8dWEjtGIHPUOibFIzH4w5j9Oq+Wf6A/
+Mx8xymcsCKyhO3HfYnVnmStCCXjRcmTC4Ekev5l+G+7ajoDguF7ZEJcQ+X0LD9D
4ihzdtdkfqLPmNRDFQy6+QqXHva2Om8/ndm7w0Y7T8+RU5xG75ADWZ1lig/8TGyG
H/FRdA4OkgnEneVjXXPcfQw2kgtAq/HCGnmUpWNizKuYLJkvZ6xgCrFkM7SJRptg
kCIiPT+dqool17uFmZiml4d7+Aa1OrXVz7yDB5QfsWGW/emcK5FMhndx31pS/wP2
KDn79SHDHvnPOdTphKzl2pQvjSUBEPgUk471xanJvOHlD0PvJuU8U+rc+SBlP2lt
6xUaC+6FFrptehHQKfuVup4KUCxFNebb/b5Rls5eeWg+dUtBPy40nfYhcjtjCYrL
L//Q38+zRmZwUld+63I8Lm49ZgG5NxV5vBblEOpIqPoVVPCN7NAXl928vvbQbkjY
/cJqK+NgLvejNt0rtKDdRX926ULH4O+1VCg6K9M3aqYH4yBXQRFwVvkR/lr+hTxS
yJfaPt8WO9NE851AflmQal3ZyDSlDq3mhspxpHAdO1TIk/0zes+8RIuBJqz/2joM
exm8FZFAmpLkJ1j8rJY68Knuoi83C8L4IweZp1zeB3sL+nFDmAutTW8eTnlnDpSw
w/EIBNy0X0ufaCUI2SPLk1xgIoLYyfuC1feZEwFy5JG8Y6SNcKFMKPdXz6SBJt1P
vl3KXjnxIOaQsyxHgqYM1g6iSXSd6HKZ9QMxY4CTm2Jzy68pU4jr9NPuAi3bhNzb
OqUYMyv+S2du8x3mkOCWeyGZW9Rfq6N0AP4nyELVeFQiAM0pX0JoHZbcSsryu11j
wZ0T5sYQxeXLp8RRkhwS8+5uAw4pfNl5OKEJvDwptMuDfuB1S2Q7RpBM2MgtTsSs
gcQDKew4eV+WaxU4s10btDtwBvM0jrPnEuvhsotWgXbo/67AZJ8jXWhEmxuNWnfM
Z0eLhiz+0HcNmCxM7VItRVg5zgatgZeyGEyx2vyz0oWc/H67L9oRC81/jWwagUK6
CYJkzUDzpq/5rFANNWoyQWZqfBVR3bXyGu0U0/L8xFDI1TmCQF942UQC7djDDLDW
r+MwLb78Q3azvkz+GkraLJIhbvIntoSv7gV+VZqJVe2s0VKdfRt2i4s4BSyWkyP2
Po07qVSQTEFeHKrBtZ7O7HcI9eNiDDG7+MJdhrSvkG0EIVjPbQ7rr5YF3DIiHu4e
zAl4s22Ea3iXb0fLLm2fRC7o2NOo2p9wLGAN4r6rr2+g+q3JPHQCdk4Gos8FNybh
OJwBtTn22PamdOueodFxZj19mNrPzuZhWkNhSiyKez3vkBPfWpzD36dAV8WY+QYw
o+y+DHLjQMIQHhhZR++Q5X2fzD7zU6IN8R+EVv6YTgMXxj58mpVo76VF+IG9Xfmr
lHure7bl2Yz5dZHlttxisrUJGjmo+ZhxFakDyqH+ug/Oqeo3IR0JOTXfVpPGkWYZ
8xsNI9AsGc9VU24HpwDYz/LD0rLlEy2AG+dZ5c2sXVyTE66DnY3g8te93A93Y+w6
OqIxV5xENzx0vyjCr6JyMNbp8FkYV2W7sVH/8Ixrkxthia+EgUdPuktcqYzpv41s
D9zZw5nVzhwIGntFNF9+dNL72cYGRCH/1iaV6wsIAWK4BPe1tIT5BfpdyOw7++3T
cqElx78BOUvmYo/LS2EcVJb3pLI/iYn1EvGHFIit9kSrwX0Q9Q2VCWNJzVAlBKSM
pkyL6k8RJsIwlR63hrdliV9HLaKy29YoemNeo2zdCvDCxSEmn/Y6WwwbO4vGyvnE
7ci6OjAVUHDPP9CkDJ6qY2yGu/D5FA8wQ5PL+udKVvfqwl3/YCuF7JLe4oMzFpCF
FgMIebRGgc9GNVuSlFbLsGHnBCKMp4djXCJYKlMHdcn+znm4bFmlSZ5M7Ng6HTwv
amDXgMLDzjEWVe4YIKDROgdaSex7gG+Z2lBNbW7lZY0KmEhONUXmWK71KDorfLd0
F5nzgYPxwO8nWxX/lsAlzq9LsTrzJYnvrnWIEqU03Uo7cFFoDjvB3zyd977E4wTe
HhW0MVSRNtxQYoIl+lYXiGZkhJS6SL8xcirrwFUpmm3FiOulBCZAXLm0VQiW8c2A
9BEIgghu95jJsjJCjQbJ1aRfejmvIguyiV5aD1f4foHvysIRujvnLNR9us17IPfL
LA9UxQBn7YZuu3iumS/G8MAN3/2sRkSaOewokdwrkM1u+auQ+RADGZ+jOikfNcpI
SWpI2S5W+2eoMTPSM4ZJgN6kafroipw1M7mU1A6ttjDbSeuVpVwr7YI/X9MqAQIb
q6QajPw3YqZReE0q/M3RyfWnBUjA91DQ6WpIxUS/dltNylc2fNS7CItzY1ViKz0j
Mp+YT/HkgFQnDcTWPyfG1WE8a1R81WJFOV9mSOIApdz7TpU+XAqs1ActyjJFoYE8
EcCVj0Wqamsb/82BMAWw/EDCLeSMW1djsGmTLlFrsYNdZqb4m2QWP4jhVljSPobw
5L+1EV7DdTQLIwLvp0DlEIVr0f0LFATFWsch85jKcHRGXajQTCT8loaVCmTrHdTF
bOz/BBOplAQYi+rBl42id9hjA28SnyCXlUctO890xA4hEyZnKhn4n5znAl/XVu5s
zmvBIx/IIK6n5jbQhm/XHCUoi3lLD8Oe22In+s08auv/xyzMUgqb7HJC9M3BAWbM
ZqHyxLC1G98rmflXBptbjA25XqgX4W9SQKCYFZKT5h+7Gquh5lSBhSnQWq4gwjVU
MBcIf+vmrbV0dRonpMh7gJH+MU8Tym9p4HoAsjj4II3xNBOf8ZzRcsM8yhQ+mRLa
SbHoRElYXrkp7C60DMxIw29vc+mAhGQ0AVg1qtGqWnNsuORl6TMX/16EzM/lO6k/
8O6NbTQQMwVdBODRksrKG+WicYLN5WV43P/9XWYAC0Sx42HeIgd7S5+hmU6OQn0O
rnR9460fQClrNmkb9jWWx6LK8K1VQ3M91dBPjrvwUr7WtwL3XVIstDYRNCGN8iAV
7vQMmmO21YzL+rg+9ffeSXXu86AIUcKAn/bIVKxeRaS5/bPS5m8cbpJ0UD880krq
EenXheFUp9VEbam0Y1i1UuILyxe0H73T3APeREmUSnncrRdSRqcUUD36mYhoQx6V
thCJq9B5VlTsdEUycshOPQe5PDaLhZ3NdgXzdrlJ82nhSAiBM/q2LAKiUV2tAsbW
GZPlH4Cf0C5UcTrimhsP0mNEMibj6RQavbn9d8/ifxOJD0qX8mnof6NzLDffaORE
ixbL6StKyZ6ahM+EZOYfkpIG4Q11S1AHJPGdyvgJ1N318x7q6HxXVf1wiKRaFleK
JETt0bqUeTBrL3xn62pT8qBDwp6tfvCEY60mb1UGK2dqCHgbu3VneIzxwRiLS3T8
nb2dkLVuBfVAS8SaIfpOzPAQJgnFDleDN4HzjPJJJQC2R3OWwh6WiG7s2Q9CF6EH
vFDqzJ+EYbVElDXbGbnUwHfCL1PQopBZwXZAHW9lz0mgn5wnFgHYxXiIAV4P7WVB
lEvwLJ1vwpOxYWTpfWi2YRxSOoX+7Edq1M1dyAIdiAlyux43c/ttHDzEd1+95Vp+
PP7Kc/V+7kcZGSRSMQeAF4qX4dQ2ICYppQV2m6RJkJFtOVi4zgCctUpIMkUE7sDw
wzpV+X6AnABUhE/3KoMcPh7CkX1zh7ycvvjdh8MqiuiVzpJ6mlVUL0Bjrl30MGog
zBdgCgw1rtVac9KaTJ3e04SOcB5D2wjGlsm5zXrasOlFf4CD1uED9BVGFEUZjSMI
ppKaRfeqZdF9sqw3agBE6YxpNZekzxU1c3C5V9U4uFOkhrMgLgh5Whu+zj8NDtgx
gOfMigpNUevezowxYXdEwhyc8xSsoZx3osZ/MqLJV7k9tuyjC7BSe4w9i6e2fiH8
1C3VQmB6OXxq3VmMFixyftb1SRNplVW7R7WmHH5f7oognOXlYP52eyEWun3oZafd
/1SG/947gAoHFmBxSA/5bYhgeQc+6S+fmeMQDUzHFvq6Dac0CpsK0b2baj8seIWk
+GCG1hn3dGfnOK+zsXXQ2vz6TcS4gIxZ4YxJgKkp95mCmiuZit0ghViJzenWlUbK
qTtd+qExoRWv/luA2DP0b9hOvAK8g1iKEZSu9QsGGAEiraAf68G07Ix9Kvx6eYxx
oAwrpgOgQ4zo7MuOZIENWWjYQqAWv8ljUAq3Lggy5klhxwD39PMHXDKWwW3Etgd0
iN0LjLRFgeE/BERvw2gxq/appJfAxKypbrT/8YoKnLnABU0Pml6pJr+DrrOIcCfq
R6mjkIMd/HKa/gBEWq7dfSl1asb1X3Yas7olRVsETUidnWrfxDOh+q/UzDmD53AF
RMhZykcNIJXJpCujX08Z2KjLrMBKChQLWt48Yy3qgWcQEu1E4a50ngumRIodBNTz
td/lEqZpDwVVMzILSRZTO0xmAGJS8Zss2NTvgrYO2ufdbMXOyp2MdYWgkVqONAk1
fgDpF4PrN7SDP5F1n1baNaTq5eusGl1mYEBS1k8l1h4HnSjZuFf8g70fcSMi6gAH
DI2fo4R9WeqPgG6xKULtbixfW5HrOZ7XCULMzXbckO2Ql9tqpr5B34a+7JRAMusk
YrwMyTNue+8J38zj9DcU34zdKfNKkWE07Gf9RCBgCOY12XgvIAlUoNOFsxxTzamH
/5IWDc5C2C78JpfUKviEBpziDkpKuskyLaE7hRzZl25t+j3TRnST5orvlrECQN6V
Cn3vIcf8ZsA2UI9hCf6ZXvKEJwRL/5VizZe4tjyTvck6fEbavhl7GpvhCvUNHIGj
f2F8LWqju8cAwW3Zxmqh9M5+YEY7UFvh06oXmQxv2VnNv9RRXOECVkUWRwBaIImB
KwWllTDdGFlIqpAcVUepaf2bO+AolZ2j9lv9o+5xQzDYUc35J8rv+1VaIO+YZjm8
lDCNTAgsfJHc2/KV6MQvSVbQpYWKJghSjykmwqIn0Sram2uJ/kDEM7w4cqvZ0URJ
U2rWKZbk7nRbYOrdAcoT5jOrilg2CvKKPgCmvji9ADTHy2zXhtjvTJLKjEx9O/g+
MCr1F7c3bRVJ7oucID0lq2M50ktT0/bbnVwsicRLvR31XC7yJraTxS3V5bLtUy8T
587fXSUusa9LvB81MD78jdC6g4cfs2Zab3EDO0e+0EIrf0dDe/iCkWmi5iGiCbeM
AWf1EuNyTnHb8zRKyLUyL8aqu7CiolpsYHiEefrZOt5JStIj2UdOzdUP4GEu6ysL
GhkU4Wh7ef2FWc4JyfzdS3bSC4xQj72j+sriF+y95G67ysQsvJHWiS/Ce8jBALW3
NTCXPUdFQyeapUHRTBQyo02BKDziXtR7UB4gNM0aY4Gj3DT+jE14Jh1KM66I0RP4
l4M/FMRakoSCY9KS7kyhoFkxxvQ7/mSYrUXYVCpg7j9dFhJttBEhw6glc9Pq0eaP
2+XYN78MkOIJ6dLwQylPXImYPXhW3Usmzmquqzxdy/9JhUgI2n/3M7J6wTc3L9VA
Hr0YiYcpufZUCSSC1sbEHuRgfWcC0ro51GPWY+AJd2gdGSPfSwb9R1q4wq7CLSx8
1C08lK/gUMwh4C3h4qOvyleQgEhrnImhy9//Y4EFSToEqT0v/YVPhnPQ2OYfGfbF
sA/XcEmraypI2/eAPpPir8T0o8htUR7agkAV/pqiZgZXAEdrrOBzhp+IQgGHvVpI
sapeQEuPBUP2NNMN8VvX0WR0g8DNjsQyovLygqluYaLKyFXP0MeHUVBBKCW+5nOe
CuRrhk9RQU9yqpTU4Em3bJDbYftsMGWzFEs80onZwkcfMGR1/cz1m3WssNvEEH5/
j3bu/p4y4lsxdNlJoRTqJ94wQi9q2tE6/1CFzseJjTc0c7ygwnFyEMpvJV1oFpHC
59wCgCLVxmjLKYUrdUDZZ7wtwqQOJwfzCL9li7lMtJIjf5i3JJy7+eYMxthuOWj5
2eGWaBP6EP0W09hYRfvqMPYxSy+t04MhUk7t7i19mpTTSYmdWcwLvogyh1Rtn+Ok
VxiMSoW37ctw/6eJET4EOE7eK99Ydu4aJgOuy5ujqXd8K5WAZu3FsxiDIXQ5rjzR
pfbIGqCH1dzlG7Eqma1RTDoydbMh0I7TEBUKrpWs+fuIU8dAQ1hqIGGQacUw9iVE
MHKoGgNtHTRPVINb53yMdpZHXPKzkZNs3kgC8Av76TMWd/SvaqKAV+HqYYXAJZja
7MtCDSPR0g4eRuQvcMZgSfpSyIOSKurJwvXxktIdfa/OamokXrkIiviQpI4d4A1Y
86IZcCBC7EmrIi5j7mjoiksKfoASwMskkFt0vLwJj+dDPIViPdpar4rHRkKZjA8c
lBYU4wMwJt+qX44TdNY4kzMRZxIbdMy9L4SmpL71Nih9ExyRbMsuqgTIXo/YNUxk
FY8prydEOpdRwJ57ZaGmDeke+Z+OCG3XDkH2lQM3l5FlBEbfPD7LHucZkFfEYLJc
OZoEv1g/NK4in05XRzzdbmFPbkOqtZRTwubhUmFrD3gZpiEqcJzRk1+1Q6NQiyax
ldhkiI284Z7YY0t6m8MncEZCO3THya1l/np3U0oIcNiN2EqJi9W/681SMsZVPC4h
8UF1b5kQQ+NZiyKa7yj3bJnrjvBDCwz9LH5y7o6Lb0DW1/9+gEM95Quxj2uyoJk7
4dUK4yq7UzNdDhrQf8Y5z7zOIrc/NvQ83y/r+Jq/c1rk0drWqYYzZabC4ejAfjws
IBvkPnC/rB0NGvgmBwnXcrdEaQBHbMjDqFwl3PryR6NqFpAg/HJTtpDfxDPNXcb4
nlst5B6osDbFIjx/4goCmHP6tsU1x0TkjW3SjVJ2aQC1BQat7I84puP99/liAvkI
ILf/+o59mC4H0N46p542eKPy40AkAgUYdZap85C2eHqXq0nR1bSQs3cwZGzEMc+m
99diR+7uuXMXovqY58ue6NcgTDsDsnmTGitJtYPFaaXLK82nChMkzgwLyhKy33aY
qAIz1kdCecBwHY/+sKJQB/jS/BeftuCfamD/ShIzFzPmHLslvl/Jjrr3BeHpICDG
wg/tIyTjrTPmh3qXQOwFV/zHWnTndUWBbZp7w0WgiwO2nO1jum4ZziK8jKLrAD5l
+WR74ep8mKT3+uVABR8ylTAh/HVWPuvaU7CzVogu1rlUGMuj8HrpiCl1ptjMhgEC
4M5/IKhmdVAwTaQxja+rzlmfOwP5PqE53nSobL4zrH/ZGvVipk/198N/Wygroagq
Rwd+StBBRd+77P7p35qEvbzkZhbrrMVAFr/xf8hW3et9RY69B76Zz37RU4Nb+n2d
6sJMCtQ8PXkHlG43LROWIPYvv0BiZXdhZTohzcYDPYykBl6GwgBjO9Qt+NWg/1T/
u6m6SyYLtfwnqMhYdmVqkJiVDXHEDDwKQT5w3BHTKZUrScFxYKu4Y3ybhfNacBDy
sx/Hk5ZgkfbClXNkHh1teyrKEX/FA2X8aSCpcl6/x0AB9oAFPGruBzD2WxoxhM3p
kckUBQwc1i9ZGTeSwuJhHozo9HcnATLLihWt0BCJur/XYgiNYgIPVg3Qd3KeaqQV
0cqSx4p6moOPAadZqZt4h9ECkFrqHBo3xgg+ZEtXP2jiI7yXQFxGrLMIC5R614oF
86RjZ+E5Ww+hTuUTfkP8dfHLbzj5DV8osdMSzxr0Bga2taR4trO3h8+njRWwbuy+
LbSNni9fx4yDQ0PFIZyTprCy6H5w28E05j7YX4RdUPzBP5sXP/EHfB1yTbF+7GWP
B/61oKrg3ysLGAu8kwKLFK/r2NTJp5uXc5S++jSeVh51XHERIei2FLXCL5Sl+nbH
e/oj+oCtbKTEjPKceLwCJ4qX23De9cdLtN6Yqnn9JSkdQ3zxqiAzk2GZTgxmKCBn
K0nGDkFVFJOlYXwZcU1lInI3XY2XLw5xwoJB8by2ZkNfkFb4L3RO7ZyYrsCQJb8J
NAbYQEnRXVQxw81f7f0D9J4/IjJG9al3fLBD899zbDYeF/SVRO7VG8+2qGGfVgA0
Opg6fhACdywyqJS1I4HbdhHOUCFI//bAmjIzU4S1TY1fGUoKnf5GTwbY+jtEYtcY
tORwF3y/byf8DCRVZ5SiSOF2GgoIne81xzQvJUr4hZDAxVXiJx02u8MXnX898pKy
B5sSR5WklvvoeoKinyA9TxAR3Hkn8NqxJPna7gR6rnzsbuWbPAYlum0AhhuOl9AQ
1niuuF42PAJPt43Y2mmKqrQ3HzO0ATqa8DSpzq4XRalv4Pu1Ll6WWeVB9OmkxWN2
ntdElgU3bohI8BTPRtr0G82GFJEiDUlVGbqWFrBNn8mQRdWgRx0RE/8amHDyP95Q
e2Vbde7eIh5c1LjLslMKSENTskCNRLG6mm9pQHGD2aWanGvWril9V1WNWt9D+y0G
o6ew1JMVymRHWmM4n1AXpqY2ZqIXAEqTnYQin5keGvnolhtyGSdk/mdW/Efgtgsn
cgtoQbz2vZoZGMXU0e2vd/EMK8bR0i7+GzSLiHpnqf22HtRgNPHffdQ+L4xIaIHI
pdwjCehIZK8wWieOE1vKsIKwkxpuhyAK08PuhgVMtWTfcUsOkqQ1etn28yhpn7JO
GpKSJu2Yn+Or18VVfrybEME9RsZk5dMatuiLJT0qujhBPQkBPQ6e+bE6RsdXZaWP
tOryYr3iam8efjoLUsCrTzAycvxGuRHNsqD7fhZGfI9pc7Ura1NiHI7G1Sq6lcbh
8g4tDhfrDBmUNIrk8B5m9R3gsSTrRPzej5OedkK9BCOFUgs7pF6vZTzdEL93Nv+A
NVTldLSJmBPHM2mzzA6po/q/zsS0zWN+00vPrZY8oTyVRn62lKT4FXlnxZdgX3bz
yB8NXlft6bxn60QpAot1/pIKhlumLX1VmPQ7SddDwoTLKXx7p9yG7vul/vHpooS6
u48QbiJoA3LBz5ZX0u4CjqTI/bcDQLepchJ0CI1P0Ic7lBHSZrNAoV1c/vAJnys+
GLTHPGsD+QkHLR+nydKMQTf0R6YRbVnlNWTrBGnL18Tj6mkLYHDKR+W7cMtSja1M
zZJjQwD+cgvBKfbZ2XF99phwFX7NO7Rj3/G99s24DiHOVcyNuiBX8PcN2uzk7kqh
A8BSOdizwk4mR6FZCMQZ35SNW4yWtPLg9JjxzL6EqMLWetxwnSGxpEqMBC3UqP+d
rlk1vUgDfJynYa8jEs9htlGDDCL8wl5HebMAhvX3glO6h2vazBY+2dER2vmC785r
YL6axhd6P6MX8Tnsa/dv0Hd3AD2XvoRK6/fhN4+xOSFl8g/gTeQZkuffmCvdZRTv
knUKalV3VbktZnroiTBcVyD07huJzc3KZTEmsFimGcZwYvxc2kaYIOrZceDZfYB/
RJgsSSQ6+HzSPm9pup77YpGKvqHfECSnylKm8IBh14/DwwGthjJt4yczb/zwIrTI
GvKSMczMok1et3qdNezFyGfsrT5/hIPcBVnfAduK/jbGQWZy3Dthtym9T2RDY1yO
jUQNT5rMG7/5gAzZHojYndrRSwb38FLUxUuy70hGyVlXdLGLNjyO4Xd0KWpTWA24
T/fTjzWI5zzflbtIjvJtKyZn4E5xyUGUGQqZkOKmQZ+o2CcCh6bx9D+SaR6xBid4
C044UZleAmEVf9ojkRx8qVTihkiv6iiuwGivvWkJbTc2g4jNQgF02qE1mifKZD/V
pwPrtDBe714qG1AorKYEF64hhYeegOBkmwwTzofRCbgDzVEqKitYwn4I+OkWHU2J
+eesYsRkV2h7l835un/GSsvYQsnVMV5ZdDWG83JjBxfo6rLsznXrB0Z5/vPBl6et
Igz+Kb0ZirgptzbF05JboDh6Tbq6lIFpAdHZH8faNwsTXxkS/Qpl8r93o1roSgAS
cB+76ZO/ZNgx4YPTg4VFYpdeU7ZDKX5sHKGN+COS2jAzl3Crx3bRtDM8AJmkrYs0
Lt3Bii1jhkBMq4VX0v6O0DCt4oU/mMyaysh+9pixP4iNEfo46zcDnnpe+jpHlwTV
l95upm6tCNZcWA/fzmdtCpXilvqGi136mhXYiui7MKCh3OEcjMNBTnFU/3y9hfJK
9G5f+r0rjZDVJqOAcUrPwoeWxEIkZZ9W9rJqF+yh+5v+sYiN7cDDK+HzMw8uFYFq
m9a71Hr7yRhYq7QHe9gQpw6y737RY1WhtKILfUHFr5Pz5ifcQiu7WJfM6Pj8we3j
AqsTs+/+LrMpdFifcPtfthA5ztotKACgmtTAghNWrT32FLdZCpprCjwM+fK5UbkR
jik783RYgJAqbT2C8vNoGIVyuJhw1H7kWVr753PTjkv6KFceH/fy3gbNyu8vPPTe
KIIO575FrP9UwjScMHFuwy8fNk5o9/tMl4bJggVmNDtQ3WJY94HRPoVu8z99QgzJ
m8PdPq/T408wdkA4dKDpFE8x0c1Kxdrb9t3NH1j6Yk8UtH4Sku3LcOKcKa9uYDgk
Sd7fNsmWFMGr+h8BdtdL/dg1KFpZBtGwC35fZZzEgCJ9W0yESl5HpEY8fKam56k+
J7BWZl6Pomn0rmfgXgTG7tDCEhDurNftKZOARJQde0dgMPCq9+diN+YlBt8kIDH7
Ss46GhZMCiwc6fagSNkjZadN4WhDzPsjP/WHovXPRiDfAOec1IaNbNq2GKAZwjlq
jibTzrRWTAdyq6x796+WVR+fokRadFFUofwrJBNw784IbiU9bmemMmRua+3JeHfs
E4ceMai7HqxwdSIAWfjpKkMfh4l+b4aNYCEuJLXUJ6P0nxgjXjwfkrCdkV0d8T47
1O0b0htaEXhvdKgIZroAOba6K11bahMy+haL4jQVJM2nlZVw3d4PAPeEPewBpCiL
a/Q6C9j06LPTLQfra+i8GA5A2rIFIkfYTDbNO1kQkgPGXW9OPDIv0jpsAx0Km1tC
9o2av3IFl4iHj+04szQ5UzhtELROks42L1U8nP5AZYwkOZwHeL/g2dxgJxMkVQvP
zfBvDhS96mX4mJp7D66aR53bTyh83JZQbr0ynqG3ZjjuDFig9EtrbbS2THSibvCU
6jZi5dCnVLfOVWMP3B09lATjgG0Lp++jccEvN1F99VjVCmK3oscD9C2xGq3HQwh/
WB+tpng4PkRJF9LdySMcnJlM5EyjezJ6Y6cK8OYZpg2XWCsxJ8RXkwrV9Jaz6QdC
aZU1j/Jyej+FF2uDc0R1zQEf2uPVXtbdxxREiQ+Qtug3OwbdLf3jqSHPHF9xOWge
dAW/AROWD9QUyzPxqvnOotHDEBFoj2SJ5AcFM/p99X3ikAUjGAglZbPCxLl9RD2H
wS6xcUEDxlF8LceTvelh3UgXJ8ip998QzIgvnonSjto1qwMkQ2+3Cvzd123nwliO
c3CjHcOS4CbvJE3zczdUJRckxGNKEvzhA4O2aFEcShRGX6nEJUZAxYDRZwsez4lO
pJSbuNizNVSh5lcJ8uPo/UVzbkVYErRQGfULF5J55kJCza2zimVzMRhQaLju2MSZ
n+MqjGaTNwlvbyzeImc6wdSMLt1Y2EReJtiMfV0uzpYv40tkoIFepNwmkwkJSDzQ
a0/Cb4wZS7dFTxyQpfl3V3LmjJXVRMWG/Jda5JRzz1qmfSkRtZ/0vEfZl+eeIiRk
xirJoHiuqwkW/DlD4ToL2+8p+0tHAfnY9dBbr4l72URGPHmQJas197nfpZEpD50Q
NgOxo4SeJx5nZIIFlgvoOzhV8ki9yQkt72Ux8kpSI9XrbNxPQDsMMpIkemvDPayl
oSxF4V21Ie6snSQcCcIdOCn8zVY5M+G2QGLW1inQIa03wgUzMQqZ6MNFWvc1ahkA
jTNnSTS1kehN/gqFojGXJwmMSaYnlbzyi08YPugi4pMn52RoAdI1BK7Iu46+zwDF
pJ8kcqzyy7vLjUBEBR/QxaevZ0tW1nabEbt2lRr3CUMrG+hLjV4gCPO+RPzzn8fP
+dxaU7AwgNmkyMmCDjNnBbuLcptY4S803ejEf/90rkxwen/q+Ry5ZTW6OSRFcUxJ
TwwU7eiUT4p+RUDv90qz1PxiLaJdNxePdhm29AK8lyawMHXuuQry+ZQPTUbBZwVk
ek9CZwUoQiRFewtAO+5dL//vkiJ6eGMJNVv/stYL0R9XmPiJRl3rtfP6xXKwQ+AL
qASUAOdTMx5ovP2K9vMK9InE5P2YAXUhc9K8hB3Qql3DvW4dDUkHS1n7sG5NbAWm
LWRXhUDYsTgqEXDIc5N4UdpdTE0WTHgATZN6nrkxmwx/g68bLJezGWzg9FMms1am
SMvVmSh6fh3TGUxq8hGhHZurLr9LbLzshHeQOZcB1SJyf5rV0856RDaXcaxO7HCQ
yCx1LzfRq3iymp2QfKk58Gl4eDDYS8PiU/LF2faS4que0z31XP1NDlfe3EOfJFDO
PhFlmmu6oQN+/JFy3DXvb57RvpS5mGeoZq9Y0kVY2jptJ0FPHvuluJdc5yVZSkRD
I7hkH2XY2e+rvo/gtrziOZ3wJr52ifbmXN8bW5ZQxqhgzgLP7snRHcYoZApcpx36
SHABD2k7FgtYU2Hl7p+84ZLZBfQvtZsFDFp5MEyH7ppoKETz69u8f8w1aTrWpkHh
PCcNx+aifc3Bxc1Ub4Q6lGQTtRJLDeGXZTDh7dYkSyM5vdj20TG2SkPQfGnJg5tB
LoxqcQpZCDp8oLiO5Rm9BR1U2nqq+JmX6JOgIIto50J791fCmr0Gng7uN1IfzUlp
iWzyKHOsuwe01tyOqNqodJWaIwZ3OaLGG/CpFdcFsO6lUxg3hFmvVTqtdEVJ3DR6
k8WQy83iN82KUPMPKBE3yyMlu/3/0LXNTwR/hA3s9f/OdATCGYzjnxUxCliF2QAV
Y6q4ta6+pk4VPsjPFPy2N5Axn0Y3s/lYPhIBli75T7upfWnaY0o2XRr0pbivp/a6
dSKI/PX5dTMDtFkCSluBikWb0OiTEBte2/en6mgh96gsuGZI5s3Vp2BTbDm1fJ3k
cdMnjYDD50yYBxlMo1Mtq9gK/dmcBOWr2OSaXbYOEMFMIhcMQDU5CFBXdQuooUr7
xoohk3RJMuIYbMWvYDntliMlB8M9ZQHm3NRTcXeZ9tKASQMZaUjNqgfWrlD2xdjx
2SSeXOjYAXwBK1r0JO3TA/Ta6B4W3gMhHOsPu44vt0H7xOQRsRHwpgU1Hq5HfRPS
0OMTvDR4Fllp3BUlxsXUjMYB4h5sqF2QyoQhQrBlkAi21vaE1YxbUThNgP+ILoOL
L9+HiCOehGDlAXsaGTEny258N/qAAi7+rMjPS2smaY3vTvx7oVjVMMA4c6FSXmjJ
9ZVZ5ReGgt9JfC+TO0ZgJ8/SXwo+jY0i7rfTjUj9PQJCMJPxQPjGUImrjLDjeTYe
KwTDW+CH5oyAnvhFDLwskZUrMxMjvNe/lTlor402HM/uX66KIwotkbjymgCIRlr6
HMwRx1qOOIDME3t8p4rN3OpmsND6scOvehqzZH3/W4GG2ojqK6n22iFPgwrfBaox
27WHBBFMOL/Y80faEi4FNupCQ019G7cO+Oex6Iqd0xvgCVK+qx2JhUX/+UKwsW25
k+UOh6y13m6sy4GFrzXkhEUqKwCylCXvVQoI2s43rawTimwO3eeqKivB/BC9UcKL
lPhuYADzkPc4LAOyztazNTSO3nofkS42wKw1n8BpOl321V0lphwvaKY58uwWkkkV
Fg3ZR+K+jnqaASCmgabERf5WmpdfGvDosPUM0A/si+6HsvHb0K/TBGXFMkf6CzfU
kunWsKTYafLxyVyRrPlgV9gB7k5pGz1k1VESFtaLcZJAFldZUF/JJ8mVvUxYwBGv
CjlwYONYuw+3v9DiHdhOgBoWzzt8Qu4898LcEE55ruJ1xv/Gij+Ipx4lFH7Dvfid
ttcZaMYKrNfmQB4n5HgZsBiE6LK9dsmfeEjcrXsyS81BAt+QFRb0Ys5BJGjgcg6I
SvauZv4Lf6mzw95OzSyIjBW6Y29OMC6HhtN957vRhWtSA65dOmIofML4lv6PcX1J
a1aG4p42qWjj0+6k+7igvBjigzm9t44v3CYOfC3m3p9pmDlekjxhZkHYWgL1qG1/
ZLABxk+cTO8KX8rcuonaZuSky3uiu1/AedJjM/w8HIrlDMiVHwvWAnN132LmdtYo
qaTCfT7HNuSoNw68+12hzkMi8ydOwnPfW/9cR0rZw1oPrA1lnXV+4Kc0Xx4awWW9
1LXPcL/szVBZxZIYJlZnK+nLANrfHN2qpIMG8DJW61XQMiQVduvEcoKfMsjTXlah
9tF9vb6+L569qSwYwmuVL0yg3I1fLPkjCWgrC9iSNrjUYIXA0Tw+c5T4WbrUA287
BTFpq8sw9A+fmMk5Topx2kFRL8FgusXWVXjGOmz1V/VH6MUAimjFhqLIKkJvc6Dk
hgUueAptrb5IIIPxLNq67ICnWTU57gft/fi0k3ezHvYiMh7AFfMQ9EcLfqoPvily
mVSgtn3NiG/HYz/xaQBFS4gbfNb7Ju+DSyRP3LJup4M8gBfDP6g38Shnv1CJ4vQu
jI0HzXluuNwUU4e65dTGP2nKohzlY9r+fUBJr4B0LuETxox4d+x2Qd+wuZ6XF/RI
buI8+Cz4xLyPUU2zhWZbOZcc5R1sNX+opuSLsd+fLFOH2pGlsEhOGBitnT129GBp
lLETET4De7b7RJBQ7AzmKZLSTUjjlCcML5cNbOWELMg6AZqzK7w4tEOHExwaCRkR
n7FFFH+ax6J+fYM1ohb9nnMThKP/64Vc9v0QREuctMjTkft90b2rJePRiPG1Wywy
yz8dHJPeTo3QcIYConZPenQtrS5+esDeEJwzdCgWwd9wit8kaq9/ffUVBsgz/xPo
hYl04VBuyOUfE0XsXPmPADcXYma1vzKNElFi1Ih2txOh9xhXGgSn9+c+Z+Io1wnL
ob9oioeDXe7mNcq5L6EAslHgWvw2tVczWnDuTPe+qTDZdrC782dGHHklMwaUjqnV
9tNgMixuUBe+9aFpW31Sj1HDzuDa2Je2FpR6EgqULCHVH4YRnS6iszjE3X8/ztjB
QvYbi0WCVnjgZlKhccd2HveX89ZqWxEjmg42V97/2thbwfam+Zdeeq4RHeHbAd6B
hWWFTJVF779GWt09he63X/xKSbOXyb7w9OXMZXadV7BHL8SmGtbEELuZ1HL5js0a
pgA6x/9WNaf59t9o0irISUW+rerAhY+ycEoUFRvRs2tLnMKckYNKFeLcuktV0iD1
yRwRDfmrAtaZ8A5xNU6fn8C+Bfuo1I348x0kNquoSCyrU1ixEYiBjbp/Brv5bjud
bJmAD07STtFqhKHghhP5qkfX9rAdfOPmFB8ykuu+cPfP14jaeQAYIsBza/KdblG2
QohvfFGBUvrYm64VYmwCDS5GgnyXbNSC+VNAjOFfHGU/Eg/+Ko3mFZjT+E1i5GZC
5g0OmWvyx4pmMFzCVAk2F7KeA/2D1iWsj/xKzAhi4DArFa4FIGRNZTf940Xsh1Z7
sMKubxiedET4PlTGbw0XKTYQxX/8C2PX1RVgZ+UqfhNoJBMk2Zfq96h2eA4BN37/
d034HRietxlrC6mV2jTMhfiiErhKTeMVE8naaI/W8vQDcPp3zNdRnLyH781rA9PW
qOpI9/4lkqgt3qWwRcxWjMKMGXcJc2axUenbduAVdvHhtVB/XuFW+/Vtedfbg9Ae
K02ROSHq/V99qLso1lsKHITvp0tCM8vQOnnClmmhk1jvopdAIHZ9REg3bwzVQ/yD
/ydIk7AuuTFB46uO78oMq4hnYMEjfIIHFnv7gZpoKa/tc3u7CO7hKpEhSoDchFzE
24gHbTcMVdsoZYm+ruua8SGlmBRENAwVeEG3ht207Ugkv7IXLjkm5Fahr3jA8fhd
Dtg8smiDEx+BNAjNFeR3Q82X/s5nI9zTSCPGMPp8lsDbQztaWwRb+Y//0JNFaa2A
7BG/tJhQUKO/TEsnZFJGQh8PblBoFq2KagsW3pXfutTNDhstz0fxp6yVQk8qkrAE
MfAmQE3qE7F+x/ybgEPNMgvCup4Pj0gGPI2hxbGzhFSiveD48QQu85yRmMXu0BNH
ARlvuPWc3DFfXiLoclZTIpTcoYBLFYruXiy8r4EO9sFcQKL4bdeu+S/yeJv6lxXF
q0ocVwSqbPN4T5DMzanV1V1fE1ArMKULVjt+r69D9xa/jwUwZdy0fNgkOk0P81fv
H013O1Q7MTWAWARXv09X9weg8jBl6OPgmW7Hp/ff6AVhuGJA/PIg6d8+iLz2J6LY
B67xdRxAv22DSdxD5tgkpgTm5rhReTEGSdBowMO0AxDdjfvuoolptMEcPZnA8kP0
LVr9o9iEoarApwf+N7UzS6WoCPGfRwmAKRkZ5XPid9plIw/HI+AaTKMEiER34s2d
p6xJ/yGrYu1eg/jPR/RNsb2UsQtcjJj8OwRAbJ2dJhvEp8kaxu7w1zb9qGHd9+kt
pwE7Js/DcfmeT1xFTRI2Yi1y7xN8dg5jOs1znMznOMkxQXRDoa05+ym+24iPhOC4
VUH3x/SRlGkd2owaHR6Vtoo9G3gkSPEgOiZ9qfppOTICwQgfis+Xfd8GAz77CTwP
I03hjIHwaG1IpNSwWlnBIrICxtSt7AJaS0AtjcxdmA1B06k83fpj+a8S58ClwGoj
4ZzI3HbTCmHVkVVFbAWnVMOUXe7r3nxdxukWYzMGK8vWdUCRTWF035X5B6FxCY5m
UlT0Qb9RjTqR/ocV95maC69waPV0sYpdjJR2leh2j3X1/oyzQDnNpFJl6jxRQWBM
Q2oWMSSSKCx0VXdDBv56ckU+1ZkpMQ0PpzjJ/sRKD5HzyolWlDg2zfcVNOP89NaG
bE9aN6pnQYXIBZAoF8wzTRK+KrwZn0BlyND+XYsBajukzr3YVTyquh51EpdUABZD
/rBZ39wPLAPhdvyAPpopJhM2PwIvi2K3nJinrDGAY0f1w07D2rg7+SWnXpMWcAKX
M8OWbYQ8/CSSXr5SXBPJrPbJe6eWnwL/G6Hn/OPCsrRqC3PE+rf8xkzYpyyuK22q
OOEkIX0d8Pcg3+1B2Ng71Ox6IoP5IkyS9EuQwRh30wbNAAR8p1IqRxNG+e6OuECG
nIlaeE0LvTMpyRwrIOmtGbBVG0+V+9GkXQSCReX7u36JrQRlmvEGfFAzXU4U0GLJ
i79XnaCkAMZDbQ9K2VgNe9wZ0PYhL8JLWNFNN+IaD2c+jkboxYkvGcXMnFJL9B14
kwGVBHAkWsSRzUd5z+0EheLZNJi8JqbY6v8zpdgPIBN9LolviS5PXwizCQ9mHiAM
AsvZKLMHgyhFtCOZ+lkfQOHozALxx4Xh4KwNQAn6ygbi3tGr4rIHhTm6pNVXzPXX
YjT+8YXkCEbblVrdNGnlKBlxm+sLUBsrYm+8tk0gCe10r3fW0f6fbRFMcHB3KkfM
AFy3ldVmA/Nc6XMtYnKZnT/WZzIiMO94ihyhPXoT8PuRD+iGvHt0r+YlVg/iJcYX
+EjT9/4ZRO0tIyn9jOUkXOLY5DYOFSP65P2negYT5qUYGAAv8Olu+ZYpuFE+OuYg
ByWzsf75GSQZpgrQKAj7baxlygm/R3mbu1q2nViQOxIwPt6tV4J8yo/LUbL8oaXE
C9hMJZOBFtvVF4YCKF9MvwpqGRHV+JgopEBKuZeHvNROiouCHAjYDmybUx3qABSE
0BW6Opg6QpZpL5bCoie6q3dBUIUmSPazPKEOCuKLoq7B4D7CzMjsxng/EQMtpruX
RoQSpAcpa3dlUMPoJfZ7A20JoxJXla11nIaTUP11/mShXWQLtx85VqWBeHBZXYs9
0ZjgWmN67pqwodaNeu6zjJiISo5DI/dSvusram/EFZ3WSjKRSii0OeDt49vpb97l
dUZ17by1djOi1NgM0djs78kGaqcrEB8P50liOeWCAFTAaXSMzEc1ji+ChcOWr1IN
rNQg+dTq1Sa73l1J5JVD64tUEDUZrCAqvx/fYOkcT+NVncSDFqOgkJMoNrYlwHxg
+taStZSYazJH9897+iUCv+Oj89BXmp2e7h/KNMc4tzK6btkqnqqZD+ms2cI31GOO
m12YeyLrIfj0aYdYoO8+zZwHMVV3w5nmR5v0hfJLWcJyR5/qBzdPdndVZdtR71gg
FPQHCN1O+YiV5DIRwKXm/9xMKN55joV85vj774qRyOah8ZJLzvKR+roIc4haM4li
smSosZnS3PGmbne/uaUV8svMQ8ZfwCix9dwh6UV/yBl6dT8xwfRWKXw2kKm4iW5T
aZK6GeDqPtp7oAu7nUcT7dvLmNV1UrrPScrohJ3X7EFxfpb2hu827lxlhoe2jIsL
uBsXlqLcgv5Q2A0eNmtRY5THg7qHt0vp9G60NktO/pdYHpr2uREBY4+CBM70dF+9
PTOCMUsEmcd06TzMRq0YsC27m23Lut2k+wVfnFmJdfvNs2fA+2P1AYyFlol6FtwS
TWUfsXquvR6lXL5VdwYDd0subkfJvwX5PcEpS3kdC85WyR9lA9p3vpV1Wl3EAH6u
NqnGz/k4yPdFaX0xxewKhQkpjs72HHhuu9Jh4YGZ/ySdU9mxvKmsFe0YCJYb/jo6
ZgY/RSGUnY3va2Yq+Y0SgJrhYUR4/+4eZP9ZSs8YTClfrRjL28wD1fm6mQj3G/PQ
8F/bWWyA7VTL4fINbHAAiEy+xO6CxIzQXkmfOhzVd49qBfcvPLB37B0z6WNF0j3c
knA+z6QqhEGnCTm2YI7fSNmIUGRlMVxIO2c5pzTNEvf1wsozbWVytfwePPHWtoa6
FcGQdpH7POH0wup67StROIO5NYhg+OqLzTrVwmeBXyYMkSQxA10VoHKYjnD3/qfQ
qKbwbKFX8Q3A+tmGA8P09y1A0Vx+GYVY2Z/Iu0cTHBHEM8fvVSGqL/RNJsiKQl8a
3n+zQF+nzbb5dT+0/m6ZMsDMT52zls2n90SVrbDjAZr3A6d2v7KX0kPgMYiRQDO7
JfHJLz71lGV8i34oFGlc3V0eqI6KhprCwxhnsSiSGQMO1p/QiU2aw51izI6/X3/e
IP6GTOVU2PzOilIm1L7SABSAFgF5ULDnFxALlrSJkxUv/nJVnvulZrGRn4CSKZc/
ITeb22/yM64E9Ww895SGDiESS6Rj5mA9X8IONhhRQTAAG+Kbejoqw3tprppZwcCS
9y6tM6LNKvp9F4tYdDQ2m3x2E/YwWSL++071pBJ54fh69WC2RzaMbAWdE68VeMZ/
zC5p0AfpDgYy4JLCuIVOiFFHBT4guaDloA+VLM84q5josEXLj5b+QdSa4b9vltlY
uj0FKgtHGDDgo+6QlCfQ3ovIwszu2W1obQ9yjgQWx4CdJGuRDIvDc5FDOn0jH3T3
ULr4hBVkN3n1DvCKz5ju82Gatl1duMX/CCtI6GLVhNecZCBGoA0w828ksI+C9LqT
IdpDTBksn5OX2743lp4yL+Bf/n5tVzANE95CXPHGmSzA5Qr9z9+gYMRohTiL9Ya3
AWaNRP4df6o0KHjyL4h+PYzJkbRPs18xj/v6LLy/NO+MpASgxhIHEZDPJHKzPF2E
c4xwDbgci4RGcpjV5Hzv2fwMVUPw/clawl9662XymlwSr8QtRpWp3cRUsxSrZmz2
rf28SiyUEvYQIlrf0XSduJBes4ZMBX+DsS/rVraVOBGkNAgIXWLEF5VITaIK5v3M
jKhOOeDEXD2ihko+J5XPE0scvhxpOTb+tAK8U5XqHSecQVcO1IpJXihh7/zMeTzs
kXmdQNUVutQurOPY/1+Uncj93x+DCDJ7k19FKCLnkGWiigpFg1Qa6G+qgVCGq1gg
so3MdRBymmwWqfkMb5kgItX+bxa0jv6nMaTQk6IHP9lTvee/Z7NMpovfK3z9HoLB
T6deulnNZ0y3c/c0IZaBwIVo95oBxqIm4b34SktG14ig6xmNR2yk0J9TVdXE7u9m
/L68F0t1a9QoWirNHm6Lf8yQ5XZh1/BP9DqrlGgBVhdRkrIYM4DJw9ax0JkoJkP7
TQ/2+d0yuTaaYlt6Oxw4lGO47d2qybSLnjJpz2LsNWYc9Wl0Uhdkv6WWTeVaSKqo
c6bE6nTghvWaVyTyRZuLPB89P2CpfBE7927MOypzq4YRWYNfQU0ivxj095OVQ0jU
JgGJ9LSgn0rqWzLmeAWeY378+G4RE/yjgyo+uJFs5FqcLHz1UprNvHTfKzdlwmPE
K4pw+4sPxqWz5pRc0QArJ3FGjVciRNJ+ij+rvJIrz7HlEKKmvW5ktVjrp32oke3S
mgrafGH5e8sdm168g1asEL2oHxvkhN5zE92oteHQIkTv/ndCKpy4mDpqFKutyHSy
RMLE0KVaMmXmK27rF3n5D+SwKVX9+cHNetMLg1T6fk8ETMWlx2n+vInXR7NVI8qH
TlH7mlV09S/rk0X3U3Rby1rF7G5LN1qWnFWEXEmBEIGV2H81p/ZLP95vD0971hYd
fZZjMvblV6gfNYjxn77BeOd4dwazJQ/Ng+OwuzxKoWv0VM8E8L/8X1o9oRL/ufAY
eW69wbL9gcj8hLvlja8QqIEfdGAwhko2NGV0cZDqjF1aBYBk4FBj2gr2jev5sg95
idBTRpnMYvWW0s1G4uWpBcsqu2sVQchFO/5+VtCWzgqclbSDgtqYquySjBdR+7xM
3cQQW4gPp/k3wbk0POHCXD87U1obH2YcOau3qGkJuuZVpm2xseQOyFA1qXXUtapO
Z7AHbormwMjhzVqV34tdeGxMD3IOmIZLGk9f3PzdR/1bGuTX3ShW2XuZEdFdsaPT
jlmzLHXV5r7cHNak/h8GjvsXpUTUMQm/rlaGI6dA8KdTMRi2YFakdk5ZASU3eHAf
yVfc36h11j2ozdu0CoNx9+kYMnoQsh9uaDsSrtTrmQYZ+Ng1eDJQ8G64mzxY1HHo
08wmTA9HFfuMHJgHs6e5rUQp3BkJPCT8JvKOCbh1eD7WtU7EaYgcxaC46/Z2vn1S
aZNfYMp+QIa0sT4qSlzfywAzH8apZ2JJwcSWt1R2aLqkTbyoXsauzdW04MPMFEKb
mfP9ABnG7KUpvf8iamYL74ZD1gMfy0OUhqD+oQ1lFtxcoEo3Z4EqQdCA7ZjyGk+9
M3fCWbKA2FxpgcKCNRswgmK/vsCwpeAgP9UFWTMekXP9PAN9nJbiwRJ7qFnvoN2n
DvcDXhLLzOLpJIsrSRmPD4edv90BfIZ3sG4dghApHKySXNHlVNGI0zmCCV4cvdIM
svcl5+XRj0gB5oPMbTThSRKi+rQ/eC5ongvWZUoxn2D3XO7e+QqkvQ8/Hu5E+tEx
JHO7JV1bXsDpOL2SDwl2WCa8my9OHm25aHepAC4v5TcpwxbF1x6kkn1OKjLS0Ydj
Dr0ScmdpkCyK4w4ywa8ZZHJbRxZiqp+PgeKQ+BzONOLjQTRLogx9QauNIpXnj+Eo
u25l8jnPQPH7QfdyDTV15GVXoJk5ZIBBC85oWTGZDx2aw5rnOMNln1DUjSP5+q0+
69HUk9fr5+o+y3crvpv5JXlffpOxzmSYGekle6zyJCVOCawOgGr2AKghO58uR9Vm
Ldkp2CVpEe9fDFnjiEzSg9rPx1V0fNoNRVcFtYdKdnMY/4zRbRZEu6jdoHKMmj5k
l0TQsfDNFBWEIPrpWfiDJfcIpvlacYZqJPwbCOp03ZFTMMH6r6cjVvZtNycpBL2C
XFv5O0e4iaZU7/LAc4REhM9XBpuqQZqzwcjFH4lxZAF469WJ4D+sbBQn6372SCG+
JjjP2cFaVpP8kCM0Bw0orUXgNA+XSLz/xPIBqjZM58HCIEW5dEDbBUP0qr8FNkQT
STa5SLjlWujGn1h1Ac+i/LYWuVv6m5I4we7WDkwT085BpAQj1HrVQAJ3fCaM9yxy
h+TjjYP5XtaRLSZzn0c/Qgz6clTGQoWiCApT1uaur/s8kwgJgneVOl9a6Z3LcKme
sy3uIk7J1+Bkm4lIGdHzwrIhsUkAkQQLwJ5DRb/cu0ge5L3z645GAcVcMQygVhhm
GCuoQdxDMYhRqGOGoFRv97f+yZrKzrdvZKf0wIWHcniAw/W88ZJ6JOlDqw67xA7k
DeIEmw6IYryFuAYQedUmeCIyzZulk21Z43Tcsu1V8D43JZFCiKEaDVoZbdtxWCKu
Wnx36CSix/HphN87GEWIdm2Rq+RuPQjvIYOT+Dv9/OyR7ctpRY5Q5xAIVt4cAI1o
rycwU/Lpn7lCt00M/0o8Ms0RXXKj5Lcxgp1gxMXjPGsGg+oR3vXWSDoQS2T7jTth
3G1x/aRQjQdoEJjn/l86HXlkbn2mPOgR2NaXHd8k63nRO5WE9nQ7lgUSwJFcZpKD
24SD82W6CN5NV4idjdK2GztlLpHKuzDwT8MvsRN8wPnVMVgQSWl2cu5EaYbc41eS
Nggr8jcsbbrXmtCg/UFF3bm1MnbkxIc6SkOajXH3Bsy/IhBO8pErgCCT+YaTDhyN
u7xiCZJKsydsGtgBcEaRf+Y45kxZ4NRp3VTMEd3dDWIPyMLRrfO4lMrKb45ZRhb8
PLyeJlwd6URCftwnXm+ySfCNosmrC6a7lHMOiO7dByLf1gKRLz7vmrI8lJ/Tc3m1
FbdbUfnTcAYvWpxKMQRQCbsgQeUjf2hDnkfIVD9m2x3bv9Y6YDNXGfk57Y0F9J3k
jJfKlg3tYo5UIUTNUJeAURB781xtvpPEScEomEK+CZY0V7t9BoV3YzP1TXF2/trW
ayYOnFIIpA1YZFLBxWggZyhEJv6lS2lRHJ1lo2hH3g3JQxnpgCuq2ntV9FwOYh4r
B95bEAFVIB6PcebqVHEeAe5DLagxaH2AvJISc7eGg0J5Vrsuh1GUkPftsMROBrwZ
LNItUrkyVaNcelV31uew1gOa+FZ9veZWRRKZ+TqyIjJDh4lITrEd3Y7gIxkh4TnV
blC4WYJYtex8aYzYuDtCWCmWG+dJkuNsphoVPcMiimrLadODmKTvnjqy9ZuEdyzi
uRh6wdyD6UX9mnm9enGct5J6/5tkvwLJTLUytC3vhYyQxoaW4+iZtPqlyL1yOLpX
8mqnDwAfCVhGK1qHhVxhBrPK6bAC+riR7txkt4/U9BDft+cn53J2bXORMP5XDM+q
JfYNEOF+k+7M102BO+vB7O77/oAlUFMRhfjq8rmvM/Xl/xhxEudpiKCjI/rDGCPi
Wzyfz8N8Nc1UyqRzsxwmvETd7WAiiKWuSgoIPuZOmmgrLEM6aAvAh5/VUkReXl8T
wYmwon6LKjqPPv7G6ETq3T5xlLflXx06LJf4rWJY6bZp3t25cF9bbXC9af1i2EuP
2uN8pZ35uA4Okd2YTCXXFgjTaqm7JBQ8CoArGAmCeSmr9CgKGX5x3a6LgK+iuGpK
SipXmaeDKhbZpt/BR5tIgYsphcifra/re7HdLPrUhD1iEmSaD6a4HqZk/5codKN4
9yIYUvRxNDu/damX5QqTa50tVwWcKYK9pQ+ljd10qxFYH2W1r6nkUYM2UzB4xDwM
Jmr/OnDpGJhxmjPiYJTbCxKfQ3usO2oI9piUEy2FFB8uO1PRP6gRWRSjEgFnE2uQ
pXDGQo48CCw4IJItJHvme8vWiDwp9Ia4+lXDZDjkwjcoxKs1xegya4P/AjaWoIpM
+5CgeZwKGLz6bpHJqOWhT3I5n+iKErIaYZV3EZIibcZo4gZnEd6Iy3ZJU2SYmAkQ
m9+uDVtZ6s+wnCPYn7VJJFra/tOe3Y2DJ9RhWBECl3fREfMemn2XFE0JBwRbGl9R
EqXdXrW98XYP3vmeQlYzht7UJsb5pV3frQSctnnHCysvvyO9R17M5t1u8Bz7V/yc
9BYZ92t71D2eWb3GQvjRGyIBi2jmwyKUPJN7dEOze+W8UaD8pKjU4TBsk/N3b4x8
IiWd/QlqY5LDHcYSiUzqYRRD5H429kjsyAe5mTecfZYXfxAQhN6KEPAUMUf3DXXy
mI1M508YaTVnX5shXVJar3bUPrgg7KuKED15lmUXG9McGWIHumCGbyfkI6K6BY2O
1Zcfoj/evjUSMECJjWSZv1CNey+UmV5g4OLko/gaPY7jEAoxq3ejTOiDLEg1vfkL
ttXnEvvvPYutIiYK8hxCoyWXTRfWSC9JDllNY3eP37PzpwAGHjbvc+09+w9cHV38
wKFjA1m2TXrf8s9OA1O+6ntAzHfzZ32BG7V0+1ZrLaloEpSdL0NItllTa3JFn6mO
O5PPvPfZGl312ldfW2Xebrn/9z5O3BSvA3THkTaOLw8Zoor4XWyONfyjFnlpjhmd
TwIaM1HqQ1GbwbVfBpHKzuhX7XDQG3XRyo0l5SxCnEIMt43dknTQ3aw4HkT5A4/b
pV6EG0SspBQRBOipcPVA9ABhkEYI3hWlUPh7JiorFATGPAil0nB+cgUcR23a+x6K
V8UIEpBOGV2VO2CIiaWKt+uxexdp8qC8Q7Dk9mBMJMLPAhc9eaizcRqdqjErwPy0
yTdbTwALdpPx/L7CVjPbLBCpBMq6fWdrDqF3Vd/UjAuhLAQextroAASa+veVucAY
ekexWo5FncqW8SzzrLzoAwkNKFvGjkSPn3a39/Fcphvxvi1fCJMst/Fhk++3CufM
gOxVbsG0Mia4cz11ieuHtnlv5c0b+RzbNDBa6MKyDCOZycYBFlM5LEcK9zQXWFeo
mo6lUOCcwT7ASc/+B6iavEcGAWxmACHmg8gNRtRjt50LE+HcCp8cfnhRPHKon/4Y
2yhTIdmjKC96jqqgrp+rk7EYDOLv1OkSKZMn0CMhxZnsBNkB6CtBUROGoeZN3G5F
0q95TvjFVxYpu3wJLguUS9X86IBxw7QRUsmkdZIEEV555ZNxgtSUTGk+YtytvuYj
/cSdeqwOKORVof3i/XV1FVgSFGpe5Vm09D9t9tKwsNE/+YNdlsBTQR7u8kpzxtk1
egZo3mfhOykZUJ2gDyONEwZxZiaQgtgzy4mo1M/mSGI4nz6bJv/Pe+iCeedlFfMZ
f6rUaf+1OmBlWrSlVZ9Oz36jY+g+N5mgIWqHJwAsgAEuKc3MBuHPhPXkhw1OTn5Z
AG3X6GtkfD1IIuvMa+VreUQ96p9cwui8rnrlmB5fwZy45+qJPmaMgGD/Q3dbGWt5
T4cMGz3LnkwgdAd0GzKZ1FV84Oeu0roL5eAUme6cWqEWoJMg9h2wR4u7GzsEHgAO
r/AsN/nKDU3h5JeUx5a+Vb2lzA6r6OTsbioCxewmcCMyNQGZ81bFgTzkcQv1yoO+
Gs+0Yg2LII1iHCODgIUinqK3j1kqlPAz18fxfKaOOLebZsbnF0DB1hPeS1NCxFE/
C9/s4g5ZNencK2AlRvH4JzhHnTOqr4u26wa8xClX0QQftzrjFkzUSIzvElLeB9lQ
5q0tmzgFE5pyoyjUo4ypG79AM7xWnaFsxgI/LgEVqxIBtjqkPUXOLUaA+uaD8Fzf
RR2exZBPT+T5lGpuMWnvzWARc6F/tTYpiFo3b+hGAzdefJ43+7Y2BbD7F/PWcQdY
9M7a8ZnEOXfTwcVlYf5eVYmvhmJOyRSiVWDr2/D4/hM862sJ+UB4UoI3qvNMcVjV
c8EZUfVaojxM5nT6L/s3tB1F39/BhnNrKTwYcqKutQ8dfCJn/kfA2/q8yxhnwBgB
HA9RFLRy5ZJUitkYLiGHJ7BZYBt/FhiPXMaqr72iYqvXvge9A04Lc35D0ps7Q0Zo
gNXV3am4kys2qg6Kg3eed0z5j+H0o9ZN1q7C7Te2vzynP92YxPE4KE8EpRTFx9nT
qIqJEqZP/AgCGcxJdvmHDzUpqWUSfvL4QUhs8GyJM1kN/xiU7BdKkjaXCIbkqv7v
jf2UVX3/LcWEEIsaBtWgYybjKtZfcfrUu/dv6r8SUoDFmr6b9aP2ea/xSC/Uyb1t
ieADTN5tfOAea2IEKEKc7Z5TdG1DtslXjQUa3PfMd2l3uJ8ix++lWmPAqyPAz2z9
UWExB/d9bBtbCfvShLqlVFRe4n4nlGZ9j1KnvJ5Bcx50O2Dt471mIxerdzFWHFBy
8Nx7vV9wZ8LlecY3SXErJ6Ffe5y9wh0Xd4A6IeAwwQS2uRg14DhXW/5UXSzQBcT9
PYqh6zMRytmEiOunRlFl8DPbe3RRD62vKcZx0zMH8wd2sVw3xkxAoaCDvT74X/ZV
Tcj0fvHb/ZKkV3f7+xxejxJuHzkjPUuWIUVUj70GWr8tXWa8BQ4L9Z1yMZT0i4fe
TiNt9OWtxl14TXKBWvEIgNb4pM6qTt0NGRQsa3aI3bRYyt7wVGiu/5UwQEUUSCF9
w3Ntjz48B9bPAt1vOKOta/4HXui+2IfGqYiqMMKCbQlAxsx2tnk/VKKMUq4R9ywP
ymcIN4HGJ1eH92zFiOKGgZv50sYoS1hiawHFWWQgYYoYmrOPPz7jlt3ikHsCvxeV
PLMr+tVc2wgMJKYxkS253CyQj3wf4M0trSb8wbiZphSIAGe5NqyAG20CKMsGNTx1
LLxuPOye0WWrPmJlY6QXJ9PgDXVT3pPrIfwlOYAe6SYRVRpyC1L0pzTzMTF6VYmU
VbOJL5gB3eu8Z7LcX/twIYnrb9vI99fYU2qL0wUUbptZgEN0M8tiv30BWco1M7vV
Cep5UAg8Drk9hgyNca8D0yR6Ucy2SbB45b3l+2ZSw69hx7V6lujEVNjZ1Iamt9Lk
OPwHxXymtV+UEIm+W7QISpGo4voerh6tpLNGNMUKkdjNfhc6jtBFtBScjs3OAWfj
hBk/JAaNo4ety+KwLGw2dOyUxcMPSi+qfoTZC3AvXTLycYdtXjjw+bcil4x7vPpL
mYbodEeIj/2n6f6WrdHUw9rwSWPLrFsyPY9YjlFzSwUS0bbroxJ2znkMNMsITGTC
1HqgepO4sRWWrO7wNZyJPiNzRNli/xsglrsHjYwXN/jlcMpHd5nAlLR3GaOQRawe
I/IORp5AJQfgQiggWNbgQRe7WpA3LHKQ96hEDjh5wFOxV5Egbxtz+iCR0ZjJUgoZ
/Mc3Yx69dITClOt43LCM6r2lgpksRdwO4f+Qj4TKtciviKXZfBKusX9ArChSZTua
eog+gBy3Fz/ptMyQVxffCs4ovXguT7qG4XWpErjYTPruuc0emYUFjOjY7PCcgfib
COYfHPF8bDIVL8974zi5AQrSlaSEUjIwSQvYm9tjFzfkInccFTe8czoyjsLlcXjd
8l5GjRQwIBRFbksS572F7AgeFO+cTlxQughFtrHOjlSrkEaS5uK5owo6rZYPqtCj
QD1cTlWUVcuGbB2CC4GiUGHANo1KKfZbLoXk7K+S9w5O0rEQW2oxTsOWRd11gm19
0bLiZEdBfhbgXVSi2+9a8APs5Lw6CzRe36ShTiuB9/JResmJ+GSnK+arobRQyvdL
U2Bl0nW4gVW9olxLdZKHnWDmZ3GhlBZLyyz23zUtLSgRIW3U+al4jZqFdao4zX8Y
QKb0vHaT8BLi0xFO3m9V4jeI22Wg7HB1NMAMMVanhCrxYlRz0Ze7m1rXD8wDPtfn
HOtuG2oH3kxq8SDY1j9xEKQa7os7Y1AkhBBJs3nMMmujNtSRuXucrv+A4p5SLaNR
6D/n9OzXNJKpejpR0HV9Cx3AZbbTxUCcLrachoMYssuThzsRmxdsF1kHEnmo2x5B
A9ReRN0EJnnriLCDmc8Gr3zd1xHP3brNLI8NNfBfRvAEPgSIf4MEOg0zqhDoeGe/
Q25djz1/8d741mwgwj0mX7kM7ay+OIHUo05pxRZk00VOZ8vmljZmS5u4WV4xxorp
o1JTNtE4VQDyoiFv7KodWVLBNcddWMXjy6DYg4l5a5xyVBdItxR5TS2vyPhkXspf
XlUy8ybRH2fyhUQfIVbip2e/suyGnNoQGph1fBO1ORhYrVG2BW5oWGbBSU7z8Jl7
vgAZhgBM8J1Qza19Ufg6nGh3t3pt9CLdTQRezcie3qI4Aq1rStr6E99sWUThHSUn
jPkn9qR+HN3+591X0sm9g17MOU05wALzZCvZnzjIuufuSNl0B0b8HRMyiBwZgBJE
Ms9xuWvNWjy0c6pFuisjoBDuLKps/rWoWR/YKuxulz2U+p6Xvk5DL216GF2T1Nrz
D5+ilNH/DKDRfOH0mP3sElQCMSh75pBf9MwXgj2grskPj1OOHnHoOwgnCEmYYp6o
dk/UA5aKBKo+VmIxGKJyS8kw5hZ9bx9KnutTLQDjcSVFBvPfBuy0yJnEoUZck9fX
GUFZ3UEIyztxebZG8e19xnOxnc8J6XNQjqwaD9YgFbLtuNlM4t3ccdWSeMrnTivf
a4uUlOfIcMQog0UP4pFL7w0PTCSZmmeCykYyK6CYDTDhCA9/3lV7OM3mw8kPlt+S
ZSyrZvvUzuv+8DdW6XF16WSD9iNI0AXmkb+F6FtQtpqoLMRKCLJnzndWxiS8X8Yg
2XlfbUxCfI6azPoSb6UIql60/r44QzQtKCOebgI5yiW9BWgMtersPbZqH6Wvvtoq
KT3cBlWfMdv6v6hYUD7oUy2JbXewFt9Sj1rXdMZm6wBbhdfaHWKMKV6SaxxUKolw
q7HfRtwBwFr/J2/Sid0oud7vRjeSDeQk+1Gp066cn8FyOxNee1+6sicNVeWpoI4T
CxErZG27h+t7xbt1+YFWS0nn9ccmOkeD2qW03CTHJXnz3lbqn9qVFaXcZv/YE87i
DMCpa2uEVQ5rYLdpAa1KG7IdIntdZfLPNToid9pfjXnRhZUrA75hYO7kHcGFDbqD
eaOnRnyVhiKnosq9O+WXVqdzJw/bKpyGlFUoTyI8U39afdzkqNsC3u+82LNdZbr8
63zixKkELVIcHhnhJbwXh1A7fxNm2mZBtljPdErsnYqIeFYaH7J/ZuazVIzzptxy
GzRZX42WNj/BzX39QzFjwI/vQv7vwrSxIkKM3oilqVe1bpnYfl710TDdQKFlXyB9
P/qAApqOxwDtHsjXOSbIzDahCiRySQx9p0P3ZiUMVLIw2NJe/OImsaseryMvfcB+
tYb54m+8McV9lDDT0Et6orI9KuyqxfR9yJ9u1Zr9rA/PvGGJJ1KDb9ZgAZSar9Kh
5cYt47Vz6BcCLm13E/aGAbtEVKR7vxerGd8Qn1LSbW8huGusVVeXNTp8VoaFutWu
esfslm3L4LLGZ2sksiG3vrcHg2pSZwD6QyHL60AK3SBydCsw/csF+c2JFkGuD9uh
TRZTb5A5+4J5Gs7Wh1GFH6AckPm1zRG9BCiA9Tp7c4EfzlUECAFluA1C69KZ30YS
epMdAhbCmhDL6WelOnyI+QomFQ025LIBpz2C1C8PQrVlwZVrCntq8PuqfSE0s49K
tmXnvqA04R6FNFoCSO1NAloDk6+Rp3ccYZcvWNJvxFrJtD4om+x4wM93ddMgz6Qz
Q0bqW3dWfRV73V0B1ya0cx3tDkQcUgXzVQaTQ7Pg6FSOdjbnLrfHSGWfRFVtbWrM
gl6HbB4lmuXuaK0VrFm+r/VPpc6KObcW/nfWCrcTey32G/7L8RV+gQ2PYkHNQaZj
P+oOGfNxyk7I/AoH8m4No8JUwuyVL+DwIWV21AuVK9lbDqak2tOwyBZ6UZd4JaG/
HGdc8+p1nKciZUotZENZzSs4GOmUkD7oUXNwO0dHkU5bUrU1tooybgtzVeLwN4OE
kgJHPNOw3VBoWSWrSzu3yeq0cWgGt+nenjlzLlCUyqFWfU155Q+pPnn1lDntSAIA
OHcPT5KBpqPSf3RmVORKAfWw06S/hJ92fSVaDCynbe4Ls2g0Kio+BBlTg68/I86J
VQay+rF67pjcx95um3E9MRlYwxYvzWk2FLfGxERydBUKzZYqMy5wWxgoXliN42t7
dTm20Vuozt84lyAeVjNhD1Ndb1+b3XbJ+LuuMw8ibcM3FHaWD4qlywIYewy4o8Cb
EzUvaEvoji4/tnlYMyJzpp05jkRNiP4kbacsrTnjVRxN1s9EAkeMB6lZfoke3QAy
enpd3gBMMdIyp/kSO6JWB9p+BgwiRp55M1uCdBmwABNWx3+iyVwXa/EfYt3UkmKU
FyI0X6x/pb/oZx+XcP22SGJVcpqK9LIeDnt/H+sD2qVUKaHMQ5plYGM+tjSjqqxU
ig46IAeSdRefd/OgSIgaDOS6FcS4v9aAk4QVqtNsO17QokdHmlzH/myEvkSr+mQA
jZmvh+AcC3VxxGx6JCXntxyKy/LEKGzVn1/7jZSLrI41wu8xF3UgwE4jz48vKKN3
69v8ID97r9rKP+QseIr/CSQ4Z2CKMTZaSq3tj7JJVTvgSK8Oqwz7kDamchOV5I2Y
uG9Ktlm/A1ef84eB8+ZCGmplFFPjGS3x7ThU2QnyHyHmEmqDBoYemRuqFgmTCFzT
dbFKteb/cHz7jiwbtU5WuR8/HgUZSi0XutrTljsmqtwYo/4Ie86DkeC0w1oSikEB
ibDBKuyiUtEigtpkdZofSy+cYkTHrLu4ff3yDkfF9dELE4Y6agiuOqAvSEycX4En
/jAVPKg1vbZdPSUFe0y11aZeCnjjkh/GJ1AbOL7eJJH6Q2LmCt7FgKwBZZNh4GyR
CJFGsPFdLAa2aGX2UoP/4DvbjblHSltPLRbml4TeRDzdnNpbSZwZ10ixSB6+ns7b
DEFImNfvJmJwgcoGaRwtsF+fX2iR4j9+RaG6D8/e4N65uoTMd8xlZFeCATJwOWPt
IcKiCUCC7o8ldQ73FmU1hhF2EnWdLY5Jvj2/EPwoCBjffPBhcdsqusSR2mjSBEK4
DBG+Y/AFYBnjlhkDYL7S8CeeQ/cU/Mm8ja0jSRK5yBeDGOt7oTJIBC6pQQvYsvL7
zl8kuK5ScBxXN9YY1LgsDh1DrYpOcExBxVnPoRgpN1YEq0kJJ3/pk7ApYYbjWo4I
Uwul/baWdoPXwCnrrLuzyBoT36m1COwlhVqPqprSNtmUj3KzpRUJlTP2tXPGdU0y
X8RdOkm3RV7rr8RUOW63Y/hNEz5MlyacHa4+/SUfCAJcywQ5qE6k/Cr5bSKObDt6
ZRBTQJFObrzl/H5jAurQ8/Mxc6XhrRZu2YoZY9yaZlBc9uR+IkvWLJlMGRwEcOrZ
iBIb2w1v9EZm8kWqVjBalniZ12BRciuasqb1Y5LkhriIHxuTPRdJ75yfxmAalLDU
OGR5KS1Uja/WJma9O+t4IqYpn72LAy5RHvWtkVoNrdOCx8VWx6WxSqR2I94NyKLd
EvoJtg5n5/CDGMy8BhsPqQJi6NiOn1MCmwR2HInTb2tCDQIJ3FR10PhpJ+bIuKuv
fUMBKBZC3LubpUFaEhDjHVQdeUBtRZxkZudGXJJru2cHbV8lvYx/XQ1w+wTpBr3X
qHCajIS9qvejj5r3FabKNBYBwmR13h8c71Y5YI8IpK0iRgYGJdJGb72T/l3FCA0q
gaaHikgqjxG5tXS3/5yIELa4sAqtw1BN656GZiyhUb9SJwjqci9GeHMOVuB6TlOX
UoOCQwnWSVy3g8PDQyYJ/2OHwml1Q2xQZOqKDmC/pl2GU5HJA0knehfUop70S80/
RLcBDeiMQWWd3/5EVGUnR10VGi8d8WEeINhBtjR/hu2yB/hblVE+m3Nw5GeEsaQW
7DWEndUi/dRkaoecLlUIDDrypv+DWf6kphmhIG2qm1xdNdtFE89ZZb1ByKgpi0DJ
4ETnG5/7Yjs+GJSaH4t2aiSDagb78iM3sNf/GsEwdX0N5kvKpNcHnQFAl0IT/Vdy
0IRf9/uWh9AdNeI3CBn5PVfxjHl1i3CRaHH0pZnuyfZP76cuxjH9HnqcniFiJpsJ
r5p2uhfuppemUisbeSp/H3nrI6QIOPWEomBtnXnDb2YJdFz+hbRJg7E8giOOhtUO
hOlkLq8KoaVZzxU/PMoDWSW0QVxetPDevMaMZ7uA8/cf/TyRAnr0mXhRbDFykDJO
PnrXc3EoF8qN4xvlVogM5rI/zVjGXH4sZ9tLRQrq6qqVoZZxkHj3GDfc6GmpBGTg
Y08cu4Ul87y2849sZdFvgqEiv952EDfj2x9gIHjtWUj4yeVi1emBK0CXEZNj0VM8
t1HDt1024NSSoy/hRXO1ljEutZvTZoht1gbnTBiiMD2HW00pVh8Vq1+EIbNfnXSy
r6+zqgPnDrkEoVU07ly+3dcJLUVhqA6B5AldIpz/1GZblcfb1e85yvr0fOCApvV+
9MhVLaGcj064bLF+jdjaly3s2m9+z1f7XJomSXCpUOrHayblrds8eaf7cpTkZOWh
hDprLpaSUl4y+ZxCA4y5RGTO0ILm9732znDocL36rYqkwD4X3VTERJEUYpdph4rd
NkgqsZaVzZ28zLDetWX8sjKGFmEphKW2WpICXhNlpE6btQarupazpyJF1VpX0bZj
VKUqUEW3Vti8KaISA+fUnprGq/+0hhgVknZaG1xUUqKGh+2laj2+yt6rls7CB6pA
FytxR2uDryj5CKI4NDCVjMvAV8nR4brUWBWLl+C/jSYH8znV5o/fTIQGUY2qPX4+
kdpKMpQduCb/Jpnl3TJPZI2prPySgVNo9ubCVzNEfRvyAXFpvpHqyLiEt3GVBH5Z
opxi+s1b1Of9vjRmTc7yApsowQnJVqxRRmhsD/WfaC2C3oM6hh9MxUWqXCvUES3x
V6l6HtHhYLeAzMApRxD0rw8AE9d5EzIGmmPL++HN44V001YeYlgs9oVCYoIZMKjo
iTbAEooqC7O2Duo39O7LZRagrtQBOyXJ6Zyg0vPQMLBObdUAFB6d1dtELB5byp5S
lt1P0gbB17wT6IOUY5gNAz/0IMYWeD6RGA1//PXJKvyowJaOjp3aGpNIMIuugzZI
8MQ3po2l74oxMNqGq5/AL5lpDzW5C3++6pWiZi6Hi3Sp/0vN9meb8DQjjru0B8Ty
6e2xqlgll7d1BjKIo/zIYxH2GExNAF9x98V15hf/3QIVQ6oa6W16VrmZc7wPrM/o
oJ5hLkz9QpB+PXA1NQTjGuwrm1UeeznOiEnRTkHqGZFh1imY9UuPLpeFf81NzutN
ZjMvnPljRZVF6QsLXp00ydxGSunqN+kqWcI+5yuLUhU1tvSsIMREcvlekZgA+8z9
iMw5+AnopPHwApilj9KoBpWhNpsenLmXKZsrrFWZuMVXDxU0sZZoS/vmZTPpQkhj
kGETFWey8LuGvicRDIApWeFPokGn7TDbaWEFyzz5vGFGpGDNyGKVX0UNzvOG/1nH
Fo0yxDVM6eYaI63M5rN9UjdxZYkMPhghAxYHfxIMKwilXQ9mgQMY9ftwFsFEJN/f
pMTTW73l94rWoUTFBwI9WDz8vVS3Gakqpcl2M/vuw4qljD1fQ5drUQyuQllx8b8N
W6BFkCY4ABbon8uFPKQr06nFslbFSFcVP7FGgbBdCIPg4qVG92ND7LSsCuJF2Iir
e7MlcrzImqcfNLAPHlGVVuNCPhF4up1F4/20D3kuPABpXvrEVuOwJQlQuU7VeCX/
B6ZWhAKNPPOZjb6zgMOYEldv8PwrGDlVxsD2UrX8+SNWG1XPjCY8c7YwERWNE1IW
rr5a5rgcvKR9KKzpZnPT3r6Lp5FZHGC2XXXiHGk2qP8STUpepcP+llacKNMZfpTO
dLHB1VELdWcR/WjdEdtXKkZne5LTlFxAP/X/lRagJ/xm+DnWY6WvCF+kk3PpuMfU
ZPwxrWsnDvqgpqx9vTT6R3xnd+dTv/EkI+8U6S+6zFlYEDrWXyrREApCztCUlpk4
ca1rJICVMId4arjSQLKfgohxfKP0UPuAFsUiL4Ak4K5kcyr4RNmRi9bSWXBH03Zo
aBXkHBkp9sRAigVQL5l/DB/paf8dPX6VTNL2+NuolYq4hEVd3n5ePrTbhsUE2L1b
HZKVugdLyTYiFMdOiprw4hxnd/ECH2QKoO0xbP+HT8Uu5GmHoQxuMKJ7q//AXHMU
rrsNtS4mr09emcIaFUPwKSp2NWHXJ0IpgoyZWmxhBsLEX+RXl0KNZ8KrcAM7q2dw
9AVI+yuf6wpebIvkM+kYStY3G+23eL9SrMAVAwzlH0v49YSo0d+ZQLcO6ts3xhvX
E7RTS6qiD9H1g81MrR9kpZd4/OBHA6uqFMZpCRsiHl4bsj+De4ZTjAN2gO94ImOa
Wsjby+QvM6556JUGENCFZfQwQcCBoRSqcukkqMsLt9HOrE2uOqF9eLhZLiymv7vs
PPwV4SptxfuQYNgepdUt/H37HBIwYopX+cRPkqXaVdaq+W4+/JwW3KOd41ACJp1S
B7k9WOn487f/XC7GXYb+wGCK97MucOF9Tul4gG+anMHAAB9uIykP78hcWqEmRKdh
oCrIiSO6zDusk6b7K9938E0hcaMIdohtscGoVXVnt+wB4gJyDrAt8a/PA8xcs3kJ
VkYh3phnBSvHP9iBfbcH6xP8a282XEyCKWJOGwtuDrmri5NxdGL9cwqfOgKE1/Kh
R5IHN50CQKy5PS+IZv9CgJ7HjmwSz0J8T0kLkSig4uBhlXLTDqYuPCKYT+A7/fpQ
TfYi3N/BC31ToewGIEwXstRYet2qySoGEXTjvys4FlXpO488KWhsbiAvhhOrHxdl
N3GmektJFQ31wsk7bzIuUkrbBxoAsmnRZXU+PEyeKU7lY0RU1bldoIzgO63AafiT
IIZnbp9t+8GiU42zioXqTexD3gTgXX2COHCF96PuLvf0kbNJwjSw4bpPTwVzLEYb
AydRUAc/2JF9TXnOdcO8AEWbXcN4nr2vtuy7TfKryUYMFWXpCeLL1I6lMtzNq6oy
KjP/yUbWL3sA/+l6bMK71Z2CbqthlmQVT00mSwSSuEsd4BEDpWxTKWY8eGPDCXQg
MFZ7oc9/69hZ75/ny//jpGiO8AYrkURBsJVZ2mBUxC0YWWRXF/hbo5KnFAAzNocK
wzO9Pu9bUgRVh8gdb42ulUhZ2k/Unu2S4u9zRY9lwwKaHPB5j2C66Yk6bXpla5nX
5DL7b0D4jZqFVVuYXlKjWODRCcdveAPAsW4BgjPhHTMxSwbKnBx3/1IZDLSyzCpF
0+2v5bLPoFlyWwtwe/Qqu7E072FZPy9AnTh8LNVkhNfSFZlFFu2VfveJJBlKMLix
jylw6JsA1D7MFrsURR6nS79ug7aiiZY7BZBEhhLCBQDWKzU9iCwHiGfhCma5vRVk
7mYEVHUYNbsB6tt+rSoF1lJ+xFAEnKzeEGrt72AhU3w6bGGQ81UrOawyWs50Lz9M
XvauroXz2SCHhngvZETLgSR50tABLDYTX7fy3a8fowVdgoy4KPSVZwJCsPQ9aOll
PshzxUHeJYMe0wVjkqYZ4WAfFChHTCwieBaeDmdMXGCEnVBoYp8xkbbaksmA2Bsj
NCJQ5JTRDr0gu8KetrC7u8kO54Iyn08ejkHqKe9fZWCRxqEBCOUEJVK33BjRY4Z3
bctNKD0OuLyNFmzNk5ho+PsiCpAr7qoItDAUDM4TK7S7EqzfaEwg08v9JjVDt1Wo
HXkszQjHhfLhAQnrvU04SVKrAoFetQcNuhAND5kF5tJWQfrPqDyRbdPT/MUXVRia
vEOBgJQhS8jDbdpaVEFtB4Ztrosw4E/k9UO8BdlOnjoxGYlb5vWXK2uHsz0ESGow
b2rLt/J91lj1ASAtpHfCbaAb2rRYyp3oZAXPchPbItB3Bl4Ho9GIDib6KWCi2qap
Q0KsHH8KjU0kiY5+tTxKdAmCpEmCFpeLYcbHJd47hgTIcJSiDO4FpJHSQChz+10P
iN/tDXRuKOdJlagfxBIPxRQpOLxjr+FThf6FJwk3FS1lFou5h72GWY85b3CyWFGu
mPImw7/1vcJR3/c/I21uKUhuckSzVv7AtrCOQoaPWc+lv3dxdVBzsbdPliNih7It
f+4TDx0JElXCg85HRfQ2oRimv9ZM0O2Ysel83ZrB44QC164yXCf/3qT/M4M9Ch9S
1qcYaAdGN7AXJELpaDF9Pi8f2sJt7XrHFwcYYvR4VOcXP2aZf3OrsxWEklllONrJ
B4n/sAKULJ6dh9Dj6iTPDU0YV4lvW9FBgQImNCklYRwBq16ywu0ehCQ1KEfurYLJ
XsmM+cQz2jGlZkCE83ThN8G+m7ubZPIrVR3b7N+n/64tZxLglgOU1+R9Ua4QPI8G
k7USib57UMkQO+bsfkAvoODNq9aogcO64lcDDtvk0CBzDYh1Vbj91tkIEKk+FvOa
JioWtcvtJID0WVTpHyxgU40JnnYkpRd2PycbospSt/i4FH0YzBHXlIPP06IedrCb
rbSrnAJ77Po+wGpcQwoQ+AOWkCdQR+rvQZGVqzWD36NGeuzdam8N+DwCIzTTWJ+h
b0hBMeT0ix8UalX1RDeMmPF44BPvXu4D9iJVHqD2mm53gg8swHNcwCdp+mLqy++y
n4EjkyeWHCT9HiK6O2ThQhT+9kT3v14pZvlwTj1ilDQt6vM8lpNee0gc5+8QEKqz
afw3odB6gE+8GyQ+GOavs0Im/LldzQxoR4N0wSAE296pIh+I0cKMKM/KOGA0fbOz
qGyAJan6KDhgKvX4aH8KYm60jJKa1FgbiUm9o+hL5IVpeWYJo5KfHNd6iKbFhZWw
afcwaXt8HtnxzetTBqqkdwmUPwMBiaJW7KlYQAz6BuZc2hcF3vkeQwInQhe0N+Gz
YGEMReF2+/ndzDtia3h00EzfXIBqZ0m3cSSG/YRYFrR0GtjvTKtZIuQ3OI87ifui
Rd1C32sw3ufbBzA0zkaKrzjEJsPh00nA2wYBFYL6kTMdk4uZse0rL3PJ9s4XkpFj
0VyTTrpIo251xNKjZxNhobdr+hkST8o2W4fIezBnXzFK0ERoLJAxSbJhmGrZ7k+C
ycLu+M5ECWqEuRG1Q4rWo7RbT2+DKurIrm4LQCBOtSEQGnzCY+NqgWU4ailGZ/Lh
K+B6Nhr3vUetMlLDuJzphnKp9zZcuZibZqe7WMyWxXP3pk2454GHpfEz8JWL9HiX
LydM5EZ0YRGkfdC+bIfCWYi9jUbMUZoRYr+SYfGGLzMdcRP58FLjA0zwHwPyEczn
D2E4CqqzCNiOHQbMixwwmucl1RybbfbK2CpVIYsYD2szACE9yexwH5YS4Me8rR5g
BOt8rV7ha75lEU1kGZ8McrKiOpEp6QJdh176qlN++UhcJPMqUVg6dGFEuHLx/i/f
2b9ralvoj2ln4i4JqVBYhIRSbY7WWxVXSiPG9oHFLQos1ePKwkcjofT0dxypudxG
+ENCJaApaaTVEAKUn2lhEiPgWrOnulz6iS9qlBm2F6VMGd9Xdjbw1+Psk9GVm8+d
8dWtNGNICcw6Svd0viTWj1CGnEFLSoXwBLkD900l0BnCM2zPV7qsZ1Mb+iJ8NpmX
Z/39vzmHkwyYJxzEI0kLr/akCgbA7kjxTlMrL8TxL/jXen7W+ZozCNQBnOUDylQt
ImjLf3WdIuZxk/t6D/DKTAPyYq/ZV+oegP3/6ZRtNgmgWnYEk5aLxOmU5VwHURW5
o709JNCRAks7Gie3UlyyClM66afhZgfs+lVZTazpfYZ6+RKah8WagXJwULsaYkvu
xRwFrNLdSY2Dh4+wXhnLnUUmz3NdfpCekuaYELfB6fCDmce8mWjWOZGdzjINBn7a
+/EHPSz6MY58pmOUBqIw7mAZDT5DnX9EJBUzA1y0SIf8LdzVU1eECLMfvMEz+Jyk
hx4qILO4XuBRI7o4YGeYBpplg/QMtlia79HW2TeNk1lKEdix7VVNT8MD7kz//uAE
rqQDq5A6bZyCd70M+aoTj5lq4jxWUt7An+eyZNcSEB2q3w+x1bNLg/97JaF5/4kK
WR6YOmfYQIFQYZFdsUMvmlMvXg42AD1qMsrqm2VkJSZOAfW6GI7pgTYjN3HD9O2M
ABRnxcyeyNemW3K8ocpbvjq0+I17A2HuvQEvJUq7+hegfMy3k0IbdTbMq6xoskEj
XXEvNGaf6ZFu+ehr5yv6Q1QrOf9sO858pyVNYgCRQZnKOyO9wMWVDwQak5lDwmST
ES0jG+NpIPkkdlTNWBWz3DBtyD1igKMur9c7LNTRF1pEgWNikmWbzf+KLiam4oKk
tMrbh/3AJDOVrZ/DFhX3xIKYq6Yq66BqDsRVqQYnDn/YghXZIs6x3VirPuS84xic
wJ9GYc6MYWMPyoZH1zrOGQLtAV1WKoMW7ETBRG4JiEtJCzjp6SfYXF/LUc7LOWkv
KM/xp7SRiyPaF0+cBCUTC/tKbjcEpljiTSoZpVAEwbTSFqShZN/2saw52tGSaWl+
o7gZx0dzNJc8mLIkW3LEIvrjvCLiJQcfMHexMCa2ULShO1Hfmh4J/WXWfYroS1m+
LgzGrpPmKyPSbbucIeM56q1BG8WdYruEtl1FZjHuxAFl1NhhL1Zm2Y3psky0PxTp
1g9Po458HdueyzPhlpYDHnyZoveZkjI+3uNXhhQRex/xVYPzHRlewHGWiapn0xwN
rFfyZUsrZnrrW+/6gS8s7zaQ0JyRe3s04edZrkZlTC1MdWu0hGJiaify0Ofha6zA
H0TJtNAcCtF9pmK8a/ZUVtAISYla8qFIg3wReXo82NNE0nYPp0cyWTXo0NiGSZpH
7ekUIu40CXJpcJ6b1ia89ooQyqSUUgaBK1aurUk9ImYZkeC1iis0lI8vzW3UTdEK
iHpECBtyjvDp9Jhj7qHqUKsUchVXffvt5pUY7Tye5KpBabLhdUQOCjHmkIRlzOLl
CbwqSg39XzrV5YOn5xtGM3QPE8l3yqcdoWDNtXm+3BvtLSVZ+1xrHXkvgHQkwFiK
oj4NXlXiemM5vGe9RT2mzLmf00BuakDzvtM1MAnJieeZATvJMondHkhvRQ+gt0sN
FD56QPReCdfRV6AvnPRPhJDNm1avGJeOTeixXCAcQgbXOvYgfjsAadLESyCO8W7O
dOegbCWW9eHqMX4JMNF9hGl7v4TJksvnKgtyCypQhiaGYKtlYo6NJqKXngFcy4C0
fdX7BO0kt93igr+ydSvNp4Fke4bGt1SSA5yi3lVrJCShritpeqbojgohNrjec50J
rfAs/g0ktmFAJojkIi9HoUPQFx5iMy3tSJ97Uy7bBq7W6mthd6AMZa7DZBvuCkdI
Qwf4WVpLD2rAVztADS7BQqtSpgvB3OAlWtQKfrbyEbrG8I7n/b+3oD86FSHAPluh
iIcaHnWD38JC3EShGkTWRcOK4KyQUQzNvii4IhvBsgDSBxnoFFabtwwRoAh0sLNg
Y6fvC1RiLb5+nSw7cK9YQr99w1GxK4a55fANz0A2opPBKLCnDRMWoMGR6O5zEG1q
DgYRZ9AjXVodYiTuKgkknSUHfoOWw1xXpzAtqyPFjxAnfQeB+ERqAI1PTDbpoofT
JLylva+FwJOplw2XpFt/USii37tnnl+WduNaaUdAPwpNpZzky0wX7fA5IndCxNOo
lNkCOhv4eEl8TitulWA7uuRJY95SwZtOSDn9opOWuaJs+zTmQfMNZ6znpzMTX1pj
8ndcBWFVVkFoI8jm2XkLFAQq/eGXhEoZ/Lyca1GbVpVSn5TfW2wNBnvQSO63+5dv
UQq1ATx99/NLecJ5/5H4n7A27i6+3i1oJPotAXdpV/W/nes8cGxj2fzlAYJk7T2j
rYtOdp4/HfStf4tTsviZx3HLoHm28HJYX4PsnynY30Fr0OeJfFFfC8VksieY6Yw/
J7Iyt+7ytW7BTrbJuctVFvzpgFc34Wcfk5OhlkWd2sdtyBCHUtSy4CQzBTNHKqkC
lHfdJg7X9HFj3evt0xREZjyn+/17IrcmfPwV2WFTIRPrvVJdHPQ5WybYSUjKO/HW
m6gga1HnCDPnEBAtjnwr4KUm8uw9Cw5NYDzVlPtfrtjChgNU+n1a2ne1vxDoiH/8
Yr1lJ/N236gelTE9tXAsx4iKGPVXXfepehkSoQ9JWTA6nya89bH1r4qKsNXnichb
ZbgE5o4/SLccD1Vt2F53ADl7YkUIZ/HrbuZ8SAvbOLJ2jelFb/S7bXsNwbG9EU2m
VfLH+XOpB5NuNb//JfzXTipPM5C/3MkIn5XqVLyVadc21cT4UaXJiYTrYOJzNMs9
3/qnWKNHQH9nYohDNY0rtr1KRs3qv4Lcya6QBx2eMrQYyadrda/Unq0ORvKSWHnc
lEUj1C7S52DJmywE5xlkpwfkuOitRF4G6f5uWDx4d9O46pF8IDQaNNJaqIkgbBc4
53V4HDOKBhnusDkxJOS2e30iFmrJzVHmooJzDfSD/ICrsPGwe6NNAcv8Xs83voDz
yIOQ0aSX0iXEYU//qMXVaJjKUpartzPGE2ZOupKzE6yvNUeSsrwLJUUhbs+J1qzP
IfL39anBgJFg234EB9fUJqbivCZ9Rt6K1bMFMo92qpu3FaMRyf6Jkn3UltMMtIl4
+UUC1Cnj0xvQ7lGYAFcHH8GlHb+CQHi8zvSHJf0kDytWH4KHWMGnHuHlQYrohdbj
l/Dmqo6xhZ3wpdz1LjBZ2MeuSZ6wq7w4H75dX4C8ELmLTrlVqHY1Rz3VA4GC1Oto
YU30gKVdWDmoW60Jg+OOpxHTp5qAcVPfQ2dT2dWQLKZFjnjWeWUrPJJ1bxh4yoQQ
absI7wEkmwNKhKCawgyvKXRL9uOJF3RiLi4jFRuKQvhrfnrIyctiz5ggNT+QIFMU
wY8MrE2WNSpTfbfogSziKmVj4j1sSSBB+lTBAUJYwA58MzyUPuyjrwEQm3rsDmrW
67WhG0x9583OTZaSDlD5KaRpO7t5Omz8kNBDr9yU6OLdGIh4FmkAAYT0MOnx7hoX
DNlT1mRnKdZpvExP7CbS6c0K2jpo6ggmn/cUNtJiejzBEHPpUvTPMVuidfual5Mr
rlkc/IWn81EqeQWQEHjtqJcTi8LzBNlYnqUdX5JfHi59TBGuS2o9BhCwKKRrgNsa
L44jYu/ko1sF/K7W0hhdl5wVO7k6QpTJg41E28fwj/HVGUXIFUvmnIgla2Cq75C5
GilViYwfKBVIabpF4pOLCn4/MfxA9VX5Gxn37CVd3lvHKFVRR3QzJSytTAHt6EAM
nWRwtiyS2Z2YoI1oW8BTArCYkst/2XFToSjlA0raQob62c/ofuZwFKGi4dx3cdx8
rR3uyIupBOMB7rJYVVn13ZiDmS3DS688lLY1jIdIcIVwsKCn92WyTNqeVbuamP1I
CKAzQd5tm5KHzFsTBaiI04JIJckU3N9AQgbhZl6sKOfjLjlcd516tQVfCI8n+Yy9
icfjHrkHAQk2uxZm1LN97zzf9sBGIO2mPK7Z1nzJd9CZZQL2HaiAbbsmnSGFIpFK
MUCNN40h8YP9zYwoxNLbyN3PihHJSP8ksFRxLMBEdNGQdhHqS+3Z2Adocps/D+hR
4qnYd6jG8gWo3OTDD5DqQjyM5HokzUlKohxFVkYH1wD/lCMCsjeT4WIwMCNpGqaY
NXFkzDFSH1NWhURJjixkkUwEb0ZRnmNF3Ya0FLz87RAFV1tyMj1l3JdEvHtAQfCC
piGtKbbZG62yJq9NOxYjnSSrtQRp8uewHQbtmb82v84X4dCv+z8n27xIydyeH61E
m514SH6aY82dHHRYgV7JMcJA107QbO5PprKPF7Jl3Uue3jIsv8fRRj2eOLDYLq1q
IskQrcdXNlhepVTXSdXYUBwUfC64OAUI9BTExakYLphkA73TEVfE/Vcq+ps7dMiZ
bX9j2YQDUUfwqtradKgwL6aLE22JASarxbLRWOhjYb08X/BgzVxgKK/cmlXUDEok
swSlHAxzxVEh8fQ8lx1Qr05x+BmceC2YpxMwSnL5nIwahKASyy28qz47AMVs9500
d3uqFWZtDDCNIqR9GXCbKKxYpIMYxH9WmR9FU4YzqTxtnkyZa/FIhNgI6t+6yQHK
wE6YUMRKZl0khqQgb5w3vIXTpH3E6vT6xrm2xM7ldq6hASQS0i6oG7zgnaFNHUHs
4WW5gQ/Z+tyuTp2ChQdQ0e4ONJGagkpvRRM4iMqEiVc8DxXeKGs4nV+IglQYzHIe
jLU52EcxWKlpVQmWwKThMPKe7wwVTCrTLT3WuZ0qgMQu8xkudpgESzspsUKWP7+q
6viGKjuOtobcTzq2rArz7Vb5iyVyfGzV888wXWpxXC7fIM7NM7gz617s7dpN86kc
405mTTHVNczXvtykiDq3o1LLy7omdpd9Zv9OovMMJzjSPw7TuZQamOaB1KPXuHOZ
mmLQr8qjasn0bWrULiC1GyVdrYGhZu1hcujHk/pwgfwMPlho/Kr6R+B99Aszqd/X
/dTb2+j9SVuXrZwnYXXA0TSA2hBtYNvolwc7rM1laf8OmYlAVOsv71a8m9JB3iJI
UmMuYfgO9fcvsH+MO4yeynYLbMdJLe3Lx40m1dXs3r6eeP2EbHNVDQpomNJixwu9
V/Cvt7w28Md4j9uHlpJATKo9CSYKCTP6NX6UT2vywIbfToe5Gya+uSPPZKYt9eud
o3shlaNcghSn1qEOy3W3ZefaLe3JlCNhupBxFh4OrUznP7R2/T0F3xJ475tTeYjp
TIuUEEKIAFt0Red3JJgjEwqMHMj3MpVVCSiWl/+CvNSTZrzPMMnZAcglupAjPgJx
CHkuSByfgSme1Mp55jWqo9GI2eQUEhxZWLh/JQy+satf/be06ZzHTFBwc8MJVcOQ
ZBolc6vYkkf8wIS/ymu/7tAQKm7RCdjqeE4waKwesQcP7dV9QiwxtD77dcZNtf3s
RV9Hbqya9+jGMCXjbA0pkd+opHYEzMjn0dRRuHW7I5gr99Ldc9oO++zWyNiiyWTe
8X6NOMmiqR722ZdYewLsSV/woO6ilSeMCl/v/iEQFYkHWoQWZM2q05R0URGimfGG
eUzIN3lFsC4uxu80X5PUbMtfXKvzcyQCe6kTuUF5HzdKJgju92o3LAWVw6BQms1+
l+n+noLjq6IRYkz9zKG9VZdEbTpk5E+isonPV5/Nwg7TmnQDNYNn97+t8u5I+dFa
NXaiDijNVuRxLU5vdzAEOm4s4+IlK04fcYPQt3ri4HjFkhHPXMQV3BPS59c23A0v
e1EeKX1KnmYVWEZimDZ6uXwrjAPd7dK0UHr7FNeMpwWs35kXD9IAamFCxW9QiHGM
NmqJG0vFny9U+wubHuZtZUqh1SweRCX6+6k2VRIYbqouBP+HEUYVCZwEncmqCFH6
JRRAgrVqPfqEB7DeUcmhAUofxGbrw173JJZcjMa33C9wanWM0ePoSOQsffAC2jWy
zaEvBP0g1le1yK6NoNrZZ3KVOEGN5t4k1GSAkiat6c04NZkFjsbj9T0ck0yxGVqM
rpMTV4KaqxnJUo/Oq7Rd91bSvmrJWvqcpbCeV1LkF3GBvRB/5yJeoy8ceXLZtDbB
tZD646HtnzgPoDsrbdQm/tMMExhClVpW2JuWK3L/5EWUTmLjAgMcDJF+jnO3Ipwz
JbRcov0D+P/AsKII4p3OrJhtI44Z7aqmCeVabS9NAKqxAmzXKStVGX6u3pyH84D0
0zcIfYAYsbXFQ9MaCsOujIH5rkaKPifpL6FL+Xgsrbb3iH9psVaWhOQCbWiWWmYg
hPxIo+xLyJl/bPSFMWTZ3zF9KhfsSPBDW162NZnGdb+et2htA+3GmBrWwP2sKbPp
Qyow55mx7VDhLtHYFms1pjWaNapZbXh3yZNlDns5h9ivsxaSUkhMySKXXKZHk2L7
AMGnL8MQwL1uizhyDtSoXUcts2qu1B/nY1iauUDJ8qVGnuzzNJdNYW+D0OnoPXcA
qKteigQFE/ZtFEYk+gfG+AzSS0/SRU9VoBUc5dPJyXRdJsExkKLOLjERScqG131h
PXmPdeB1mNzy4Lpvw9vDnkyM+536wBItR0tOh7cVNIdi+o7mqn4J4Y1nuw6I+DE1
JiwzqFgHTbJNdQ1eInTGlpAZeLo1qWwiDZ18VIeqoNMiQxhTtT6vf9QNnTaMtD2m
0iqK2RVRt4n2JL96mPJjAzrHkIPKN/DMjbMwjTggYSSjPa0BlVT/hISkm3YR30sj
oDHbkvqd+iTqRTz62/khqrpNJQioXtcrWdUIi6CADpCo1PIM4iL5JyeVVWvFQVjF
ktasv6OD7V+DWg3TdwdTwGazt5YRgh7rrQOlnZQnG+bwgmDGPUpUayT6VHCZn+xh
CAgNAbW6DaR4susc5wkztE81YnO5YPv5P7mrKmIqFIKSLtHxlGdUl2b0f2/grUXI
bb2wzTPrXmIjAUojJrdjnkgPzouWD0jv9PxaxJLRGgcr9GsywxQ5yP4ULWAXeHcJ
YIf+QeKpqRvlFPBjBUEeSYUgT58yzqZuqm89Ka6VecmXkaR1Tuhpd+szI1w5koOP
ARt/wyeLIZIs5S0gOGfRVGGKbEjr4LImUplaMdiZyYQjjNUu/wLmfP2IKCC6uNjs
w9tyia00XQZizUG3BGirxbh4I+HjwNRYQRN2nWN6GpWiZXDSmUjHVaDzVcHJeT+O
BKXeXlrGTZp9BMBsHUR+iyFCbpq5BMrEqH/uGrLllCo39nwuCUXaeRMORK2GstV/
hWte3P9NlLGD1s8tB4FGv0KjlYBlvce1u+trrTBVxNlaS+n0nqzUxElvR+czKUWs
X9v8z74h68LF2RtJ7DWTk/J0NrJ7cmU8DZ3zKx+wWmKD/fsNWDXQYpFbCi5q/UlQ
64oq7Oha180h/7cBUodIYiFnE23P+I5hYuBfi+eHq0pePdKRFjL8YfVhcu/s2d64
cZK1V0uh5EjmBPsVbXjEP0xjxF4nohjgpSrRXnZs/z9bxryY1hA1cCpr+YcwSUD3
wFjKzkAtkGtCDAvSF8NECHOz2CiclAvn2ocRjXKVhXldZCXCVWRB6TIX6l+c1jPw
up5wzpodxwEXZtt2mhD9ka1TUrOpzd8xHr3CdnD1DPzOSC+qaoCwEJMQvtFTTV80
uLKbLeP2kjsc1WwzpLaOUlCvMricuyFoocegnbmia17RZI8ua58KrvatZv+cgr6r
RBKSTbr+5Y6MQv9LDFtoCDbgb9Uwq8myJh3k939OdRAhFSd+sB0MSgZ7i8NI0mtW
dGrUITbA2MV1jF5Hj8PwemzlwX3IQ1h10Os2EZfSr4V0SVbkosd/jbPKWflEnJRY
+vPoeoW0jQuynvD6ZHXOdzQr2Z5YOkxdGbTnK4t7fEFupgknPZqv0K7FJ1nGyBY+
a3RvdugrdHuyaM6WiKvHxYHbRZ6gaXsZthrvBK2illlSCioja4LLPyRP36lGDHl1
Kamp6ZPr2tvAtZhvqFEKw+HKp5kI2WexN2kkJXYZTxXEvuVgmLMU6H7X2emlaHMJ
TToMWJeF0MYF0Flp4HHVftMv0iN7Zgx1uXvumIPWL2Pkw32Tn1R8YclEeQ/Nbtn1
4uHi7CDxlXBfgxzMD49Dyza8gyuAozs4Mr3AaMZ87RO7wjq5QoWrAve2F1gjcfUi
+GU4IKihHQMWq0tKsWVqECFM4YQrLy+6RTqFVmhzt5WctFFChYfv/yDdMvz2vepW
dxwxzGyJ/wcCHE3teKDf5pWzRi7gr3DFSPg5CpoiBETlmunNSSZxdreBb7yTAvYC
glUzuu+WAoWhSr2BSppmF4bUjalTeudU73X3PO3j9PDzhfqIX8LSt14JjyHNdm8t
bAmQPUox3figeqhvbfc5hb4AtU6aQvtLKRYgg1AZ3tSxNSDemH7sXxlvIU++GWkb
3f/4NFkLuf4rFxlGekZCcC4aC69dnmSTcdkvyrJ+cEQ0MPDf2SNHh2sgW34ufEdr
JO5duZt4u2yqRKNeInTsACSjd2zZlb55nPdhkjUFSyGgMVHvsgSJSMwkgG/QFGgM
e4XPS4kcq2l/fHtN9kB2H0aN8QaDrBgiuWWjzeIN37oco3SfCmOzUwvoKCyf3A8j
2F2YIWbBdppx5FBr72gM6Dkg7khBYELAa8kQo/de/9juoolYkdgnu+GRwmWVVfck
N33E+LJRYioy8/pDbGnuqn42ahxHNeeog/8hmzKOJZXah9AjpsUdiUA8AAvj+EdP
j8i0WGbZNHmCrBMnYmrvwDUqysX8BmRQwxXV1bqXdOTx3PA9LmBfsNUWCLENpU3L
dmrGzlB6lZ1mOyQIn0WFg0zapa/+W5ij97OIUIGHvtp0JlJjcwKPYjQvy3g5zKNH
7Ruz/CDrETSdX6fEgFD7eXJuj5w9FouCkyzIo1bXykkEYdl2LsxlOSdnTsyxLwZT
p0AbKNAqMMegv21Bf3eNUQbv8/BYji1yAfn62mwyx5KAofWO8Ou0Mdu8QYWW0u+a
ZdkA8wS0uDgVFgAKDE4prJDMyFSJTBFz1JbsOEWfQJC4oFw9vqxB8Wr7tugqfcR9
EMAXGH+gmdnsi9lZr/hyHy8BhUs2a4lOIqyjt0j2ebJFTrdXh6LEEEkB/D2oYNPG
fns0ad/VV378tZUzKzCJR0UJPpTq51RW02AMo6xmrAIbqPDOSCZb9KE8jlXv2GFY
yr2mK3M/rTLcsLqPh9S6zGUeO+VrapnZNTU5zb7u0imBoztihC18PyyT3bhtkSaO
Na1+ni/89o+TThzuuEpH8J3Eh48s5PAAiaq0M/UqP66qLhWUxha4Q1un6tfSgC6a
ZTJn3afW7SqWpasGTneziRKzUQXUjptpyje7SY19p5lU8FkeWAVhbZUZIPNfdklp
UuMtFsKChHpcpjNSlhxDYbJ2T52+5RJNofjxCjj4qchlYdYiuGW5N6sKl7e82gEF
8O88HUZmwnLkw3CNGVjDzgi0aU3bBSIcFW87SSSe32qWEpskTJCBFw+3L59dZ879
s6rA6+Lzxn2algR+53IjqFRm7y/7hlaqCrGfGLljEBiE5XnPM05bbpbK+Z7S4iAO
qRDK8s1WTeDAGkZRYiQSD4DbfUkqTRkVgTyVSc7sqCfAtW+wr6KNIXnydX6yQ021
C4XNKN37W85qF0VFiGUQ1weNtXTzxDcvaxUuTPR9uZuF6BsfPt4k3iabFsKC45/2
u1GwyT42WytWEZ86c7iwXeQ12hASHRZOJwt35PgA/xZX4Oh7lfbi64ezIOIW8IHV
c1TS9zqwc7XwI7FN0Lr9YrZNLchh+hrJyYMiD7d/Fv6jhb6D1BOE3VIZ8O9uFFtC
qtqIDs+yiPHQ/xXLuAnybfJGXzC7+J1s5CsgxY0OhPU6EQYNAZ2lo2foYe/n1Mzv
5tA7zkSK3oDzmWRJ7rRjsO5E5F0ufFiquXow1Sa/KcDRhCETlT3Tl6a01o1+/jzG
nxrFXDf/kVlPBM5u+pB+GdO/R65C4d8nZOjWaBA91jdtzJkMgTvLf0gWlXw991iQ
MkG5mdwLjuNCzQlPBEqJ1bEO71vhqPrftCztTQ57fzwLji5ygE5GyFNX25cmXY1E
0hIiXLFECwRM9Ts2/1+ElMEt4eybcj/dTe0FVH5Gl0YGZTK7r/HVRB8L4USHPJ5q
e++zrqwSdJYebzUXWLuvtVzWlWMsPffEVGV8dAFIE7xInJ4ajMP5U63dvLwtLKwn
3CdDTSWLK/uJHpjz4e9O52I5u6BfamXA9Q9J59vhnC39yda6TVa9h3i57VHSzG+J
394Nl6c+Phxkt15/k/1Pke8mJgUuu1QR91R1GIeiuxE1YTDMyzeBOUEH3mjRcVED
eYpuacGsgKRJcouy2LZjEdnOoMghs//j1+rvMg3fW940PLCTs9ESi8xMHYZiJdMh
k0pYngXCdITpuz3qSB7ps1Gb8i8d7P/XGZ80IVeHAbeieiFI034VKMjwtsQjem38
Fb3qKj5mx2hXsxDbvxXFN755DQEls/zvJOLXRv+IVTzSbCRDh89bF9JBjYa1XDAi
0WtsJyQmcmEMpbrv+qCQZYPwa+muNn8KDfOtppjwMF5NcIS0Us0egtgfNRs1mJO7
iSQ2ocAe3mk1FdGT5eLi0O0+SSGpio6v7FKdnuy6YGFzvFs+BTU8wpQzyN53m+bI
ST+bIuyPIG2goAO/Af9hiEv1issMuW0hiMnmxkTb0DRAD5PAYiJVMIyuR0ViC9C8
4ABtwkw9ek9pCu9HSaAqTzBqra1WRioGgDGMaYixuNLYv0oPTXTAM5TuS0uDy+VA
0oiWZy2z3sw868E8eBy6Bd+2bGCy4NofL2tQImPibuJS3ntcEinbJ1bG/lgf7PcJ
CwP5pAOcngnOWeYcObQAce9EgRtPKlOVXwlOXz99JMk5UcEaeu0bF1T6HASZo7QV
KMcwmxReqn+2Ap9OQSICtlslqL1+YPujup5eFTdsiPxu9dcJl2uDMZDwNoi5ed4a
bgwv+BLvu5dlSp/8UOWeJGnn/2Hvpn6A+G/khiDtHQ0MRVVQ7Uu0MfpLHaloubv4
p7EHSTh/VU7alpHF/7LqEbkmHOnjsPVJ6ZURiVbhMbrvw0XUsnAIxFF9fsIcjerW
/flAki4QrVN0YeIy4SZUUNW5fXHF9OppHH/QFhZXo3deOI18K0swmSS293igCLHV
IBYDowUc3QDxBXDZuLzZqMpzPCfyWpn0wzF9IIIwH8ke+PTjD3mMRfv7Zzu5dJNI
O95UYRNrbP4XoSIwovwjiknYkiK+oaVwee1OERPvFKeCaGwxVazh6QhjTMj7hRKt
UfTjuRqDqgD2ipOMHP697t4zI3eKUoyeYvoS+my2Bx58izmPLi7MjmxHJE2xx3Se
m+1BTZSljG8obHrVHwQXajFyQ+cbqMHgW9qzps2l3jGK3JdzM0LJPFinraTe7+62
vLBubohFmwwCYaSyJdoJwth6pMWDJ3tTuQ83s6cnGYIm1qYT60bbkOVh6ERhCX7g
k2AhIjEmDb/8qf6J7Pgvv4o3p2JgMZnHZ6livdC++iS6FGbM4uO8ZRvJEA3I4LdB
976zXiWXlBbbzsj1HQtyZswJCU6Fj54SofcijS1S1Gr/UCkh1HdRd9FRT8RTlJzW
l07vj+N+3riRk0kVqAO88FL+TahpVFXu/cjujmx1ggB0BVDgp3TMIIKxmGvc8hJA
q1iRrPNIVgDLITPKXWcM2ZvFiyZlOS86vbK0fT32Bh85QfrEvuknKfb4KyHL04in
q7xkKl1jaV6a/2fu7K3JRmFXycriub+MBNerN2vTplbVIUjM0QpGkOuDRsn/vJKm
2yj4ocHAdTg4MjZ0ICvGFTbzJLn47tvZY+lozI05ntiKUk7PqvC+Y1dCTHMCSejT
hrNvY6D5vZxwERy6f1Wzl0MdkSVh//dZ6OITAsZGJnfW7Nwhq49EZdHzaER39+q9
/YBL/mKZG9H3tVik+4pjH29EN/hrY6UDi1qh5nzOdqlYXm3HutP69JRdx7qNvAOC
Jw0ToAfICe6sscxkUukfP20/iCD6mLsXlBPCbrEPPf1IqgHc0aCol3tD+2JzgRqc
p8ZicoFks5f+mWqlYXGrmd2f9/V54wLVL/5YEa0uwVfaujfzWiSyKH76UWnIdb8g
lZbyhKLCqIbkWiePgBYr2kZ+YaCfNL6aH4PyRHAni5q0kZW4ns2OYilKOstBRDcf
r4qrAfJ6Pu5ZAGy+XUTG6IyT2Cw18gqqix78e12pbb2TS0mPm+1xG/IqcdZn1F3Z
HQCEGLoUYn160QA9TromkCGy6scPKj8UfXsCu5N6N+yHjbhau5Ya5vDt1e6fPpvr
3c6Cy1a9eon23RzDYsOue7pABghzS//fXOl83nC0L7WXnys8Vhp9bVzKLNSJejgg
wzXDXE6xgX+Q0EK2rcw+IHYlHCUQZDuInj5Ugsdzbttef7KVHnYTxuUokwvaNcjq
Pw6HpyNvsefsFiC8TMEwA+Tc44CbfL90fXSQ86jbkgc9/z+x1Bx6m9PDLxyqMQcz
8h34vfh+M0iCs15diAHxa5OwhCGMKBKGdW5WrYRa6GBx+jHuEyyxdkwOxtAiqsT4
GTFmKFjo3nK5hGsMDSq4EX7e3Vc9coT7xI5g5pHwr34VbO/N67n9ow2OhQi8CQQB
7z3sCjEbt3N4oPjtaYPWJGMxcpmjMSvsGcFwt4NTxJ8LhusRnnSNf9fCmWv7CdvF
rt6M6pdx6qoLRAksTGsbjYFdz3Kxq+lD1+qPVx+qdkG/nalOdWH/W8D3h2cPdOoV
pOtqUyTgWVOFja7SukSkX2ejNaQwFm1NvwQ+zTMT/Ymyt8cz3MGtrx2yZPevvfZH
d0Ktfv48w96S92zkpWgLXij1dpuW5096cU7/aT4HCA6Qt5+D1PKKTwBnCKrKQsba
7+bUr2W9sIWsF/t/bPsCQsCDJi7FG4U4Wd+TIxfgKxNTGvH08Y8CpcjSyTuN+/Pv
bL95ms7Tt+c7Wg36vMk3NuEklWe15Om6/RmK5cb3jMUHu2FpxjGOD9XER2Lt8QCZ
geNR+qRM1bmRuqGewqoFfrKUDWEKsvVV0AlqOq2fp2TtELb17SpNXYgwMftQFmxk
ujzv9XuOk7NKvBjIo6AVNNsE9ZoYQ06UWE6jvjCFC/y5aAj/8wf9es/njUnw4Ihp
8FGR/o/ArwaCTUlwTFnfoF7/xh/jju3XH5+UGlJ+JbCgSIRagadZsBiYySfz+gRB
BCl3oHHBWefa1K+lQOvUXjNsBqd6x9COOe76NlYeLwmbacOutBCAYEMSBbqucphI
/PVJE2owlLOqNUGe4TLy0xMqL3NPBL40QKxhhmndxDv72LhLXV3ftktP9Vd/bP43
RRd9dLk3G1ScWfbljobXVxL9l/q5Qu8Kpo3DhianSMcLdOw33hFLsHrC03dtUc9l
lxeyvX58JLi7LQaKRsoZvKIxOJzWUhum4mbcMTp9E9tG2SmdafKasaUJ4YFGZ0ja
fmrKIz7eNi4rErmNwYf6oRQLUkZkH1erfYT26/UY9JnuZ4R6UABzpiOZS7AiFdzk
V8RkO6QENXghW+sKSPxbOnjc+b3hwJBzmzEHbJnmwfF5QuDDbyay+nL2ShPOZESM
QP6XYtAsIMb/1XeqV+ik8CbKBVWqBnQ/nk7G8W9c1X2jQ3Mqi9yuOhy+wvucpU/q
569vRQo2t75dWdK7GsfFvDfYwTz9Ty7yVgfdagNihLw8Sqtmd/Flpu4i07+ZfwAq
+SxE00a2ZSBhceR4peJi+VYiooitE5HtsfU6Peme7iPwl5nnnX7VQeEC0K4rsdKz
BsraxC7B9RS9MTkz29xTn6wwozhmZfQkePdJxIrPPknWuYFVUF3zH0baMvmM13Qv
1Ruv0M8YKJE0qzKAM5rEwl5k4oOU1qh6FblqlSY3nhm9tln3XwKvUIv5sEA8Ysct
fY4SLnc0hxmSuqwUN7rijw2ehRSoWCHlLnGEJGKpuy+nbkXlf/IqdU2mZUa6Bi21
jj8RTOfPVPtxusZ60tYo/gQs6dv47NiXcq8W04Z6kPBIBjGz479PF57Kae9XWSyj
WgAJG2Chod27vSx4IVA+ROu6DySGOuEooCdE7QHbcSjDT3YgDWv42kdKIENkIhh4
HJ5tLhlUrz/Afz+vEwNhS84dIkO8MbcQt08XLcj92eTsGFj4m4l+JhLwYehyZQDM
doKMEpkRZJp5H4iYk7Ku1bjRkpbt92wGESzT7imSmos/rGM18nURQ6Y31CCI0F7j
LwXRIpbQLa20UMNw9E1molTwlzQvAL1GcXct3mljTp4NZ6GmTy1EUXfMOcHUnZAY
j24zt0DdxW74vdNkfHUQFnlTQMafO4IuL68J5q+6QbjziAEXxSisj0YoI3ZK2I8X
oys4cxw4hU/91deWdjioYWDFDcXPAhWAkUclwLbx0tZBsI8B0IccSSqeJDK8lSAw
8SHasI1EiWTvHEyKqkUhUdjVxoH6DpG3nV9PgPc2yplN1mH+uBEuRsgcLKaCrCfN
v1w5Zy03Xh0N3w+XUXp4nUAsgs6WtZuB8TaEGC2VXy1PVdZOW2soPcNoR/q0H/TD
WlFk4RF/0ItLdK1n+/mbZ8BhkKI0pIn5Jn08NqXHTl/01NCKEkiMLmJgvVtRz39o
RsDFdHX0/cx8onWzqeO9ZoB2LiI5UVc7qLF/SaSlgS7o/5gtFHtaY0aiCf+op44z
GxCHLm0V64o3drW5CYDK1KOHnD226QeEIxwTjLrO9UgOK6YlOyuL9Yed/C/DQWP+
zANN7T+yDLhHJlwwMilqOAUwGga4fcXpMEWy17DoSsPy4CzWvC6bBjfFYYUGwxu9
+WkYDMSQl9hYpxmqlSDxJyodfmj4gR9PALbQ9zi0g+cy2vNWgEdY+DYjZzZMjsKh
dv6DsUaCo2PpSfidcSrjII9Hk3djP07no7uCBLWPJbEzAwZqc+83t4d2Zwmej9ws
23/vp0ruBSq6bTebAY5yOF6i4ajjkqkgGWzv9KUVek1zV/aYeWz8FtSHxgZrmqm5
qFsGVCNdn3T5EKcfU0YMz3XD2zP9XedRrAcPn5u6gYJnY7iv2e9HBBgqqyvh/DXG
fDwmBjfJ3rbrtF8HS6X5zN3OZNY06oT+z4dW+YXGo66fDjpp/KwgwJyeRrAofrWF
iBLFHSQvQQJsXLdbshMO7VPcXbJKUwIH8kj95KxfZLxxWKr04tiEl96Uw4vF+UFY
wpQW7MplF+vhnYPskL96w3FPH0YKADQN7HT0QGhsS1Zrb2QKhekhv78HhjeJwsfl
huL/d3uLijva6Bsb9QlnN4me1PqfHaZYRLPVcn1/Qpr1dTWUP/2H+5qXXxlhOUpD
im4H6RDXI0IsnzyC3CeZeSDJW/w5UwJCs9joUO4TOsbmndrUso6eGhihjTxBUKJl
equLqltSuMgdybc+u9N73hfKj0KEarrCwe/iGUssXZSs+zT5in++bjh1tGFJm2kx
YwebLOqOFbB7Gap1muayl3p8Z0h3fhkaysyG7D3vqLhotha0lFKLAwzeALhnydSY
qPX8f/cXVJuKKfb6FEs9YM5N67HesRwaQi0deM8dsnMH/CibcexyMxlYdJckQuH0
/S1y9m4PGt7T9Nj3cIgRKRWqxnU8WbFeaZnyy8eeSv0/xWDCr0hUNbHZvp32i9zN
tnfeiRTVBurMfkS11uXIhEh0hgwyQVFO+f+aAEJztOjRour6ICdYX69aDdEGaMtO
iORAoKYGB8OkyPqTOQ4dElnk3VZEkFLRRdoain/XIhsKsNqC41y+JFYVAS4wlSRi
h3/OWWJ700EJj9smBTKL4V4bg5uzkHOixjoOo2bM7YCHT2rixZMYf85O/IdBn+Qa
VPBg4aeIXS319tPk5BmhKnqrBcZYLyv3qLPvKSRS/D7v1JIZ/IoN4K9niLLtURXh
6ab80g58lJa+jq2Mhz+7TNk6w+oM2I37YTpJ0BF0w+IdFminHakeinFLIKm7fFv2
LqBd12irqhmZjusqRXCO1CmQ0i0ea0EfMSKC3lWbuvQ4Rk2UaDOL46NhEMXzPCb+
rrDoz3PCEBAtF72KIysCk0DtdsZrdImPogOxqSHDHTTLrkH0IB27rCTL2vX3micF
INZGL7K8vw/W9jjJU5x6BA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAsZ1ijzmzVmeDQ1aP4I+37L9TCv2tWHx4kE9XL7X2VBQ5S3zf34zSQPBKQORW83
4ro/+m6aEPugfPUZRjR9sjSkXPW0xORbdixEx44Jz7tZp/4X4QUC1P+qCIyX+LbX
ui9ffmakfvTVU4JrAWOYff/ZZjmP07Da86VqkDEPlBGCL776JLza+RSjk+ferBCi
k1qaQrPGxcoxNG2oZYEncQgg4xKykZLTphC/s9/YZVzn1ua8PGoLqgagtni4BgiL
I+Ry+6uGLclKGt6wxtUHyUGKC2YjrJcirWcDiItb1ThGtCzN3DlTL/FdDSB9wjsD
pJI16aBdQa/FYxu0ImimS8UQ10eqfB861U8FgB4VxrqHCOubFRGTGBtbHFyV8eAk
Hu1l14KWTY2IbNuqvOvMj78wmCzT+tD/zkBxegl8dyjLGlEYQvcu994fp1Eox7sQ
50Fck1P1knGdD5cm+z4Iof1XJROHCWWiNCgNbGEqbVcxvW1ROyqaP5g1YHiWzspM
1NqAZeFGWfvYVJ3XBTEJsWrfxzCEwWqi9vKzORfPfc+hvbPP0veI1l041gVof8Rv
JWgzv4DyUnv32ryxy+ubABQxuNnNdzVKuqWSwr7AWqYfbXlw34FUEkJHIzNAgpki
CBy4DZEcV6f198FTPhSJlFA6lX+uGu9wuK+vkWizTHwcCq/BsTNrUBFa0LXcdEPw
7+wwOlzBH53/VQtJX04NoXc9a+UCqSXIQo1AlFSRr3ckvHoSs3D4UqgkNSQlk2f4
n9w2B5FztWW3Nr3lkI3VUZRfVu1TNyHGfAcmfBedr/bZcNOoKiRkwyjhbSLr5Xr6
hKybRLeL1v/shpXH64vHITNRGpNM7g2E/MIJOMkrweQfwKT+47JvWwd7t0Au6hUL
ZPUibQZo4XYbfF5HegSDiBnKg6HH860bUgJDm7NauQM3tvSMl0FGc4BjCXKGK/wD
5D79HJWW06n6fbS1dY8PT7yfdAK5pmGQmFJHRo3osl7RTA5DlDM4RF2BAK062puq
NGt/aed5Vha/FoR0n/6pK5EO/xKLTvOWVLh8/p7bVyM8Q/f7JAh8uqQzIZMSN+id
rLm6Y9NsX4Lj60tqGNno6TVF9TNUBj+EXiqgN8xzox1g/d7jmj+iFzt40jdlGOQV
ROiUUpVzlMajboDHOLS6R5XiVbm8J24T1ZnMDGmjpqKgPtQRODRpnesrc6znAnnm
+lbA/urAGRmkbspIfTBL5J2XaEoDBfdAFnkL9np2hehLLVBfNmCFDBGunA5XziSo
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGsj7s2fJDVOhtaNhc0Y5iMOIxaCYsdsC3/f8uUjzlhVw2nDS2XzLLpAtFWQiEdr
5JR9Wct4F9Ubrvs27XZaVQpZbPQZmZKTqCEA63DNFw3VCQxJIjxsUj6cfYWpjYaI
cMJJeGKO1rJn9pT+tCEr4CJlrrCgA9CMSdACVg3rz5EyOIihDDeM2AEtTqicxRFK
DBHz1nn5pOoj1gBywlRoCbJE06Mhb76qoI/YqbBBYRSPUexEALSk3WGnL0/+xcSR
pg8FWBCx9xM7hpoTKZ7rTSt+DattD5zq0EuGWT+L06IOTlvjEo5Y5nLCWOdMtSrb
W3mTEVbThxwaOZavzv02KPBP3Vfo/6rK23vL3ee6TLRhZJSD5QIe+UZagBu2XrwB
9uBGVWu+qoDcylErDAze3iN+wfup4WV6QPozqiZlnMUxN41wJC+m2ffOn/3F5sPn
9234lSqWQWJlHKcU08RPrKrirTSFfuS5ZTGgVgxM42jbIuBf8bax7Y+twzlHDkXV
ryfel6ncEmhg48pnoRA9EykHt2NUm049sGCCGQipCpulxdFPHlGQJ5fi50o/F2Z8
fyQVMsaGzUxuLgH28U0m20UwDccN/VKTqSQ7cQQTXMeNNISRJGVT/nW+h4LVWnjO
atBO/N4X3Q+JxJ3H6QB749pkym/5MO4MnCf7uH2kf2NS23e3NWaF3P0r+0aohqa+
GKoNgKATdp6UnVW1JpqDljiNQOmKZSu6Jj9dWs8ujYizKHqf2miuv6gsAvRryQga
Q84BfACrJh1ZCEJnoUyT+Y9h1H0iohPwESIQfqSeYtYO6krXiyR4fF8B3izu6T1K
xYgeNv7MSjbiyiOjJhOUJk4+pvC3jpEhET21PJBVWdw4p6K9r2yzqAJrRaOSCFuD
DXJ7es11qGMVMFEnZFxWe9dbruA6ZxJ2nEtT5AZTV8rL+REY87KuZZds1VDBDL/a
LoAKzEEWKdj1NRF6Ki5eGy3O2sofkTeLjSJ6oVLgBbAGOJKxTGtO48KShF/96346
/nCgBJDysl+vLX+Yz30RazFrFpqafcygLx6o2A0310pHSPCczxg+F1arWl77iTct
Ig24jplx9Al84ahYVRjuwTSyh6qbx23iuYtgWqIB60Hiu4wz6i+Tn30X5hj5Yw7a
2u7p5pHQjyqIbubYhrLaB63D11NJRF64ZHlDjbacT0+uMvYUncb2e9/T4N2tFIm7
Dwq+gGqkogDWA3ozlE9QurWbTYemwInLQjmAnRk1i1F7suWvRqlpAkLX81kyRVbe
Fqz0kkFkQjaR33vMsOT0woB4PiWaok+reks8VcIyf7s1T402fIp//wgigHQEhmD7
xeUQDpgt7tnkMR+Iy2JCUmJQTYfgTM4//l6cdBgF14j5s2woQcwMwIT9ncHT4AFg
6GjdbntLVsZ0FcFt9/eQLg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UqZE0i2NS6fG5vvXypDJIuVbe48GbJKgknX0A9k7VS7HnaWBkKbXmhDSLeH62+qu
h9wpsQXKbUqEMdq6+DqiVzDd5Bfdsk5sQm+ehtfPhfeTOiJS5GluaZa0imhX40Gm
7Rj1UqoY7XjpEeAoexa1zmVlhQxl0oDYf1EZLuWHP8jdnNU/AKub03c/nnLjTy2Z
1sbc0pP4HO/A4ufxASC7wJ/pJsxk3UVCB7LgU+zXHekJ6tgP3qlFU4U+wnF09tT7
gz8QfF4Ddy5oXVwEiJXi/SGx6kdf1IbmuekSWUQN1VPGRIPWRDtZYVDuxTfVYpoS
z4/YfkxZdbnuwRdFSPyK8YOFmyjTQRjcu8zFYMhwziOQ4FEYQdhEB20wENfuhOt0
sg+gD5V6p625svlRyEy3Rv0ZREUEXK+VvT3NvskIi5w+hEu3AzS0Kf8yCEtWMyme
Ig47sxWNBWdWiy3OtyjFRNcc1g3LumZXGiJntRK2kd12+S4wCtEZGnCrWm4RV27/
4dK+huQNl8DiDTFJr7N4E0VsBOqDCVuEAxpNAcJJLCt50PO2yLPP+nOdo61eUmAA
5B2AwfddxMlwR5qErth98KTbIY1CH+ov4NZfnIjNN25hfagUFsQtZTBLd1KrZoni
ZzQn/n1Ea1pn3b7RdsKO7rfpkLIn7ic9wu3RC7OtVbvhqhyP1+0huoNxNvSKnDmZ
5cM7AzKejrnkoIGshUiUSQDLHDLhfyE7dDnmSL/bowbZTtTzlgDVGrJ2VgtcdulR
580WQ6eESE3NKlJ6Hg5hUzHUPhkaNCczlIOCBjRXavVMFVoeTcz7VUpfrlRU859T
0UeN5OK9reD/hAHi1+IEUkQGXKGNGgIJFnwyRgR8plLTWgKZe65ANbZcyUzgV8tW
MX1PWij3u+tyMVOEep80RbsoGfrauwhqGAkI+0RLW+DvxmK+yxlVuG0Lb/PX9S6t
foUCoRHZlYKkmaeoMMHJ9rLGLOo3UriJFkmHfs0gZyYr6BDC2CeiygIibDXVl71O
UMxDOVlJHi0h5lRSAgbc33CgXsDCH0p6HFF3p+vD3HJvcEGW/qaw/r1+ATzQPTqt
dBw8hmI5BPlvAtf/S00Rkko0AKD1QYe3UhbCmzuPgOfeWIcK4/Xy7mAdvLKv4dGW
XuyPQHKSpft8W74fucXl/gPLixFa4+qZelFiytvO18R4WfBF89r81WSruAjrjdpW
PelVn0UFm/1xk/GfwC7tRHbWYehLn9n8IL0z780t/wn38V+uAuOCTLxs9EGRTJ3O
dXzuAUySLyLlfvjAB1MUZcmjShXkIU1+prjdN/d07CpTnT/UmqeuOK1hAF2fGCbu
xvP6w7WGbz6rwYZr5C3DcFG5n/PNKGMnXq7w2jnaDB3c5vCpJi7RCdgSmRCnFAKo
RY1//A43tQskUUO6vjxyXQ0K6zYeyQuAcNK0oaTEa7OshuEzEfQUFQBW4WeeHW1Y
MBKfqGfYJjGVbg1dJRxSK65qEZliKZgXfQ0K5gJBJ3Q1P/jKcm1T3CvJr9uCP7i2
fr9hhbL40l2DqzsVvKH9WdAmxRr5e3hwuAbUPH1Oa0jbFN/pQhbTbihfmLKxIBsI
8yt8syKfUROE/oOtmuo6DWk/3IEfLaqtZYjBoCx5L8ovy2ZbNg++KrJQlmY6LTI4
W0TdTcGFobznnsN+xqj8DemR2qm4V1lNBK2sN6wCslMnTVKSHljBrbraoxnc5gfH
9cU1kjJAUJ981LBtFBgy5GIFty7nBaCHObQT9DRo83cqyIpL0R11B06je1l0WY3L
OM4AS8cPwMz2GTk2G+QC98uF5i4YrETd9ILzmJcvSS9Rc/bLYDjcoB3PMvckt09C
uTZiI/9fYnZQymwkCMBKbAApBONgKVbDW3r1764mNkOcb97HQ4ZSdAwoFs16ie2G
uz4P9EqFj2mw6bAOf831JMHqiLHdK7G3BPTjRLw9vG62rAk44hA5n+7b89U5Hzhj
znG8nDDT+5us85qaI1G/2UqzaHeU5KqCf/ng7o8q8xkrlulPOHyEuwuPEZDDyGat
k05VdS3eDJv1xGO23ykW71Q7Ehm9Ho7jZd4XGp0yolYDCaC1jMkZ400mRQpyM0q3
IMeBBFA1PKfTuclCTUv7o+AxQhIyobeoh/So8FSwCusc89sJD6V09UYY9qVsIBWK
6sKzumXKSP/eUcLZ/o6/yn9vqpws4CmisoV4nfAPX9QF1mvp1XE0kr2VApL9kVK3
tmn84J99u3sVSjszAjFDv/H7l5rHO82LG/Vjir+vc0Nus57lMoJDR9ZfNodwofZh
us57X+nzJ/BhLujUx5gbenWeW1W1eFoX6IZ0UqAyS4r3V83SqN3yOAnKQzrHAxEt
eYZtbp1vTfycAS1ZmXzRfCMyY+SK6P7DqeB45ibFsQCaa40Yr96s/J4okAoQp2Wh
HDPasK2/0gL3RLHcJkp8dGnQRKJISC1DlFDJmYVHcbUcvS9ZDmy/XuNdwMCOkWtI
e6LxSUnZLrolS8gZPeRa1o88gy0L7P9T8WDLdi9bi1m75r5KTCxGbaVkhJNz5hj6
+tpKd8QTT+/3GIBzDqmCADZP6fPwwJXQpqducqMGmzDS5omptHiuVp1n3dQzgCfM
kU1fhpAN3JRKV0uRFPVp1HMlVK3XzvrwL0xPcdNTnGGMHyIjPTNgp4PDOJqkrdxw
uurx2vB6Pj9qVKIQunFvTTA4tcKe4Oufejg4vpr7sRueJTP3XThohqWzpvLE0EhH
x1S/tIR+IacNpQsY3XwsY7vbwvrJHk+X1NhJF5RmldRyxvdKHLM4MmKdWkqOlLaM
FBXRMBJCq++28QmCus7SYSjpRBWBxfOv1RGrnWqytt9mF396y9RL8VR+SykMrjTg
3bBGY9VnfkRoTKffNsLqgnmikBedwEg/UBOTVqM0436M5mGkC9eILdB4nth+6vEh
GEqjvaWC8mtTV5p38TeJFsulbqODvQzU/lErAZclpDuRIS9jaarZJTgebaE+3upJ
8mE6ttm0pccCmBp9asTPEmn4PIaY2H6w/EUAkXAja9AERt1h20/vOnV9TmLe9FEX
sltERtNfw5mGKJSo9AHB/vTmDc+ZYVBVoPdlwOD5GP8Zxdaw0TP6Izu3IVBBlQTZ
Zt3OJlsIqX39DxCi2/2ImCG3RCXYHhQOGzNQzwCbtmMO8MsM1ODEievViRGNJz1H
VjNl7tMY3fXNBDv6oGgOqrm4lNtpfau2iwBLoZGt5VGCpNeYDu5WoFHFe4N9Slx4
6RztvtGqKqyJFUeVgJiUhp4ec+cxhCMTZdRycKVoNYqbQbMZKZ4EH/j07TW19k7E
nMwhslTTO6BiDFpGmuCI1HNQDoFrL/PyTDiI1oN4O8BHOsOxSqWnXIAR7R76ylpy
ToE7/2hExw66rD9b9ZlM4IzvM0sXjCEzvzvEqEH4PC0W0zIb1GOsRmW2tzciO3wx
uyCDf6SNbL+7uNT2PjNCpNOFIQy/f9snk3/oithODXVAR+b68Qe6cIlUV+GfLtb9
MLzH0I5Sb/2ojdfTbMKNackemQRpIdYWSyx1NRZVOAY14eYSJWQkZTtgPGqOvjmg
CCPdqXrYyZfAxD886zFFx5ZYcxAN8OOA8B42zTTXJuhJujfT4mGBRWzddnIxm8Ku
ZskolBRVCj0UZ3Lxk+XQX3PZyInUHE5dRDAhyuBIbC81TwHTMvjqoleRzmyKCmla
DjoJuAsYUBF0ctjOaKmpmdTOYN46T7dhPWJb5dHrt0bKt7wVk8zo3vAlYBIO5Ypi
zXxVj4LSr+YgN2kn49Y03R+WUV0xj38b+3DYgzrfxRke5WI2GVB/C7IE5F5RG6rH
ZKY4ayOPelzsXpplkM7aSttiWAk7eHtx16Z5EuDHuZVs4pw4OwY3973amJY15koq
NNay/6Rbmflbcz22+GbinmiYERwGqZLDx8bsrO9nTEkdL2WxB6SwflOz90rJ77TH
wpybw2L3r9kKQS2qdTc7NVWiPsEEXcRhFHsnFKOdvqj4BnCBUJL62kGApOZ5Qd0G
0o19KlPBrhXBEpx8WdfehVlY5jxC3csVh4vgdcFOKB1+yRt5bfYQ2fFRfsM5FY8+
yPbF96xs6+MpvoOmkXU//PFV33kE7GCWOfHfo7cgzP9eIPxI2CSx+qJ39VxLpjxs
7BF6HuaTIYwya0lG+AhCgACTVTTWw17w5jntEbR3zGvWOo4eVBk6sOXqwSbibnoh
dwx/fh+07cW0TgmJ2TNN+pYnW0MnCdjmEw5mxJJ6cDfxx4Od44Q8L0fMnOn3k4mI
ShhRBQQLJ07GxwgS8Eu4FB/7gez1u7cWZSEOWhzy65Y2vLHoL9iqBeXZKzzpc/e/
RQsgdgi3O1X+JYRTSYm8O3B2ahk0u6hKk3u4M3uP0QB6r0pXK2oCoTBeeIOZZ6IH
C8S/mVIEiKhr4Dsy7pG3r51x1mYVJtHsJAnRd+1oi6i1vQXxS/7o4KkGO4CTr/zB
2ohxqdfyqn4mPM6C8K8ex7bvbLpMjzp89ZQAu057X9JdpmhEEwlgT8dzY4JqGRDY
qZUjS685y5hOQ6lwqr43LQsbw9BydAM/dHrS6zJQBK1r3Ex/tOXlFgeIiBQcHDb/
Hsye8Bn+LgcL4G10nFLH8hVSZRlsajtSoDA4nApgQRkBl2vkAzGyoqnI7o/VL7S5
nsbd7IxlVoLatGl62iGuKSKMIEp3hfY7Xk5EBCSftp4srIQrbt2tALKCW7tYqJ+a
W8bs+YhLmPj0L+PNY4T/KPiwd6ZZ9+0ApRKGQO8/6aBUjmuyqYlUj6WJbbHrdmCX
On0BdELxUtZlyTUoMYBZiVHfs+lqX3HwM0i9qIb111v8HG12P5wxsa3MUrqK5nCI
7ewZ384XSFefeY9HLeVEEupWMsBdElh89nZotaXZzJI2CdUoZ/Erk13woK7bCUo1
BfMlzau0h22uTqW8ShQUuijJxq0wM5hNMgbsYecLMlMKsGKs4IN47QqZ2N9l+qqe
u8zalyT/18tidfpOtsIIr5+4/rT3IB2e8e3n6do9I63lkIePRcdy1HEfrMJxDBXq
VvLIgam0rvlZDj9y4ThpwAgvoREX6ZbezIDWdYvfxEu3jYZLy/rixBD6HV9dwBBp
FBTYJI7pr5xSw22bqZUCS38BhqbrNQdOL4BIn2QI3JOuCgHW8TZMjLladYDzSDKc
8f17ot68CYnJzxy6C1+z+d26PjhbcpH0B+E3CKifXlopuD1bdLDozBiWF3aHFSKP
rHl0VzhHp5mx0wisl0lvuoChTc290ygL/wYElasqDwCSCOFVaAm3DCckjTdwevPQ
f8IW8EhRTVmTPBuzPXvccyKwhtBp33uJ5xVmKY5f3sHOKMSI08mWyikyfUb9PtE8
mUyFg6z55Q5H4DxMgssOFejBu875yqCLOEhyqaDlZKv3JBOJuvDbp3T10W7xSKLG
bDfPxlBL1D/1pgEbSVMGJ2bd6/Ll89wSRcVBU4wa68iJ6HzK/+3i9n9Erjj3kGOv
FI8gq8UJ9PU0ui9bnnZ7hAuw/iT4sWkOjbWwmKJ0u+EX404MsK0Im/t6jimQnsOP
TnXLFAHKSr+GaJJW8Ohc4RpDHmNI63Xlkj+28zz83/FJHmgyoPdQnrqtdyHY02tw
tZ0WipAl7jbmeL0cfG9g6HeiSoC29F/UQjwVOUieIUTKyKVxOwP7EExkrvm4a9my
CgT303ZrRBKX+8K2E7U1jSq+dzlVeevv6J3fGSY6NBKQhK2kfdwaTpA96P2yb6Os
GlPs+zKQprI1ykmFSuwmdFFqBUAolzMIz6e6uXAaBDkyM2T70zWWsVksDjQkxPo5
5IB3s7gCKQRU52EUTtmtvlQrp3tR+wsKuZail8yt4KusNlJCzWp84zfnuGFcHRFi
2ckA5L7iUobHiGBjftc3M5m0sPDqMDU8EwXDuZ+fQ/UrQLvTpY4gQnh5qpft2DIL
HS1JCA+TpCqZk4xfqbMZj/MjM9//8M774OIDRUXG23/zhnITCfE3+xha7xfPqdRg
id+/GncO/Nbj541iNjY/rVg5J7gimHc9mE4bR3rGo9s=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/QQ7cihkR5IsCMwAjlj6WdSuf/dZ9Dc9ty4HfpenFFEyK0rwTVN0A3F1+HyvYMV
F9AF5JCVJqFKbQEodqPYihZvyAWieUXXvP9ruHkTKunQTHTv+5BeOD4qiACgQvWR
2XG2yT9u7dSqXXGRWGJeaNoOYo9QsLAN386iei9+mqjUq+7cZAs1c1jXNgCAFCoi
AzJLznSxk93us2CPIowJLWIv6MecLmOvvPalT/OKUPM3RdXYAUHO6OTOcTIVqZrt
T+1FE7PIWaTwCyryuijRjd8F22oio98oTqjEvOe8HDajJqtp0FhWNKq/Fy8LDAoN
2bP5Gwyxj5JScKcK2zKmzOV+C+oA2z8WBCm1Bca7GyniwpR8unpJzMRzNgYL11r9
DzU6OegLs2NdFmQ6WIHZMUmAnxoo3CnReNJmpVkpPAgdJq4g5dU7SdICUOMi3OxQ
9aVZaLZEXGRbjic4Oc3BUAuC62G1b4FSA7zFs34v4K+KDBobDG3HLuqIZR7+d0P2
rpc5jSRESky2yxhuCoUBbQ9M5XzIT43aTi5AlXX/I+KwohnHKJkeM1DUR0dAAoQk
p0jPPllkErTnzTou7/3KG32PYk1yBHX+iNwpCVkss2eJiIbycvjqeV9OoB8YXSQE
HwnAIaT/lXu8JkI/q3ShMPPv0nsqpzYMVxrR/tCjdFSY36LptmVZ5A+LoRAYiFu8
MeIrWvQfB70KdKTIukrg/pA19I0ViqDflue4HTSXb1Kj4N9+WcdU7Do9VAM1vf3t
Jtx/r1aEVeolcpEe+VLUcVtbFpx6Uj+ktdc7D2IX2r8pJXDOEJ81PKDHhSuDIOB2
EouE7RJ2nbYVTSjhAjvnXPrDzI6mLhZQ7wRRPi/bhVJEs7OcAQCugFOU5a85fDAJ
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aof8PmEjmaPLwO1ezSrsaGmDyZtJTHkLPCrQOVNS97pHQJbnikD9ie4tw++e1Tao
JGkZ58CwGt05CnIeni/+sx1/GtccEzcoobRyNyRFQWZCMVN3e/6dMXIJkA2+O9Bl
lM3BnJYrs0Sm2TGR3dyMLOBcZu+waLmI5xMXSaUlOzvbG5lX/kX9celRnXff6WpV
otDmgze6v8QOC+MTqy04GV3KbPLbCnwIAI11sYyNPi9s/DRH5SI6E77gIUk6et2R
0yo5l2OY9IIR/M+fzV7FcH5qN/9h+YzwgbCrniN5MEnNWoRMwvQvJ7KmmE1ih6G+
AlcAQlBQrTqhIy4q84RlOpWVY7kFz7Wk/PMfKMK/PpCiMfhJ2T5Tf6btEOTe0N41
0fZhJopDrkWpp3OGWq54V8hKS6hVffnnQZAlzAijsz5cs6+ilTTBsSGGPeP4dBP/
z0nTSSEgGi43/GUmimSpg9TBVJAiiPV6PcA6687vQ8/PXMrg7UUOkOL81emQkMw3
01rnrnIlxYm7mzOkLD9Nbk5Rw4cgbsUM9OB2JxEtqeyIg4RUDy3eq4fadWZ7+Zu+
YHqz86c8Tpp3D1oRPTcjDnj7UP/4E2S74hkco+DWT+R+UAsado6TEqHvxDWrwf4G
yDtLp3HBAPFuS/sMnxqX1+JEFXQVXsbiBFdcs9iYe8hamaPuyuVQEBcQDcC4EZ0w
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+k1vCuCa/THyv83tjcc63GBHg0AqsAt77gSEPcUJwMbN8nYBAOCzfXYeNr/y75B
B6qc0RwwL4hOhk8SKSYwefs6ZmuLEiT12hYCv2Y/9PVhnUClNcP8ApNtzaxg4+Ro
QfOoJgvoSXnMZAMfKK76vzApS2IsINnFtp70M61sM11+e2bpXYOm0ZQW7BfWgOf7
UE+BoQOGjWhV/hnzBj2BrEvOBEIAjF6Mszpgn9wvp0ptxqKTeU8p60BXhZc64/aU
AXuMxEH/ZjQc5CUokhWuJKmUzHGHylBBBydOiq2Q9Am6s7kpOnil2kAempApHw1f
qNg3zHembpgyV6m3KKy8l4eK0ETRIaVEWE0X+pdqILthHi3xzqu4g3G2jpgQwPlV
YlHyl2fZYUBLy7TRGbBsfkTmmD0vIg8Dydrm6lREMhcCHfzBHuDVMgkgb99omRBR
7Y5/ZWkajQ3nLuc2GCxOjnb/VKK2uGmQCSEM4w+uK81u4HnKXKFS8rkzmY1htTY1
zCRgLAIMRttdJ4Hgk0aG49wzVh2AAhGC+2gYJ+f8UQiA/rE5s414YqtClYjEKbra
HX6VEY1fmQN58ym1n8yHpo9qPwKPHnJakLgj+oNGuzZ0K45/qi/Mf+QBAbaiOHMI
nF1haRUE125WZ2YxRsW5f/LkHd/xQyS5cvpCYGNOlzxcfdYECsYDXftOjzq4p3WD
RQZGaAN/9Y/TVDMRqtXq6PJRjTjT/UGx0z3Ps6VcP1+6aVVWFMQsOKd734egKUZC
PIRI/ZVnuuoNcx/k6I/c9k27WMTPwVLCsBxT6tYfB+KP+Dje82WO+MVGgOarxlBh
ug7YXiA7B2syb4m5TArtcv7BgXCumAyk47GLyaepu3W++y1MiT3su1Sy2bavq6yR
YnDQODIhRGkWvlESm4Wedz3MjmP+qE80/b9AM7/p840aS/HjXMuKEZ2b/aF2Tps1
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A1IY5Djax2xBkjsEduSbj4gDtX2U1WXAe2H3/THLekZ2CFvBZwQyqyz8P4fDTSIX
hmWUYRgtKNwiYzJ1maDVXgZitbxfqtI4q3GoSV0Csn9fIyo4q40TB6DUhzkrRL/c
fF9lDg+Xao1BrB0SJ/+21530+BHfO/mnX9GokTiOIJdgmX7AFhaMWhATL5GRkyIt
0W92B1k8DBZy8gPOxft6ekbLP0bc42fQK8lrjRhUhRVqPEZ38r/Ox5aGkcW12FHs
DZuAqfX4+SSqxaTySYOuvhEzmDvrJ6jlsWaBCqQYQTlBDR5W9SxpaaN+sir48zrx
jECVcTn66xG2ESF2mNgsTT7Wht95+sezMpRL9k6U8fW09MANcoBPkBvY5uMTT4qU
p7qAbhecBzB6o80u+i0IZcyvCGwP8o3PKWo+Z/ISovOloTtIptMRNmzRtcgS4vma
t6dUSWboqSPxotnd/QQKVM+9QypQhvz1Sbu7tsnM+Zobztn9Cu+4xDqm9xveTOh6
3BQiREdNKHw+3kxrJNXpOByEonNrnBZu1eCDXVplmIdZ2qDxtUE7rPSAT94llkSs
wZ7G6sEm3H37zlMdbxp83goLITljxpqjCuOaUbsy5HfJH58E2s6ADhj9EiTmubaq
HPF2YGdnTclokY3qRUv/JY0svQyv40rTngTY4nmtG23MbOAzbMuweANAGUhO3vYq
dTK7wJSLOiEkD+n4zwuNCoJsU31lUpYKY5eVW0IpVAdI8wXmMTcwFeMamKI2UeUa
c1yAKGw7U43w9wiEKFcCcB97xUXo6JU6kCgRa03SBhk5ueK/bepHSWhYm/4sJYA5
CRwqeJWy53qZklMHwdpFRtIIo58oHYIrjaumqbVkB/oCQZwBYcBiexj92r2iWZm5
hFmTY/tDire7BlVaK9m2cctmKFqehq5JvXkVw24QWKdI7MUO7kVfAt9/YOblr7Pi
CwFLLXnM+57JgRgs84DUxGLNmu5mMPAg4AjLAfAPsz6RwuZ7l/FEYUDPHsNHI6Cl
390is+sUSNdD2OYB4G/PvoPLUnHJf623H0bjVvLLBqwtpc4b329hEmPfXFVVzqeM
f5yFEkV0U0jBx030/7JsjeFQJFmmWg5foaPxjSzH+dcclxG7vORrKuAJwT93ZJnB
MF03+sQAIasxWPtqkcQKLDSOAhinKgzmNgTFhB2NuZAmIi9HHipc2Mc2Jnsw+25h
MHYwWIAhZjxC8njp65AONF025SKJ9nYvQ/aHQHGbSXwiWMkHIq0mtEyAULCe3EqC
kSj0DS11jpvVaQpjqiJ6I7I49fMS+feL1zaN8VfRKz0rR0O/eHz9p7AAoBUhrCfw
UMu90EA9w8emOMjXQBGMkdXjewiOYGpC6kZsZcixa/ZbTb2LUBbhEGx29OzknrtL
ffT05frzxeX8TInbvT9dxhSWGgoGoWi7S+LvL0ORA0A9r2rzPwHZXBRFmwq8DN8w
LX5CqOZ6perMsRSBQp6kpbRO/oYDH8EPHHFwRbyi7Z2qK1tIUhyY4O8el2ktbLhY
Gvh/AXNY1IY2wNJ27xoR8Xeikc1twHwcu3kWZoeqFgLVv/JI+qhlxBu4kEr3/SYU
nPVkOVZ7uct/fhKJInDyz0SwJ7w5+Xb/obkZDU8cGiQLX7foQnBTF17/9S6fJTod
zLuD82uA2Fg7KFLz365qR72YaS9jfOReuIwm2iNXWt912aLRaWQSBX4VE5W5g2f5
1lDggTuE7sI5kxmpS6HtybZCj+qaUau+8Z9D9H+6ndwaTUSGt7oOQz1cCo2C03z6
+qiRDJZoLRfAglN+KWD8Qrsr9xyn9xbdFgW/Hm/FF+7JMfFNdoNIAl5S2tPRbAAS
y5cV4TAhst6kfepbUOWg+g==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0JuXj3V04U8GIhfdgK/ilvTOcGWyicgLg1kMVhtHRNj/QK/E3WunLRCoQ6zT/oN
Qiga/prBcemLig8bMQtA6JylpqTdNyNNHYM1ldib0WAtKmoln5RwFXv5DU77bqoF
wxpaPE/tN1dO+apNfJDm+LtsdUVgDL52RchK/sYFyacUHxFVovYtNaz33JKzptWF
/z2RTL5T3LZHZS8ZCDQ10Ikaw56MKII3g9INOpEHAKuyOR7iBUnyvhW5qkdtMcBW
ktbj416HcKV8ogOyYEROR23HGMwhNq9jWzswk/XxALJHOXASJ/bCZsKEmSn9eVIJ
6nkJqcfTD5tVgILkF49EbetAOPc9qayrNhexH6cULqEaIBM8ty7gWxyOBskYWC8+
tooeYH2ymE/FDVCZ3Ipt2lgUlt5b4vuRLuua25KGBbCEpdnf1oiMr7+63hSSiHlt
+7uDW3bxsKmDLdXTvs4MexcAk/WQyGbM4wZPci2K+d4M6do0sTGxz+6/b1UUkxQL
4wUVRzkemUS582ns2k1VI5u3GLC3kKn3KtGtA+iBmvgLFUmZf9XntIfyDxkJQNAQ
IGs39MGgKf4r7vvh75018xP5cCQz3rW7wzRkeAjAnLBUBMf1ul19e+WXQ52JGq9K
Q8FMx7vALgAnEK5+yjL+BST2TxfBRYx8bqRLr/mHEaREAki1cY5NCW1UoE1jJStc
FlyIo3SgZsM8pzunamRKk8uBAJSqcFvfPDC2tkOUMGubDIvlfa1unombXP/gbfLr
uHTXCyCS+aUqFPwx3FZ27Q==
`protect END_PROTECTED

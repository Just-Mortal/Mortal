`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZvRBVek0Sq7InLwuEwQLmVnej+jWHPsL7Mc1rw3Y7vKEogc1hcVWIBAQAHe1MtSs
gTN+FsnwTz/s3DvAvT6Lx2hVcY235Fc8dT7RIx/WYqaNwvhZ/yOd2fz4s/84Hwis
S72CAHf2oFD/EHltEYuyIgzEmzLSyLOMo2O94s5meTkishZvljLaO+Iu55QvoUwq
yMfNPntU9ThnLB/nz7Lj5mr6xTHCVtkz9g20VIftDtM2kHEJg1BG/1BrD42g4S8W
NKfqjKiQ3GZer/cjxG2Mdrmxv3P86NB2WMz4rE3LGL1NyQmmA7Me2lzesOvd3Otr
BaFBzq/wIXa7Y06VZX5cVmxxE342FG1ZcuN3GtfvxOsqIvmKUCB8p6TzWG9aL837
M0rs+mXRDvfILTNZt0C5alLT/sD9361ocjbR+F8105ENWgP23rQBsCdKe9FtuftR
Nb+gLUPg0xYBaiaeUbTdPWnWI+iVCtB+gpi1gM9TpAFjqmsdV5brcUOPI2/6/1pE
tLsrSYidzFHAKiV0cgOeLU+R/aFC68qVmf7UFYqQBmz4PXPbMjN9V3J+F3L73PW6
GCikwpwqC/hDCinYeSr+XwhKLttO6JXPSuKKPmAh0Nwhw9cMDA9r6o5eMP8Phuxd
36V8QxVpGP3jJhcuP0jV5o/WPWtRzBtbVFApwwg3lCSKyCoOZRPYNYI0eY4dHW5e
nr72dy8lEOS/W8bocfnIOr8TaH3hgrCBzGm5quaLYWvk1DYZXvaUHLmXtn20NK/P
hbVvCp+uJDB8EiB28T/SchpCcCKzuRWQqJgHG4BAz4wvtDqdyLa1gWjT4EPqW8Fe
80os+JRjGyWlJzYkN16DMwbiEJ5q8lUWdbONH54vvJv4W7WALWLggtawBzzOah1W
W7oUmblrEoomIw9gWE4nXtvj77bQSCOlSgUdr8KJf+hWR6xrD2EXbcnLu4SANt+n
VKo+fxmMtq+T4YWKRWeFDkREnZoXPtuquXC/QCMvkrPJjSqIwEQlcx8weNIKIdQ5
CA+XdYarD5O1LyADnKx/s1M4AhtP+UnJ1GOnlG0xde/mQGs4lkNT0Yk6MWAi9G5H
Z1KVy7morvTwUGprcOaZe+r1+XqW0gwyvwYw3LDnsKeAA928giYMyjMqFeeTfHXg
q2jASXkeUD1tWpseEobCVZBsiwgBRUXgWMilo8+9oZCmAJwOkvzP7VIX863tMc/Z
4sFVagEKmBKVPx1IuDK0Her8gkvMPPNvW+NA8VNOJ24vvDrf7H0/kcM30VL0e3qh
5pAckPTdcCU5LFmu7g7B91pU87Z5jxFebYUNoIxeXhgXa00laOCsFPWSInj7JOC1
Mv0lQHkacmus9vEh9TBRml9SHKNQ56vaXa+igK3MnMMWEWjYR1pTsseZuj838dd9
yhvMH9VykInAaM32c/RR07/JqCIgRl/q4cX67esMPjgP6HWGoruXbwSLgGTitziX
nUntlVHq+hEDCDhMmNoX3bZRhqVKOzB1TOrG6yv+7w1GpIcYwsZB6aXv89a+D5ls
KYpB3/hYl4SPUSzwTjTSCKj3HBisUglqzALY4RfTCw5sKSSLCw0tVMXSub9r7DUN
JaWLeueKx/Vz53ympF0e5i0EB5AsPUIiQykab3LTH6vp4a5RSzIMuNxu70dobhlM
cZsahkfq85R9a4no+pker01Tcd/UmJLv+nwLrTilDoGXN91oqjAFYOQC0baU2e3b
Ore19UIKb/D+uWbsdKcKNDonqERGDD/19+IQR6asPq24sXHV1QBSnsK3+JNRlKHr
RV+W1oQufiRxcDJEdlyVqDm4X48gi1Oo4aJAWs2b0ffLqJHC/40aa/ZMQClzCJBK
PJAohcu0T9h6/dWtV5jwhMndiY0oqrBivINGvFaV42WVlx4fO2Sbobl0I6m3YM3v
04GdsAKNnZMpOrRR/MxEt0N69xF2R6rH+IToTcMj++uY9ndM1R+Yd5Ld/+ujwiSh
FqsBudkSeFbX9guhAH85T1njLjX9HRGjqBdPM5sgdx38M752i1Vh+QgigloQ2/I3
vRO3gNZ8dwu1Nz0o/i8Fq5pupTEYWK1Lz9H5j9E46DkDGyqvhAdulQ2tnVYnz5jj
FGWk4i9aGcOcIknDmSImzvB+gv0OFXDQYpIdrinT8lcREhKynUHlyC7NtjzJRN8I
ol7AFR5yXIOBaAqvanKEaJjWCxQCJvObJN9zryJH6CqpY/resOApiPe5vZKy8TJY
E0UpUwaxjPvCUPI+sk/iYvKErT0inVm96wDty5bosL+139dz6sTu3/UckYh1FsGu
JDfSc0B/9qZw+n5ct+LTDGWQVrXwVCijjnSxWm6m8cWOzEAmfnG6cMTrdMSZEgFR
QaU6jl6thJzqlwOhmEc+ne2SzX+ObILzsZkOMKl7zo60TM14r74gPBOZYNwz0y+v
NRvX3q0xQegv/87e+t/c8vobFvzAM/TIDaEGaOZn8gbSb8fdVC1vHREG9PBdap+P
nmq4pVvIP1LHubgzf2CRQwR/tGhQtpYIm1Inab+aaZuRElQ2fRUL2eUvqAESFWxx
kw/R/4Ejgqd7RscfODJwaet56jada+qw57c7TorXApPq+uCSD4Ul0bUG9upVuaPj
blsAP/tVuyAE9GD9tRdlBse8k1AL5gDiOvrsPjaICmKcEqepi6No5rhTe91IwCg6
m7afNinO4C9MHQDt4azE9b/chltMSlHmX1x6Atpzv+RruTT/CZ4vFYjTpVKl2Uz3
vQPHgAsRRAVcV2bqKhLuThpvu5qb+aWWv8pbRUeGOGz7LlyD3snPhBb2CIAEVUDS
Hib37GVCJ8zl8Bw+K/jOEHK2eR8K3Hfr70Lh2g1w1NBUpsTDV22HHpRhJkvH/bNd
uKR7Zoe+FU+/M8tVKQHY+8H6xfViNXbPohHjxsAqnP9zPAGNw/HXrRzefwojB4aA
QxDT27T565XbJ7xNFLCL4Ji0wobhPLq8SX6qjvRxihqYLsPZMs1b6d0ZeaLJ2HPO
nKaiYxqN/G7g0zrs821dtUqXZ5qpa3IAormjbKwVh2e6ycJAl+/2fg72Zd3iRzjr
IZz6jEifOaX9G74fyego5DRS12/6sq+tCps1/ulG6BhmBASQhNJUIkTWEYRbTUki
r8BWD7HXp4mS3nKEbG9deJxYp1PSP/133wM3RG9Io7A7R+Kj2kaTEQybGwJtdHu5
uO06S7WMZ0lEnbOW7XIwIuxSvoDsaWzMoVZPBnatMwHaFu4blYCi+94rulw/7SxP
C+iE7+XXGx0chsWFe5V2BdHTcEidaIL6/cIpr6uRyhlIz9LrIe9PMXrunhT50hV/
iAWnKJa2FfLB5XAbANFZqjqO6l/zPIHhSQZEjcxD2vt6xKrP/CwRACFvGVWer9NS
IMRdWRKJrJdhz7GO68lnx79F7P089r8TMPktnSj8fnqgu93aV+R2NjhQpY6m/XcM
9HOlrNHk4Wk+atBgPJgMijYlxmHfPjTQ9fV7r54373DinWHiGlt69ErjNIOUzxuD
AASPIokkBbRX4/3ZUbNa5tGk9lh+SpOAnekHOSCrcCg+SALleHH51nY3d/jaHjZu
J+IOp6jJd18rklT1ILm4KQ1EFoRRM+Ic7DmPSDdyhXeREWW1oIrDU3k5E8Qykbxu
4MEjyVAbFhjP/RyhWcuy7v7mNp00D8iO7/tJR8dPzg6AwWraGJ7W9XfM0SodjpRo
cERim6tgZXEiBSK0IynsCcLnFuNGNQl0lGvkcWJ1NEpk3dE7cQnBqRactgzbbHcU
aiUDQSwH+2u9Dibl+am9K6Y3P5liHtou4VzB1wgGEnhlfRdnH/ICdHJz7G3HU06f
A6NQ1gcrWBuuaK9VMqo9WlMB8DCOwKsfR2JwbSdSLTCZRv5/CF2M1UjjN5e0kXWG
RGs3ZKBc81Rf1ouAS29iufk2tFNVa1zmHK+MFFSpVl+cbm2l4/MO28zHp567O2Dw
atXO+0pF3lOkIauavhkndnnvaFffh/Jxc+lNiQRVSh2cHo5SWq3FkseSefcXzLiB
iWddyGbOAyJISGegm9Sl80gErEPT2cxWdogpnazIl9l0Dlezg26enDJRmuZwzF4y
8szPF7cPcZIngDFSLNhyKUUpTHph20cdP2pgqaLJQiKLwNN3QoLdwujO24juA6v6
aCY/Z2jUR80YuuM91BgJK9gOSzAz/h3pgpCyPkhulehtzkCVieILcQmsfiRVOAbn
9FM3KfbpfNSguaC47J5uMRsfcixtIPuOcuk5qUPwLkr6867bp0sK3at6XUQCBvDX
Krwr9H6lxex2cXXLne+Wlr21v7r8iN6wAj5zORTliwdt4twRdlUlD/Pp2+oF2ySe
PKf4pJ6O+y4SttdrCq+IujiH8oJh3Iyh7BQOp+nooAeF3rRe+sUCEegO2b1DUp0S
OTyJ1Cf1SaiJM4AnHLFVqD0y8yyK8Lp3bTjA3KRwIQO40Yb3dP6wm6jGE1KVPS5l
RLfWxA7UaoS64URHIxJu64khoTXGyPj6xWFX9IEjrtrFFMQ13yBZ9d0Uqn5sgnnt
0dTnD7s7j0oImRcJi0UMGZH7pyhoDu+TtXupWBPoXKDOpNYEwqpZl8MW2My87h0a
66zDzu8vf/DdL9bCO6tf+2C3lbaqTpY9ulnuInt+Qhu2ErNBqpzUZZsMjJywxnS6
ChkQIKmwZWkR3lHSVGt17gVoINHCN8zpVQH6tiF/vfqbu9KCHDB+TrTccNeuFZ+P
f9iVsKi3ikCtYfiAke1+uTSI2aDIIudSoq2HbNQtCB6hqmVvLJHkbCvEIFB0H82E
VQqV/e3ek0/ZpsV/fWj/Ztc11ELkH1lySaMFOG4w0Wqi2JLD3TYyArHwjXSRNyUp
QA2E8dNCEddp9o7V3fJV5Ku+80I4A92s6eGJRJwhwT8XVnCBTPdG6xpXZzlOgjYB
bytGs4/kFHEQKxBJURzi2UR7RNYd5wZH46r8f7drXcW3b/c9pYJoEDBgoVmHrDsa
F0tw5cvjhHnbiHzmL5KudnPnRnB3rbRbb4xNGBJiPS0MWbKay+jv9ePVnoWfaPVL
cokioWZ0P8JR+SGKLsuAKoiyB/NfIblN6xthn1ZnP9fu//1w9b9A4+ek/eYDdErY
GNO6GZMrxYK7nMyh9Ooimj01tXRtwQKBoDWGe7RvyI9paPGBwWLG9jkS+4E3WjFm
+0n0xUhOtyQeIOZ8oP25JIchhqWBoUCdGwhVCyeyg2X9JGyRapaClVfOSN9CpjJ4
e6WGxmdb8iq8Ot9sHj6GpmD7C8eYVnw2wl9TP+0L/rDmL8sj1V8mFMpG9CCn2Hkh
66h/VtE9aCFPhqzKKBIlx7V9C7I5Nn23OsC6ZmUFi19NWXg+UdOx4zJWW2mBS/Zw
jyfOAjzSH0n/yyGRvLZdn5lSsW5H1aGcm82f+NZ4GZdnvrd/kcdLH4aDsC6vgDuC
1u1ns0y8fqBQPcrS05VEyOrNU4euds8oWnlOk+yW8hS22fUkPxETJVr8LKhruEML
zHs3iPFft6TlW6twPoZoSloZJd/bmn1tb8N0a2+eNgvGiWJQDh8bNynUicuwC9tB
BFN7EhNmQ0VX/3EOf3RaBKnnH4cjRSjXhIx3kqeYor/9+6euoQhCKhUw/sib5oBR
qaOse8s5QOxGVsMjkC0YXSXepO/CehXs3hTrXYc21QQHvDt+wvZLq1Bgdxh/14CS
PA2lOZmKDLg2tHXbfc1ZJKuQEeDHpY+PG5Vssp2Z9QED2U8lerHR+hQkqr61zzWp
AKp9dlnYQI2TXj7wOePJmp3Q2sizbmj+cNMB7ktx3khxQJyQKsEa1Sur1yhuIQ38
BJoofuFtDbSZ9iaOU4rM5bw6AuWpv9sCm2tYtCSKhfhMTmCUze3wWuR6b+Ap2f2C
C6vvit1X41R2S3nWNIEjSByn7DIoLwc5jUEQUOYuTuZv93ZfgwPjAeoK7DegkJE0
ngkP0y240HLGSrvEuzSAhdhma5DofG5SFCV4N93j1F2CPvpKImn/85ipt00cjDSN
qbSrvnyBmlyZMP1Q/LE4d7xuvixrdWY0wcMp5JRV1bDwa9HMEHyJ5H8PVcP8gl3x
LRpw/UaUIkkWudDzV27shYKK0LWVjccxZdTNKPg4idBN6mhJWLiHG6SJSxb8+nNT
chYbAm0tkAvnQxLRtTIA9uuwmDpvld9VTPS5rLIS/ZEPEexDs4NOJRqTxbQeI0Vz
bLQXvg1KDsmW33u1ZvYKQouACSJw014iuNI14QWdwEApB7GTPzvv/19hVf7Yq9Ki
nJAOjuPXgzg2T9nKFT+wfDCGSPmR0bwDdjusaHiJ+UOearyDEHCYEAL1b5eZSEbs
QcFzpjsHZOqaMZY4JVBn7I9Bhc9+GI9nZOIA36JnHtkIsUdJ921Hxq+N3OBWHWz+
JIz+JLfUI+Mi9g4WqRjw4Vl0BvAiCExu5pGOn21KOxHKu5tpGvSceyfGpSNLwnQu
gmAgUIlV/1R/RfuIrUL41mT06kVOusO0HpsectMz9JjGN5/kl/U4IEwfFZBl9eEa
iMl4hDIU4W905EsH8BRYlA+OPtE7TdJ6xBpw0XQHFtGivMwYqImXBs/SN8JUzW0B
k0V14zaETJyNdy26jALAx3L0mblYwz5N0q8WoaWz4QWafWxloIdKNrvKHHQOV7Fv
KLMKejtKjSIidKNME0oX03D40pYLXK3fPABfDf+7beid4MGTKkS/CsN4x88N2r5X
lKPolOICfvBy280nCNpyziAErfYjN/+OC0rtC9/DO2jjW++xxvyJDvNjrrzCzu5Z
d72Xvej51hGvPtUmZXSjfLeksDM6NjMSCln4FkEWlKu5gs/bi+plGMT0FljrLsvi
XsYHDTNuZmykrvCXIt4p1dDx7gjR05LVAtaY2rAUYbbJACtY85xT+6lAONOuEz5a
NaRZXNodbOAhNTCZrZJzatXGLNJ7M2gKnTMljxJTJCtN+UKoTpYJJA/3vTxVyeRP
rMogonMA0b3mODenq6LBLl6m+HCK5RgrT+ZIfPJIg2a7P07vG61y+3pD9ofrjslD
ULkp/oaVSHnZcTYJW0xEP8Lb/bn78dmSGe2dNMpKFnLEY1G0IKEfnmJ6uzmC4UZD
s4V4OW+8hGku9FxN49GFWlW0jOo7vYPW1qcfyzxDF3ZT7VD03vlqhGjeqnqDJ4Un
cfQYOhmRmSOJukzUm/ZvT0jVeO8zoGN+vaYkyaIeQBA0WpSLfR0rShXnoXBqP+KF
ld+XJN0PRK1GkggkVzYdChgk3FALkNE6ow3X4WEeglbqERLmOQnbPUKox3Btrd7n
0dTt3hFs7j2e+z1JMW7MHSUjfbeI+V8Z1Y22dOOVG6x5wKXTdXLbJe5tPojon314
mqVZSJKf3zY4z2P/xUjfD9rDnMDLz+cTVlBwCvE4RjTeYMNH3RoFLUSBKLNw/E+1
e10V3SeFsDMmOyGX2AFKDDFr8aJdskWXjm5FNNwc9oZzccS83Z6IwjJrjUWo0txF
Ze3xAlk4mwvhK0j9SeLqg6+xeMLVkl3Ou81bRL2yGxIFNJG1GkDVkskZQGqOA5A4
/Hpz2AyyhDc+hQpYes0INhXumBfCAoO9PKXR5zVtR9cVh/u2QsxPg/+70bLU7OT2
5X/cZAq21e2++SyvcJKrTZbsQfO/IZU8VGkHyl8IKKXQExQuovoZGM1E/T7nTpo7
2dkPX4MgB/8Qb4B9CRZSF03eFjvJPdqFUemZAMYvmJOG9HExKC2qMavZjXDsg10n
f+nMWPTtDQ7jVzRWQS4W/rI9WsIDPazqAvWURRrnZoIfAKdGJk7OygTDyDrKJZy1
nsTWK0rtmxxkMZ8qVr1JE9My/yuKcw+3lpbbtfypXolVUEzzVtRiOb2PwUkomWxX
M64/lJnRiIrwKG3IFSoItDE2WfGgKtvX5gSmJ+vNOQa8cRDIaIIGIjuciZOw8Ji3
etgD5e9Da6B3r5gmFQBHruhJrvOHzU2CWGoXFwthM2mYP3TjUxmYtda43/HDjDpn
PIQoHJ3RXyY1NTJtUQZuMCI9UhHKAxb8eqeOig+JbKtIFDgGleoxvepteAYaEPgZ
mavbrQYMxX01IEVUqJQxsthoSb74VZmebXP1y51Ll/Gavo2P8F2Sud4D1rqLdjNw
tGh+aIrtrytKFN9zsVDMjsdl9tUSJbxLdE6ORGSD2t1+YGVrPkLbyJsyNneWlb8l
9Bfy9v4LwZ5n8zI11bF8fLepN20G5IOlpwtls1Its7o+WjIXmn+jPhQhWUT/dU9C
yzd/6HXPdjU4HQs5uNU9EbsomHf4A55oQ3/q7rrQClxIbOdvUmMLK0FMxFnmyXlg
aBUUdsj76ndHlu+KXf2BpU4yv8E79/cKzfL5SISbEkE1q5B+Ssc1n7QHgoWt6AuY
mWQSaxbxTFfNbqCDB8rcXPK5BYZCfxAqiQtjcgP5X2D6ZOjy8Q3edTp56/d6vdaj
CEPVRpF+n+XnsRKWLfwatBwhUjw54m/yKfPnAC/QRoOKjgaNv1PF1A5RKflP1fbe
TfzmgIgyt14YTZ0uS3cmQS3dNCpdxMHSJBlr5sxbTbazGQTA8T3pinhGD96LMlLt
t8YD+pBheKTUEiaWP2J0SVI8CcAsN8pwWb8gkp8RkEPlcFKfy/zu3NOBO9643ZMX
ZoymPL6po3OyvHsVOB/WyIRL8vbg0lcYNgsvkYl8q6hjNrVSbKmWh7GQ233gpQgg
leR80Zm+GLmjVq/RjNhxk6oICk/uNRStkDGpowmbfG0LW947bEXsUm/LbmwmN0Qv
B62lfhgXdSDFlLEXAsT9aBXijSMedru1XhBdQfV2mc8zBKPKNMRJmNldVd6N1kFk
PXukG0wdTSE2EDBvdcTvGP06BKK696vj/Cc5u+tTjIEJc5Ah7aqQzrABbBa8kc8g
oS2Klb3pK51AhU3gplzUyNvT5tsOilFG+AafE9nsjrqv7JwIh+JrrVjVKCbejtO3
yGMX3xVuuWNYM/qnRuuVDCnSvD0irmzpAwc6Hm5lBFD4XdpJUAQ62b12NTu/pD5E
IbDqEl76zL3ef1IBoSOdXQzS/HiwsKu6r6ugi+1JE4CzPsACQths6IOgYW4RmMni
KzZD1RMA7TpgIFavAxSTKGTrXrwp8YlWE3HafoHhfYmE4GCnDjyh6/wUsYQITY7o
C61WqWa+VWbhRI6LMIlm16hCxaYIlTTvwDJR5liehTVRsB/0e4H8GALiqtCWUmDz
WSa8H3bmuBwP/pNlqdk2JMTm4PF4IBuAD2kHYtnEG0lopb7UtucjQo4qqWePD/FI
yRml/+51m82zsssr4/mN32lz/VpWAe7Fs3t4trPfXWmkGcJGLF63cA4rB+owESng
FsCAnxhJhiWIDqdovGT00KPxIdv8uOhToTnAtfGVebUD84XfJYrTqoYIwfuDOlZT
asy9g0w3ve3KHuA81rCWFppk5EiCu75PX6SS7Hm0jLESkOYk8ScQqyGVbZToEIcY
FjkGq0U+0SspQAxYrtuiOGofHPTnXNi+ybeA7ubJbYLQ+7gL+ZUYM5ldZXhEpVI0
8uyZb5aR3IHclHHIEEu2ynOAmiJD1CwOjmXUP/SlCa2+bBZnsXDDzQdVvPdQktze
ZE+EKOO6bOXFk2vDBthV2ScotsmT3YNJbzOfwqBdZfA3wEIuA2/bTwOFAlQiqFvW
XMmI5u2rUu5qOsEsrUwxNOmoL29n0g3a8jUj3/05N1H6cXxuqwezMjyZBn3KcSpX
RPECBKteSGtNgvuZ2pZkQBf1H0GVSF4FlljzRfd6IiTeVYRH83pIG6t+2ErDKQCi
hnMOWRLEa7Jh1068bfY8UUNgwTX67X/cFZZk6TeoU/kvU2yFZPsjzohOqd2wuw/U
1kJRLhoNQKe//az3b4U++OB8DGNUzmhOvYgWcu40V6zRhBmdr1ubpx8iulTdguCd
tFonC4EXjNE5UOSGl9EwZ37JMg3nSNssskF482RNXbMHe4kqyFtIOktSsvNl/SB0
JiBwaLPb8YgyLwvi4El1ZGuznGmOzoF4UNTVcPAf8UE0tu2J5tXNXRZYI0rHsRem
YLuethTAZaAA1YzPS+e7x8S3INxKXTG6+iFzEVJqtS0we1GOGLVA/uhxIc0fgfe/
9ZfaKD96XAVxTLCXoz02k9SAUUh7PRb8CE0pE8KNTEA+vTaKqhgc1Ii//uAgdx6g
c6n7yMDmzG2aj6fvDZZNBvKACmCo38diJUKajbyCmHewt6SrF2EZVwL4iKdslgP9
QZsJ5saUUtUmPc7RomHi0MqcCP199xZrJRsYC2O1DrEfaPKgf+BOYMv09tRPecVi
C92cJLJ7HhVCRECKunK27BrU/jZizQgsgZCh+mfpkOUkfZCFzEbjmd125l+ucwKV
CYgmb4ABVeDunC7VmoTBJbzWEX0EpNg5Y3gVxfFKiHzLo/ebB2AK6BDJCEV24K8h
J4WTVqZkWRiumoAC4NM/plsEupPHDC3h6PYU604FQHSh1RsPsN9ca/unWsecSlqh
ETT7mDrKo0V9yfNr9gJ86LB9IFTxw+s3oJG+mMvQK7VxXEKpycIcnm41U23naZ8Z
X5z7KPF5F07W/5Qnxeb9Ob19QCPWSZ+urT+P0MPVivEh+Ulldu2o8oI/15OxVfB9
kCPemOIkeYDmpcmyEuNAXvpi+shDeQYALkE99au1PfrmQpA51mHCn/WoUJ6QjjL7
pZn8bH8OXtEqpbw3D12Z/dWC+0AD457yXgJ/AzlfsK3n8xOf/9VLDtOJOh3DSGcF
4vvE/c5eh71nSPT4QvaXBuzBaORIxEa5E+nEjXLCwUoEztSSCEjJScaTZ1I2KAXQ
dagh6znJYA9jV3DXX7ADa20iyMbvZ6+O2D4HpJuL4GixmrC7ckrEUmInUnMT+4gy
0OKWDpO4669sF8HZvJNRB4XS67+nFMpjQvhg990nGbXxOB+IeQwAOaWzm5u8+aU4
HywXEjKaXWf3qJg4Ae3p1wLeHa8gJ7pB2mBbrpsLm4oH2C0AHT8s3ZMMVyKm7rYs
wGxTdyArjvgMk9rFtcSPb9/7jid3CssbaVZWtnsp0FyxKuzF0W62Jb//g0k8ndSJ
qVPtYXcGaAWifIqQanMY6CI0SOMIrCa+0TTEa90d/w9Osp5z8ys9I6IhhPV1jzLJ
k6MApamv7azUtyxpnA/nV1/hNOVCfxF8+g3MnXVQU8J5vmYpRmVvUtUExYdDMQeD
skGTOoi7adILOsta4cVfw/F2CY3ma7uBNC4OTEXN5ATRYkzbfWSlPMlKC6NKuMtf
cr8rg3gpuzjJNILgc/7Wimod88tDyvBrKRXOasJCkFM1r2RBIM5wh3+11nqp9mXD
C+ujZc5dt8INV420sumJP7T8Jm4NX2fSxXuhL1958C7wlKLs7D+SsigCSWsBu1xl
zXanZ74tD2tK0+WDJZHiqOGB8yUECBI1i+/8Kls4aa4IWRKUCO3OVSpfpSKho1lP
pyr5krvXS1Anrxo0zkYxNJ/TDApd53WEuhKVCT2tWnX9zfQraVTsbqyHMFQJ6A8/
yVIXaNAwXbd+3HvpYkzerDKlCDVLFjxYaVurWqU7x/lGySAWl6Dw5c9DfbJur4Cp
bnlF1YGmNCKHK1hTd7ad/vs7DovFjYVqa4i/3ROXQemabbS/b82XDOzO8u5YSVij
qe6MRsiRWNVXTzrjZHGj34CHOF081ZASVAi+rDUyXl35ePS2UzSFTKp2cYw4YfU5
uo8x6ZYX65I9giPKWLKCDcq/ebyGTslhOzsdfrRUgCzwvTW50CbOEJb9qzntCWc9
LuFxmPl8e33z49YqKVL9r071aNxcXgTb0G7EJiUgxspS/TAGNAdJTScaBmW95hJ1
Ns2537T/ngcSFHEzWUBNoXoui6jcBStlaViG9/6tGL+Mn2gP39XHXt8Z5BIqaJm7
GYHjtvSs8W7a5Vn+ZPdoNdUW913u7Shl+4nFpsZJkyllf9sp3AUV3bI0q/6JHnzD
JBQlPVhodVpKaB5lznme4Si1SD1w2FjwZSgwIEszp4Gtf/K0nUUC4Mkvjnor6fFj
fbN2rnQu22ptblEJCOnYYHuTiL1QO5EGRQkgxMGXEi4SQj5gl3p/rvcP7Q2JEbDY
GCdbcwa/Dq+0eF90F44bV0elMbJQYps4Kj/x/+Lin1u3XcjU14lXZe/h9OWuBUjp
Ra8MT+NZk4YeoZYSvCulEcdrrPXLOiunE8KoUtyhB0ldEk2fvFy9zkhoJ9D7AsIB
qZZ/A72q0Z2eKSQ1XweLfHONVMNpXRZYubUB4StY9b7B/enM0NmKplvoReTWSLWl
TJu461srFSckkP8LGD7/4CP81rX7UVPQ7lDQNUe/EHVvY/iwk1YmPTTcA7DknX5y
2hhJKSxyR6cTCuN62ZbHtB/vCI50y/kEWyn8GwP1gzhzHbP1qyJXwG4vDcycCJOI
NxAeUJUeEP9jXWX+P7XUOuW6r/PUv5LtYjt0BXRURFibMp8pd6IP8kNcHthC8R8O
Q37wBgyUF8RHdAf0gup5iATy6VVHwTF7OQuh1s+dgky3pc0blMjyAQD7GTL7IMEh
qZ7ppw4QOSxcOJCMhMRtu0Q9q6RoHbOaqGkXmwN+OyU1be1G+WGUgE3Mc+GSmvp6
lO7ryB5++JA7R3Nok7bKCRIB8HwthfksisdPgSlSi1+Dzh5dh6dpXrfcWtNW58Zt
nCuhS2pL0yCkO0fuNpxFc2daiNdqPTVBABSeGFQ4GxwTSWuWyQ8BEGxGPi6pP59t
7L63xzJKp2+85i7RVTkum52RA6/q5ghlLD+Z7MmbimzUHR08C7AEDkmahHMetLVW
BWaU2KhE08MwqM0yl5w9dPkX5F/9t88JcEi/JlEClxd+0cQxMhKMrQR9JB1G9f7d
K7vB57fDGeUgogLDySsWsPMkS9MD5VEow7hSIScKMiG6y4uY3vBDnFnMxjUpwI3q
+j/SNtSZI41ZEVvfBxGIa7GrzZPgFUsk4RhghsCxjDfbWR8dxA8j5uOC2Mz6dseL
sN6becOfMpK6dh+11Os9bgrfxrzA+hPYAzmaJuyd38r1yIXlPXSfOI3Cp0fT2LMv
N4fVPAkb3eGfr3Cik29mmXi5+tOGPqvEuI5vnqn/iaT+1jkQK0nzjs9/bwaGEH1y
+ljJqoNYHiVt+6MFN+QzCHrNDzlT5c99I7LS83kMnWX3eusj8D2109C5CQfa+05k
t7KELxHuljN/iZ9tJU8VXvoODDadqX9uvrrJkEl01rexQ9Uaeae5XntFJj1e0Smn
+E/6rH9Rc3nbp2yGZjwwIjyXYF+YTJDmEtTVj7Vf3u9xWchgW7ZJnZCeN6Muxy5B
PSCXNB3RHL50E0lcOmoNh9zLJ28beVZ9PSj/oystSq10zyQKx/VUnSdbLxCnSeCj
twhrzrRbtri+GqS/PNvlRyx138JLBsZNyNgB5wVCVWoVtU7tzkCmDi1r9r5Eaiiu
GcD+l8VvuzNwnGt8oybpYSiLUySGckSBjdXqLGDal0vLkv0ap6jaJfUmXSx8md7A
2inSjLJ6JBO269OhtmKKJap+mIfAtm1kpsWfqtkTuG+kXpcfckUuqCdxEDdWsfDa
qRpOp90SDUkodgEGC3371qzNgvklx6ehnLLz2f4OtAhsB3ir32Bc7NGSNghZFkon
x8C9rv+LCSneutZ5qSe+4u77wyRFljPQujm42OCTMFuCC3ejcnvvEVjNII82VRKO
UhtZhS9ZjNfdBb0atEaQstN1QVN155b3NtuVX5BAENH/1BTr/XbtQXBadH/KgE1n
V987rr7YyTHIjTay1NzP8Iy4aK0KlBFOJzz4vjLshPA0dO/Hy2zQRFsCwGWX4xT1
bGFHM3PzHuYXw7f+lb0H/zTBZcUTyfoyJfqv2WQi81sI5q8OOiS3rmLqNuS/77f0
Yylw5zFLXOUoM4urhoYwE2PhSTdYlrhGLVGmD1GLj5P33z5n0jIUaNDV907gTZQ1
kCNYOOtMSLw7l8p4/7cnM7gFgn/87FNMx9EMkqlaOtiN0Ic9N9oXqb9I/u5Twuy9
F9SvhjwXeK6D8XK2sskRbZIVWatCDWzbZbPYD55aj7qJ+HJEgMeS42XyjINUR16T
zJxgKE9Ob6+7dAHK3i4fySWbLMEWpePM7G1iN6eLMMlQ6mkVdWnsseQ7Bn/nPmSD
83e3mg+Vd/xnpxU3TWdLoU7QKc/JYf4WME/ZbQdvTB9pT6q2WpZIL1Y3poSGe2Mv
fBSMfSpIWaxuQRmcg94QGc+vzlnrk3KG6GobEWxHZwbKjSokwK0O+wjbx4+K5Odw
ZjUWZBq7KLjnUZFMuKESvISOapcYNsF5hzFl4U37ZJlZY+Y0HRZ3sHRCM1JnXV1Q
qigpODFmPAx5dziRo39S5g751aRMXcjIwk5kamuMJJ0UdbFCLq28IJPQfMhFaMpJ
3L2yctU4HojSzCl/6llaQTlbqm1UFrCWMKStvSegirhi4Jj3HQFxPzrBTE5/55Db
tJDzvSM7mk7n6ygrwiIttl0GqQP5YeLnR2+Cw5uqZJP7VdtjoKBHORfW8DlfDS9A
z2rwgDk9Imx2qgH5th33GbaUayElq0WX8Jg95PdSfvhrMg9OS9fFnWmbuhlxNN+N
j+I503yFaKNR96GmdkaYzq5GbfWVGhkRXIjQv40KvNE+CvgLZJYvLaX29XoPUCmK
w4R4hTFV7CY6vAWQ7qZkyItJ+qT6IcsFoaOVhCNcwpTjaV8sNcwujGVQvK6U1iw5
h51qArnTMOPXMwKsCiADA+tXvFPgUMRR/XfbpN1QWmHKDeBh6YdRjNo+kuqaQtrJ
cmti/IxHIzV4lEbfcPENf767Bh3DYpd6OStWJGX5Fg/0h1gZthh/Ae2DLKqAIq2Q
K2Xh70ejznMTdpPpBPknljCSYgU1SVXJI0nNJ+LzYkGrRGqN4ANfpKfO+DRCqUp+
Orwbi7jqEpLl++bUQdqmJccGENfpRw3eAcMcsh6Lu7nkZpw42kZ74caHaFc1szd1
RyePtulIvXThdpHUmv8PUEs4lwIFejCG6v3DkuWysfKZgn4iZsT6O5uxtv2CsamK
RA/EYMHpyYsffUZuBnZVChxDFNddDT56A20zgc4H4NqD8ln0hGN3A+60FPlQfFgs
svkB1LqLGarYSQUXKhSQbmEOxVqtVpU3rD6fr1rW1me/Lw2M3vdRVupDBcv6iDuk
odzaUeo2/xx8O4C86NBt11iImNx2AfL3s+X7SpYg4rMlSVy6Av+P0ymgrSi/zlg3
6+DYkZiAHU6fjvSKa7qA01x14iuXp9JjPSXnlS+S9X3jft+EG5jg7wvZVV8MaFzf
ubVEaPOednXXgGRvWwQSWERXpL1IumQimINf3g8sR8VzwczE6l9lV8jHvm1cvOS8
qbTrfsOVHdAcCCgMQb0EmcXM5ZBn0Ul3NllpBsHt+o8eMNh7NE2AfOLi5JeCTizi
Fe5Q8OTQxW0b/gplegQbkGW8nQLqxwuzXdD24yRdWn02jEN/3XsRELPHTbJl+3hS
FaJJAPYoGKfMpB3HyRm3bZiDgb6xG4G0UBeV0Kzn0bPOOPKkWmFAcVE7uPhABzPf
Fg2yo8HyyZjAc8s7j6Hen3xNVS8TjYZjxj56a0W4SsZWO2jOfxMMHLhBAvfVeJGl
gaRi9GlzWY3LIFv/jymUcxmySghQGE01jZxFcCftyiTtpq+TkeIF9Brty3C/fKrN
epLA2E9flxN7eJNIxy8uXv4MNEY4Fl7UWtH17eGe6V0=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYrLhHwjE+Ay+RjrmYAdTTBt6UJnpm8tifxoE6w7CAatWAG7yhcBkUh8SQkfqSBL
Z0XcJZahSuRsUYdNv2PGPaDeEfaRCYVmEH5Qj0+e80HRCI6VurJ6e9judTUYiMLy
kc4LAqrRnADOuuUtWM2okbzQxDja1e8jh+RcVEz+8iGKUFqOwG1i0E0zCf26r+Hr
fOD1oYoCgSU9QxM+PTICV2qms66Om4t85sW60LDhbWPvniACkcRkkG2tj2mNpi/c
Qyuh7o2iv/b1US1mZTtfWOoBJBNRwZDCFahE+7qEv3Xe4kOR7GjhlgJVkqAr6dtT
R9zxtbnchNWMLfoB168bbgGkNzMhE48HOhVfd4YrYIe+Mb8eXNBm1y5JpNCedzYY
COSuAQqbrvZN/dt6aOkSlSUSvnR77JHtXqH8pM9vrIvETgCNRpE7qzCTQkdxLTgG
bOvL/SUFS77Z3tzyTQLfcHZol5f+TOhyk6ECcK1H8wk3nA0d1xRuW7VGDvDBTyfL
MTrkEJVk2J5rz9TrXWfuNzT4zstDP1W0XvTq2IHfECrGPiEQnXEgExQRYJ0PtdnS
dxXIpH/KQuKEl0WDeil44IjB96MXPg/C7k7OTN0I3wGqLkLVzkhhBdzQyREeO5PZ
thN5CzIrW8QupE91mSjDlUucBYb4uGagVSzqjrRNR/Q2oG39aGIIxw39tzpi2kMU
rLlbh0+jgiw8mdzzT8qWwSGa5inEDwxi/JQwOiAYIIozoVvo1CYdPUdbYw6yccD0
4DurZKp531nQOuBXkGDgRw==
`protect END_PROTECTED

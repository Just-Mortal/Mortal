`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Am82ldHR0zKE4uiOLheCGqf/PUUtEtFdXEHZ8OaFOJx6tPek9mEUJYxwfvFRwHXd
SlPMvf1K/X/hXaO08A7Ild4CrUK8TvVIFy3bUqHsEZrw78qjit6wHS8opBw1AvQa
u64Scah9CK0U3bM3Fgp+Ec4QHFWoSL5RoWuknKwhv13RHyfXICdJkK//zwpxW1H/
pyshUF5pEDLJxilx7Arp61BxnB8Ux8sxncCfFAERzDhIecTpVuVCw7iBhf7YoLGY
10DiCzgq+H8sljNlysYh2krHdnetwG/SB09J5E18LDXsTPOzOrCl50HdSFxEsFNQ
PGQECV3ESlgHv5JVRUbe6YfBNJGGyhCF92XoDcdJmp2YX0Ow84pEEIvU0Z1Xu5FF
y1CmM9CkVNaSyDPJoBoViB6x/JcnQzAWc0dvX6vDpKGsQ2zxVJc+c8j9aN+IOUOn
70QvxhscgDMXd6QBh/ZN1qohc+7hm9vlxXc02yvG/1yJ4/xrc3EXIzM5zITSAVJK
b1bJdHklUE3pcPPT+czWNWp/lCC2ynAdTuwbLjiXO9e6ZAWGF9stS5hHccGs+dW4
fHIh3ToCELVNojPcUqTjdCNupWTg6S3zlVtQpsBvneLrK6rG8AC8t0buedZtLNUu
k4UzT8foM37n+UXpRJP9MawyQRn/uXEICeZjekKAMsrBe0Q1ZqAhk+FjZR+u+V5S
PfDbP6rs3+61yApIo8KQ/kImlaA6O3qmFmX/KnfDkmSIAr5+iGPJQrNhO9KWoQcZ
aJhO7XGA/zVGGh2SxAOzWqAi6k/Zx/leOPwJY2VKu5DdT8meJxvjnOEfM3OeJsUq
xJGhsf9lGy/aZFAZi41Povh+cdCS+aCAiL9bw3nAOCxtzG1ZcB+xySbdrUGd3ffc
RgpF0GP5hP70FzNx1MDS5sS6cTushZVcE1OBDvXIZoM=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
whHGnoIeV0Py5uvauMfjfgc2cKy2OnNkwC+cWjL6j7MTl0vje4emKb0MFoeHVCWC
7cGIkAw1iUkC4auIhDFj8sdBVTsuHC6Mp0UphM//JbVUc16Ck96EptAhnza+RK+m
zJcu9IkvaArRACB/5AP1F50JmSt1FktgCcXlxo387h2lIKK504HzpGKcZslreEii
8aXB4zGiVZiINOUR4uQltZgaluP1btUwfrcdPh1NhotDoK8DVdDQE3xB8FQiw/Q2
pFwY92eJPI2bKVS+5oVBBvcdg516idwWrR/wN6dHJ/K6+Z48MBV+zLN63MRBEX8T
IoVGXPt3ChCcC8OobvlmdndgRsdtEGBLtr+V2D11OQKEXBPovB1sCPL99F++LQc6
eLb88Qwi3lFHW9c2KPlPK6MkVmC/6qj3blqBb/aMhGgyQZ79iil+XtUQdAkQZSt+
YDHcudFkUar8bM9g88rPHN19/LTr39UBICn026f/DclSUi7dgs87b9ZhEdPcTbv/
IZagx6XH0jH9yGCuBOATAwF6/6O0JPQnSaFC4dntqMdzrLBIno/7GK0+f3UYCE0S
`protect END_PROTECTED

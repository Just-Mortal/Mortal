`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Ldm4JcYGoNGVLXQUAnOZt/vpkOEecHXWR8SFiyh+/pHaCQRSs/jFRgltJBuxWX1
P1fWnpi6AJb0qGu88bc7KufjTHFmqcE3UKHx250nv3xz4FndxIeJyV1ZONP2DJdh
icrl+y2Y+TuL3qgcCpAmy1V9upj+ByNl+i1ifkETzLEqnAmeXNUg5n18tDMg2G/D
tRerUNKD8QqZSIY9JGVjbOB/hznRZyLvUX/TMNgeCBAViicVKfOR0KbgGK5shOz3
4SxHW88PSqWWw74H1KcT6tR74suVLSmm8FC/Q28BMX81vcYJPI/xprHCaRo1P3zu
08QUAmHrblT/4GLg/eQSw97X53smYmPrsiIJx/8kzFgKgutbiyNbqOtNgI0+YDxR
9qF+Vx/rP59vuXke3VlB+wIIVqA4YW68ixpNC+wEZDKxEuwB1Os8xkAGZMPPdkYN
5s7Gb6NHGy9ieLR0LeeTUvQSf8QAtdDXeYFrlXrEzlhAHoO01MwVG6OFA9f0Bd2Z
tRATg5bDzzWiNpE7jPjqcIf2fYGpvzwDr8Uh1qA713/ma7+5Lxo/hR6HyL7GzC6J
nX0Q6w5XobuUyrsRL0fRJc5HWLHlA4qBd0rXe6ipLpkCFmkiXHS7hleiMVC4S4AX
ghHQ91TqBD9I1ZsAmkUZu8kjP4ML7Ot5/5Ggz/xwXTtB2dRbJjtjS+fYIUEimGZ2
u1PpfTnvMIzTi1c+JFg1LCUJH90X12ArYksCzX3I+Fo0LjS0baS2R6821Bzm0RCs
ggElC78A/H5+k5O6qOIzuB4BNPHoMgpdFJjLDonbyj6If1cfzwO6FjO2rDZiOh+t
WGaqWL8C0m57xKpwsCnbk3l+Lhrt92iPVJj7QE8zBHlCrxgNfWgLlbXPLYr7xO2y
mFRXBUf0Weqfz8FSBj6BUOfeEKI+H7X3w9h7HKhmcVfVYNmGb3/9xIgSMrmsl7KN
QK0eKv/nC9o1jVTdphegrpcIa2NfcCe+GeQpmZY7cbRqq5QzGrpedkZT+1QJtY2m
sMhs15AIUyAmqVNEd0p5GJ7fX9TTr6/1i/TSMkMd10hDKxDKgKsizT2+Nd+Yi5xR
oxvEh74NJ9o3NL81H4GWl//qjrFNfT0J5hffR3+QXSyMeheB/GdRLJ9xF8Qav1TX
xYvfw5eGsAS0rTe7Pn867+/Qkd5Ai5iYdedK/jBt3CUmEZ1sgQpYwfxQV41KiD3p
`protect END_PROTECTED

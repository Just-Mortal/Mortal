`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcWPju1wmv5XGRAAR6O23DcwJrzBcTCfXx/11r/othknwc5pahp2EGUCzFtUlMo1
IX1UJS3waZJk6qGXYr5CV4UTtt0q8chW+6CwH/V/EwriYo9LHzzcCWuFP1yskz+v
LZpTYYOUYEMij10zYSEUPOfz1WdCKU6EsFKBw1mARaYTyz/nLuzaZBbF33SgAZiY
CAgVQ6plYnOxjy/NCjRCw0cx22Z2vMAEGVsT0N7I41upHe778fNYYyyStCu58j/l
LmTgAxZkiee/DG6SPey4VDmO/zZnc8DtFW71KctMwIRUFzoQUBladY21eBl10K6O
8P0IgaeTbXAQkyJcij2uoLPrh9+SC8mEidpCvtbDQU1JTNUmmMXK6axDwnz1BQKN
kERUCvVGUBrqpz5U1JFoh7+oa3G9AZQY47xVfCk9+VgucsSXV1gqonoIeJ1dSZl4
gl0VpNWwZLQ9XuaoBS4tc1K3EefKDqq7boVre6B6ec4NPf8Te8xDJ1FHGnOp9Olz
tqpBVrrFCX6shVepqiI9Ytujh486z+K+BbU80Y5sfRhDyXxBQuO2rxsxmhx58G4v
JTBV/YMG2WOpn7aViKNs6WH2a8wUtU18kMKLHITR4+3lY/Tq75tDbeCHrW4BNY9P
IQjbweSmZ0KVB2KvYxx8Ug==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
keC2rom9xsjgWinVASNuKlKc6QcNaPFDpRmuslf4/l9ygomeRI1kP06fTSE22Uec
DRJHqJIyURL4ZCiOYuOT/6wY3mrn7pYcvDJ6jiOCaiC9iyRXz3RfID2c+HPI6/Ax
mXxfPQHE/xOuV6xEsbp4Mq6LwKRWJrc5g7Nf+6FoeQmV7t9793pB/x6J2lkKJxjD
3/681Uqdq7Iar+0mSYrbjuVBjPCasWCXGxw9N9+uwkR6JdsjY7Feu7u/eLEn/bCQ
VoF6Ngo+MAsoX+WUOOeZ7RpFudDOQq6cIAyxdeSvPibjLft+TVshs8Ecw8E13CX3
Gu2/utG3M9Dyeeocfac4ImL2w7egcesAPenzuV8a4lMudbMR5syMHJKN4ICDuCfL
1NTdaYHGtyiTK0IDci9bKmQcu3HlN838sEVnh+ttGZjwBtm56MxAPWZIM/M9J0Yi
sZzT/uM1+11bKqlEqwWipR2F05jaUdGHVdWRFJ+HHaWp0rmJJILiGDeilvvPAvuY
1firCkyKpJDacA16ch78J3IrVxodOEXvcTYhTuUnmjwcpAQyI0DKVeuf5KO4YRTR
n9RmNbtz7HYj30GJARR72wLc2Qpt1jMoTGdhGtbDtRU0cfODEJN7qN/IfMP7AREz
B/g/3NscoYqaIiMG+xb7ZxbbxGf9GzL/Z+hzUFOZ9M05eboo77O51zMaG2ZUSoh3
pi7wUTHjrkDHiXTbzFNFjLhKHiC8orQWHzmr41BX2m1WLlG8T6q1DKV9n+YIXb1/
VpOJkr76psAVBx8Nxs0moxtNGVwzkBkcWOgkS7BQjL9UHH917OoLGG1kckwnTEpJ
ZYFI/YyxYq7lpnJUDgsOQa9gFLMixxNQw3QvMAMRBg7s50/VbXi4V7xS3uUNMbW5
10cZo9CfGbbQ4LDxu6wbzbeF4FkgfvLkruVN/z8UfWTY2rBGzxLecGcpmySvFsvK
gffqEXUgst555yU0ZWpBPO8iGjJbtu02qkxSHJWnq/vjBac3pcwO2PCPQPPaIJAD
w/m3dKfxCfR5lazyB65OGrwQb5xMGAB2GLp38blBiKxFoMXdD1Srm3buyEtEyQJh
93buGLrvFGNA+Emt1ljP9ufNu6pvHH5oaBuGpwgMgYpYQKONJQ9BO0uGx3cJdzSE
B06lVsx0JMmxPk34EF0LzglBzMp+z3jcrqwAhNq6znOcXKFvBcnkwGyI33Cy0KU3
hsWdap6JUYF1kXapYMVELl9+4PQ+s/OLK7hzQQjTILTWuERi25nfapOG/ZzSnZNi
RcA4+FrX/k4aldxWAtd+7AA6PYlYr82Z2xPHqekNoAEKOR6qioCkOTz6UIxCU/xd
6NdGTPzugtRTTXcyhpJ4GpKlJ8Ul/cuzm+C0N0zupJUlv6sdx45EFMY9+nLv/CnU
ry2s15ZTkRxnvoPMFxTDVWd77J+ll1O16IcWy4GHI4dTpyQkSX6TpBf8Ujc7k9+t
Lb+Yur6Bi5wyT1SaHtc1fEwLE8HcM4SEa6uRvp41txUfsihrzZE6KWo0I+KBtZ0d
A/fHHBGWSPTdZc+88BWfhQ29D5iZ9nDRSqx2cMTgilP669Oxta+suydUYj8aiAWv
4KL4feTGGrOKpf5xkaROuj+gFgktoIyvznZ3xv/tEjQ9TIUHPUreuZVNQfKOB1Cb
oS4+/UUG1AyfO5gU1E6qyNXMz08z6AuueDGQ5Te4wK2VP8mJwQnGZ3lyb7P0Fylk
6b/iL4y7SOhsmx/FcnMVs5G5QBEmtSb1uLJXujkd4WmdpSRIGR7R/reFgeC++eaS
gPvdazgKdSrxVgILZQt+G5ouESOz7i1cJGSKtUk3dxETjF0noUH56P0CkGTdIgRu
7Kh+MREZ3bUyjdt7GSlzZHPWoyReabRj56aPzS/deWmvxBw/sGkzlKn7K49u8lee
ZjqZ2PCnO3LAFcytXaxl8ftiSQvT+p3g4BUBe/DIvijrXozwe0/6opiEnpVqw7/7
mmM97h7r6n4BzglZL9YaU6Sr6WI302EOeZXKulyQKq4Bh1kFbtFcoRh3etaOe81L
ULWKOaTEWMRUGRFWaG9eZBZGoWt62a9UcMYNZBA8G8VBGBRzUxt9fdbnOniwe8qo
tqddzvbkEo4IYJvOR8FLCLNHSCzq2X9lMdDB2XIarrmnak3jz8jZp2COepzFa6Zh
e7Waq1U+cf9Qo551XduDF1+/6dh/nBfZIaLNfV+owvzshdz4dVf6muWr0V7qFyBI
5Sy1AEcsd43I6lkJjdUu2LhqYEIoAnbnlin77i7t26DU0kzyQCC05EdHYGrx53Vc
vcPc35RrZyM1wYKZKuStkidrQfSLxnWpbMe/0GES6teRi7R0YY8poKzprztBmcPo
Zu3+kGRWdwnvtwuTPJQycXSPNFbyw4BQrkJ9oP0rSbZtq6a81IJBAJQ4+165Euhb
YPSjKWVhUkd45cwGBLcTPdohNOHc/y4pPAg6QIXHGG0CHqWdILe+2QImfVoWFKPe
YKPlejgJH4NWU4/hsXv2I9i4Uh2uH/lLUDvjzatq0bNrbWqy6/7gN8m2INc0u76c
hOE29IARXzJwJJ9P2C/jxi081hB5Oq1lNCQQjf1PHEnbDllIcu/yHMKLksx0ba4t
7Pzv0vHOW8yFuNhHoKSb2HZxImjnliN35Zn8hF32s3LtJX4nGxzTX5EToDDSZRGL
u2GYz2KMsZlSX7pNn7lYOG9T5zOOndNRa6AxQBMRegi7XMMy+9kjx+jzCssELWm9
p3miCiApmfB9e7sc+bmvBcAO41RPReY8fE+XMM7XEvOmH7kO3fQgxeWQiXBtzhjx
eURmodLOxyFb/9EkeAJJ3pNNvYsyCfy6KM3MSUa67J1H8owPtKq6kVcH9FeddUTy
F/Z+uF1DXoYmmpAAmZ1fZy1RXUUmb+3xOIdLgAhws+QN2ulpXhn+7xW79Ta1yZdG
9mIajVGHZjJlBA9pzgqE4g==
`protect END_PROTECTED

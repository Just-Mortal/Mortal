`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wz6X3eBhjnEie6bGsZLRUgyEdAprdtVlZ33duxgRHZCWdm58KUG3cKFm4rn81Nr
GnrcJ5QnsXo58ZM6laH53rtircpitIypXayDGqXBhGAtwHGlK5DL3FN+uAmxz42I
X4L1AKc57Hyv1m9j5KXzxEGcEd/wo1vp08oonVn5iHWOHGLyc29tvN5nbN5tgycj
md4CvOGjJFxmO2dSSl7h/1orjcO1yuTMfLKgxKmfG9Gcw54QF0eio8C7YB42swOX
lXBCQJ90Ifs0a7oNNuGvu+/NSPIhv7CiTpeyM/a6Var1Qoggww5Y7JYK4XDsDABy
VCT1LAQgP6htSR7G+BPow3khVGFhRpbedbcOlxNqeA9XFEjKG8Ri0Fr1wzQkLYj8
UywWHuhUH4SbGuXCuQg+4op31xPMmXTV5MS/Od1peRP9GlleizGB8RXTPHoCmJ/f
qTi/XSamKnII3FXpiT4rqVzD5rLa8MdYp7csg+dfZlgZscjP4dfd5mYj4b871JpV
ry2GpTUda+WRVU0teHEa0GsX/9Vlk9GPMopkLj8Xbu6vkdtrtDHlULVMzkXSvnMy
d1FAeNr7MtxBe0P3Eo5AmA5k9bp/IGO9Jq8pqfvp76t3NtIcURLuw2M0KK94I34Z
c+Y36/fzWBtbv/4ybklNvKMlRWP7j5L5PcY6nBuZshKf/Jyy4TDx0yfM7oS7lDGr
AlVW0r5k7dLd+MfCk73GzaMY8A+ksYZKXEKLhtj8dJkSIg6ue5xwSzGMWEpFlETt
UHzf557UDOagBlcZDkdjlsc5R9xH1wB26UNAxHHH0Wlwd6yBGGfmw/lM1rUtjus6
nrQVCw7UQVemOsh7qSKkMmI3xTy6Wxy9eB8cnZxuUQsf9vEOpy8PN5nPZvCFQxHz
uTHoHFhlMZ2jTc5DPIAX2hlsWL8/RPMiT7DNsEGFjJhk5W8sOyjkTaTOpntyxvBD
6H4+iGtGzWzyi5XxQGKdXFV51UumZ3IufsSP/73bwJyCq+PsMLDDjs0AU3++NaTQ
B3Js6CZbyuWo5lg2J7o8h57MT6nNH4TTGLu7+jNMGHmKuw2P5Mh5560uWcH8iHhr
5RKDtXdzzKXuHAF621Pup1P/tvFK6gQ1LeO8Clk1enA=
`protect END_PROTECTED

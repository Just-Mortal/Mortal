`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZjj5hx+7UjOg0HyAcmd/UwKU1ob4Oufz4IWG6h5IhGfOjtdq8mGLMz8myEqnadD
ZHYqkIse7zMzBuKR1bPs8EEX5GmNUc56gNOaiyQ6QEHvsMZZYp29KwrHnpasBD5N
qFZbz0gVX5DCpE5PB0C1oos0/OFdYz12vdDuwKAu5NbwIjvZlR4DQbJqcWRFUYY3
Ee5KYztL5FmolgyY4REYr3KfFo0K2ygThw+t+OqTvLILCxTXrZ0sfjcYbmGN6sWn
/1dNeQauySuA9K6K9+MhvpMGubqCjtIzlWF5P3BEn0Kb1p709og5Ed1TZqBWRQVQ
GXFGt6GqvFF9dI8I8nCgFrVjyydf/+lHNVAODHNXNMBvkuQdW4lro4e0LT12Xtnb
YkSvOU2rZ0hsVAA7NnXnx5eZvMs7PI82J9XvlIOAa3wPLL3up7Bju8WSITWs60KC
K8lg+T3COsCrnYI/Wbowd7lc85NqxhuwQi909WNEjeU61NQ+mzfZSEPASXhVazaS
JwbMlJa+68cNdJ8v88EHDCxxbwb1fWJJc3jYg3v27d9XyqzT17eOadg+nUAdi51x
K5rWph1AXKNSe17aw0Lha5Z59oFghlwRfmAt/AISFx8BxWxMOsllTpzYEqUiRG+5
soD9aoUSGFBg/pAkesiGmpqr+Bp3PgvsoV5iMsRz16jgrGhQO6ye4eKhJJvelLvD
3ZgHf4Q3mvwkErhYxm4ZTsE7fVUgbuGpEbbFveW0CBmD1nwmL2VruJxKNFa3ANqq
7057tDtMAeVzlpkS5NNQsybXa9PnuDH5EvWUnBIdwgJi6kgkXHa3mhl59cRV9sI2
PkqVRSG9f3AIkI4t2h9I98p3++Vpe0jA1I0C8T9JOkOqEZPHZrfH+pEVD9VMWN+u
1iIam85vQ63HyBCqeOmSYS9JS8QY7Oetme0PTTDXjaVNGhW8jsNA8MeaH862nC+Q
hTFJaRPuCZw450Y1sYJiyySYYhpaHKXeKudcpAZgs+pVUIsJaL/Jc6fGZWPBlb7Q
fczdII8n2GBAh7blaGsMI3sdYz5r7b05xgojEeLzQx1boiNU2XsXuixRMhBwsW0G
O8p5WLskhI+7UFyxEJrmjPrIyjp4dAu//C9ozI5R6Ib8RrNA+lp4Q8QYx5Zoms6L
SfrLrqT82bcDrbhhIOLLzq3J8/Dh7IeOyz+OuQ+kmBeMzwYpeVSuQh4ncDV7DehD
NaHP0zzAY0JLEwQW5BP33iGHxyfdJdG9RH+KDf650yhbenom4O151I/oDMNKoySL
wn0nd1iKaCW/qbXPeGVdN/NNKpzqVBhR2jb+QatbxftkDB3BD1TOtP+6V7YsLelE
ehgSawe3uD2hYwI3Gn3V5qj/PJi4loXhfgHWRL3EuCCfToHTvnCxEIb3N810Scbr
RJsg13+i4QUvPdukw9v0sRL34tLw33hSIle7queN6TjVxH7KsD3I9utFgUVRYiSQ
bB1I6d0IScTZ8GA/4q8/e9O7t6ZW8+9Qn5yVZX5B4+5+5rFUHC1BJX4qR5WY+ZRH
+62bdJfs5NHoE8/MU+1kTuou7Vus1dg7dHVU7g3MUF6DMmhIT/98sQFSV/n85dly
KVf6bCk5PTSoI14mUh1Jovnq81CvooLpUyCRnpYzM5+fM7Vyab687oXjQAz81ZuW
aocVNuNUlqXUTYg6+Yk59B0RvuPraP19yXlTum27OX8jpLvzZY8TjQcmKJ+kRLCJ
URNib+vfvV+/Mqnd9saJ3mmxbWE1ZRIBYSE6duFakL49mkM9FSxAH+Tf6dBvxsQk
XDiRsIfNOJumRyOqnnMEoWbKEjTDNTaZrSiDFtlu6eWq40hICqKV28RoqT46p0Lk
wYaEO+PY9MZTQ8LUZUBSzhxcCWPTSmgugEtOnp0nsYa9orjJnAWSRiHaoDkr7oPJ
zG8F0wBATmFwetgB/SrDrRYelGzI87S472tbH8HfguUrIkEel1OdxyMuEvEqYvQL
p7Uyb/R1Npe8rGUIZTS42uH69TzY9EM/CyC5/Ds4UGaAlkFJExNjJhGK/7WcRf+l
UasSpUFqmavYFybvoIMmNOU5oqIPkus9Dn7r2xCkAdogpPw5EjdNeB+tlR/mk+bV
lPSOLgdyBchhTwU5m7JDUDrpPioprNiIrwC7vgzNW4/ogFnqqNso3ZMNX+wc9Juk
QApJImyXoAOL9YNH/3h6oFgY0FUGfP/885PC2o18KNzW0Rb/TlMVLu2f3G91OfbP
72G91V+2IZ+BUMhtB9t58drMlyg3pYY54qzRKG8moKZnfhhUBv48VKCFG/KidaIe
IDTZF4vpfvUehsD7c7XUIlZLNhmJo5Edis4Ofn5uuedZyurl5QSvb3o7KwlJtZbB
n8G2RTi4SUyTJ/zfRaN2JSGAt5y/qHZu639D3t7wMK6d1tjApUTnxdHiMpiF0zEr
/vJTU9Sg4XP7S7enuUi0PSzU2/8J6piYcrjJOcBDtWkoMTfKNTTjN2Rx4P3gbeiv
Uv7XBactbRBI1WN2Zp+ELpsse1Kq+oEA+Zc/1U5aMnGcFTCXCdT+bA/0sZ4uZque
7lrGUoc8NstqqgXFa/iktFP3jYmOSHAxJs9rMrt7TtHL/ZAZb/6qi2SgpFT/wRUA
6gq4At9MH4D4qILPRqM4uaWkX/TqkaFld4GaJHQvaCZ+AIBxs7tZ5oOGecJCkpZs
g7QiqTHPTDIMcC96C4mnEO5es4Sf67D10FQnr/zKpAOZqXXnq/wlJUsGQny5CcNN
GmThrq3X8/49HeB9gToJE0GIXrjKFmOwH5uvOJJtXDLxRutSd2IVh2q3Tuk3Hi2a
UeSXTgHtX19Nng49YPxuP8DFLiyfPOjsvFw/mXXgeE2/VFXoQ1Ia67lU6kl8z09x
dp03uWH85eMxioKmCsIvXAYY3UhtsPzHDijxEyPQHPTUu1d9fKvOrGfWs13k/kGp
X/So/Hxsei1tIeT8d/Fz6uxDOlU2WxW4Rm7ObEwo0VahE/ebFT9W4GMoMPP5lsKN
icyf9BtuxpusF9hL1ajQFBzfnJLtp6/b5685XKsUYnySePGWkflHz2JxxQBKf4Ur
02I9YzYNjS4pV8M6HIqdvR2cMQcFXZszQr8UW1rolqULNNEmRoLma/Y50vozbu6u
NI6sUYAaQtlZhREaKkyRN1ZHmJvGxImSbSzYvM8QvdnTvGyK79lPdY8nmQuvpihs
aiSG63Cw+YCtwfOdH5VsyWbahKGpX/F/DfaoMUl2IFARos9i7yNhdK20/rxijYME
lulsbrjJ8cxNJwEPi/DhXgrR05X6YpDOcJx+jjoyDR/zy71zFYbVUqA3wPJ2RFxo
KuFA26PMEMwC3Z8IgNoSx0UJPmRNlQAsUWCJhaFpdyQltBZZT7qGO/CigYUdwRoj
iQpwSnvX7NgrFuDdqSoDHq34U1gZONpBz1HSCQ4HUgfL7/aFoE6HgZw8d7V2epdk
hDeXzC0ecyZOv/HRb4Bsg9bPec6B62rorYR4iJrU0JjxtiAXuo8BevpEwxazw+dw
QEhLVL+RqgAlMQPkwqe1wdLPZTEHxC0ODdcAG/Ff6J5c4IwYwea7tiPRr3RWN9Fq
+6ecHrX8jwjY9IYcNd0e7i1ZNa8JTdnHXEKzldniMzNEmnOuxcCRsrQrB5g/iuVz
OWaUJSbJdj1HELfJ0zhnCJaZ7CLLGyHwD1tBeAw4kzUyxRg7XpdaIu+7MmOJIxBD
OOsI0z65OW3pu2B0X5JSWm1Hhaq//WTvT8HReVIwaiXL94US9vMlztbUQVbX/H2Q
H4NFS/YBnWf5nUwdl5sOIIGacckQNCj7MsPexr+xfgZlQL+02VSXuaNqOzG0p7Mz
NuKwbe7x6TNyrPTQkuYvYPEWvfTshuFU19A5jOY2gtb8PE37x8oYgiX8V8NvcIV7
GQM8wjTxHZz2mj0y/9sIzTGC+fQkHXC+e+y/I3aU+9lQgb/Gkg7bGha9T9H5hIs7
hP1WaHX8ke4azfEpV7T8LCfS5vMkmRMvpkdWkeIukv8s4bIhiI+gqH73XT70Jy/2
GQY4CcMPYlAe7XoZVRK6DbA/fXTNDsoZoBpmxVywsAmGq3qhE5VaTHck5sOegcxq
m9ArsCVVkiPFLw8AKBwIAlYbfUhKpF8UfS0Cpwl8bvLO3csVhLC0Y39Ma4CCIoZV
Y2ZLBm8sBUiRz4JrgMOrztUXj5SZ9IU/jfpOz81ykUBJiQttlxM9Ig60f3FEHNCB
RrL/IQyS23p3Ev5g0WNo2PhNZVkTy93+KAZ0VbuI/l6c/AGTpmcLOS+LU1/GnylF
FtddautnH2AUfvnycRp4wMTOEQmSaT92emiMQ7PaL+AKjWr64LzPplgJNHnI8SGM
QAJypbcFMgoFGhzj0VAyfIkQpA4VGujcj8SQCV9B/1z3w2Fg9I47GdoSUJwMM2rQ
KdqvwCkMK4OLM7DFWsb0eav3WpjRHivRN/ZkrUeMSzRDfd4ymWVA/EeIJg8EDMIb
DsnEuGuAoPY9ak2FvqHDlYu6sR5KddNePbLB1d9wKp8QbmMebNsri1+K03+XWWwB
mIQG6a1JusysIs9Q9dQ6VHlGJPkYztSDTTdmjWW3EZGaTb9yHnIWdHdNbNHXS5Wn
HQUrl8/t5bxEuRh9Vhh33wUGd7bql+RnRkjSl+K9KriR0BZcv95NqB0UKTTJGc6c
qRJTRPMLqPEeAzCjhZUCGUPb8U2MCnyJpbbqmhw4912lgS1zi3IHjcZfqN/QIjVK
obLdDEsR5DPMsdtIiQJkhU9B49/dHtmPqTWZ8oRfHZ9BTSGMLuA8hs/oKGqKL4kO
sI3KJEvvTV1e3gJZGXSk8CGtGD8Or61FpU/dbtKYLifdbJdFPg5UkBaFFdZTndE0
bledix4Gv8lZe/VGkPXruhQWENfI8V9qZghY3S8vrU7vGerWbvu0zJ79RAwZLO36
aDQqiMw7c4VW6AZNPhw2QAaKth12GuiTPQV7Lhqb8TMPXqsOvV22LdTV8jYOFika
kXGTTCaJmrO942GUxwTHcL/yEV+00tdnzAGsFsEafdgwH+1Y38qiK5Ts//JhcWLk
4mHyx7dVu9CSvOPqbdODNIZjiu3yy++vj8zPHIjNPsuYkOX0EdnsaITLaYd8tRr7
v7fm1h2+5Nq4df3S2sycoUib+ggVvrYMua8KnHvn0XnDgmZIixhLV7fL9Q7PonAm
QZHa8w6AbmruODt1kuVlEVM/7IkWMZy4uQLYhuUhdmDDlJE4Aa4H1+cjW98b5NMh
C2sHsPcj+/cyzqNaNZCZgH5YZI8FKZa1VsULf8f3PJhWXdG4pv0V1oUsZGFctjVL
+yayXIw8//MYDPTfN7ItajNJdr92kfZudFhRDHqm6r2Ok8tjyWS0muO4ByVVUYjr
6V3/ujsiOsX700jGskAiz0Ka9cCxmRqGQnrd0rlS4TStXWhhiZbGPGXpChqJTAQT
FkXYxA922J7Ho6sGOb4h6Dqavw7RalYIltLmtxA2NQmjFfLdUld9OdNbzzR4eLtS
YlbFHeri/HeGGhdqgccCftpd0r+9Y/kLiu9ci8km0QovVidcZC8TlXMo4mYUHVUs
lgv1MqaXOyKd1znrYFcufujjL5vmcnX0qwamzmQQNOc+YCuCXWTjN8LuoY4DDXOp
Y9McnjUOCdl3cR690W9iSeC7osI25LiPHcb6nOXXS7rMMJNbIcDz1YkjFHOzhonD
4MNWP/KmsXTP+B3AGCGNaWT6Az0oAYeQBxTeLcCiChgnhOe9mLuSYn+EwhQMxT4P
/orBoKdVhk4iRNXPKs4uWPgtG2wxTef5T+XWtUJe4csRn+ghNCicukSUYYWTVSJw
QzAvA33onuKQSw7hdx73Ktx8SqWCIgxbroVGIlhveJ1rDyu7/E1VC2Uo+45r9irU
6U59TnuJrapvt/j2CyGgQFxJ/hrSla5dIvAyuwmRGS9TAirUJ+Eu/4h3mM2ePkJN
PoeqGEiA53Jq3LqTkpaWRJxCZbGozrlHT5H3lq+W2B/UdocAgOlLlyPGNntXAfYq
I7008XEK1kcMwBm9gzgUz/3fttsX90T3Ogb3F5hiIhytRIkuVuuqqAHRCFd3rue1
Ftavpb7RTLumBycR4GHTWDplasKF1hCme4MME0cRiD4imsTumkJC3eN/gvyJzmZ2
GdrE8lztg+f/5PUp4+AZW88TfvvLCrNpB5TqC0GN95vi4vxEkuHjZUTw73i3p4kJ
fC0FioejTq0JMEg+UO21lChqbKKYpqa6OMlAj2hHYj5V/vrPPASSTF3XRF1KmKdu
/eUN9jD7483yMDDPxWUAxJv409hehvysJ8zRzFsLHoIxEQELTS/uUKW2ZR71Zu7l
5lExKFcHQZxhaLB/MGK37Z87t8A6g1DRZ9QxKQsG7Lzjl+wSJfISWBtWieowErH7
jQlOC8VoFg+LuC/kSnQ+7/QlbHYzJRzpRnmnHhGNRosP34QEiwG0Ovkdv7OCXVs1
V90FDBrpSYIYAaGtKzpZ9Lld1nxrhcA+I996iiRl+d+XEeTtcpR8bkPaEaj0qWci
qgJHLa691pSbHqXlAOFW7cfWplnwcIlMUgu3FbDk1sSWThDzjeo6BFkUrgfP/j01
5EtwSkmLdrAnJmxF9Re1KBGeXivxXFh1VOR77R2rPmZrCQhlst8GwZRj9rk7bSpE
3060Lndzwg0tt4Xn6Zh88llzM2nt6znEeZySi3w7JY77M89RthcX2WYm9+LX0i2Q
KJyT4wB9z/K+lFNkJSCkbgwbClYj1UeaMBLGk9ijHb3bCxSkuZFsm8P9s45+KjE8
l9UaVtl1YSM3skpZh+4Nh0UFHnHlNxMlDgtRt2AnHKAYdQdEZRnW3k/p5E9aevFV
WQ6dVE1V/l1wcOOfebamfwYM+DB+5U/DKQGiEuTvu8w7mX4t9KfzSOprFOedENcx
q93gkaCIH3rpXVGlDoPACI5NYnzl71u0a4Be66gqc7mxe13BpOKwgg7MlmU8w5If
Xbp24AAs7+kYf1TDJq0H9TlXb/zmjRg6rcxGeujC/qt1JJnoGKr4yBv1Wo+HC0rv
9agxSwWXDmfT73RsspU+CbOIqIqwAC4V4koFwMsEI+cdoHliXrhEJd1zwbbP3Hz2
AHbvjl3kABR+Lx7WQ/+DRx+GWVzzX1LY8w5xreut56LpafPXKar7P+NZ5ipDFLOP
OHDLb5DOQ1aD+DtgXdULwFY0fYuLeyqdhzMR9r7ZKJEtY4oUq/CyRj0Pg2T8+acM
kbnJZni+sRsh6wHJ3L7Cb3ro6L9QddN7Fujxe9x25oUW6pXkFqdw7P/TtfqXld/p
+iqMwyppDy03FZNUdjwog+I2JoOO+AgHoT8T45ebX4kLPfLSyq/0b4WAfLxvVPvI
DmR8oEaOTDaI80ElVcA62+NVXp91MxfVuHkZrJW61O/GE//U2OPiC94dvpeU3CS7
27Mg+lgSDD5kcA4CJU39XfEsFKRWgXqICk52JUcXN24Lua+K0BrgDUbZVHAA+CKy
/eHV/WVFnZWbci71lIjBQBl4tP3SrymYz4oHPv1XOq7jMssAIOjqIlqdi8Oijy6k
cZs+CwlbFX22UZk8J97sSM8+3nTrt27ja2pp3gaktBVQSFCw2OE093EHi1l2t2dP
yAU4IJbKvNbACwwI3Ssq6E5a22IEaGhOZ/+uv43FfqUZOr4OpR2nuDuVN7y6LTo/
2MuXBDlygkv9pZHYGe/TxEJjRE3yIirVCi0qPYXhyuoXCeV3cw64SaL5XVTgxF4Q
wU2dFJaAEomUt6edW48QHdwmEYvHq4SahzvfNcoIOuPZlxaGnMlAQfiOawCQXYJN
M5xjTxKQu0ppw3WwMg6CTcaONyHVF8f102JNA6Xxa7UZh/ZJKnKl6yMG0Nb/utBT
JpbaGEIKr9GGcyQint9JCcd/khPjdNhE/ZMMX/l+cJbCs4nYFcOfU7qLQ5i/Ygkm
zTvpqspj4N3QiG6ZYYf0vM4jUqScvBTw/sFfFOzk1v8IRXIaze2vUSdXDXb99aga
FPpz32AdivFdmqwdhIVmEiqpZG3beONN/IG8jsvtTA9K0s+J7T5zRX7Qb2bsTduq
3LSGhIxxDUA1X/3HKXC6qXN6P+J6wyrKT8+3jbawGvvpTaxPMlJIMw9H6Unc8rCP
UMx7duvxnFnBuVW9MNpXRTtasQ6CaJEJBztIl/qyo+0GjD9l2VRETCjBOUqBhjeI
WSy+499KkUdFHZchTFJVdt4fvCj5sHO+k4yPGl3Cc4OcDT+ieIIC3+2BPMRJFdWc
qDn2xVcvc1jYC8U4YJd7Zb6pPQ+pRH98s80Yomtct0IYf+lABkvk1ZTY+hFigik1
TUleatMNzmMC1lWI8g5PStcgDEQER9g9M63xnFOvjGIs8GpF40jOfsgw8c9z+ioD
GUK/5wCTPmfWUgJ76DD7xNb5tF+khU8uQV+fo6luYlcKURzioBJFpSeg9m44lPSD
0LSd2FRbi3rqtrBsZh059uLceoQ8PQ9Z2AEr9lG72hKWNH35uEwZJtUXGKWfvgL2
qsP2o1CmvXwR5Uy7zb4Kf9vJSxth4Jh4ZYY0IHhY94UX0EK33BgY9RNNl3w5bXYd
UVzmCavp3DqH0EAUv066jF5CwZrBz+fhcNsn0psGvEC/3Y8z3gDPbFIX95TzYDT/
yiQZQ/Y6ziolmvpNrR+0DP6l02NGoD/jxX3ouIdPepegN/NiEEVuCpTNEKtpIPHJ
BByMYoXWr2CcgjtSSX+5QxHpbXXB5QS1oKu/X9haPBMf9dC7aowVgzhbZuVCd6FN
pX/Hz8xHPL0aUg7A+mPKM+CZTJaBIs2nhR332eXinmvP5xL875wUHHoJQQYwx3bq
vv0jNAiVorkZS5HOszdoBdCg1DB1HqvITwz53ZGCxgE6gxKaew5S6/+oWwYoM/QY
X58TZ8ttlooNe8GK2DR/e3OEqm/SbOAvenxmmVhTDqmSMxJGj0wrqYCkD11S/agQ
gWDSVaKvlXxubqROtrJa4SutP5Zvw0ZSBnl2oXlekBiaZ6pl0qnIyXpJeZ39MLMh
OCXCqlbfvBzpPXw4MP2hlQEGGQsJcoO9ooDqbyvBJgpwfbajFIZ/sEJBXbQu4wQH
TxH5ANqn5PAjnrIogTHkb8qTDpxFr2dMlmbfvMwKcKgzCrDiipKHuVuffnJH+vJz
Ui+gIrfkKjWillTfvpTUy7djnjwRol3GmOfFyJOQBoxxCIv55UnlHv78ZEPHtR03
9ik4Joo+3uCFqzLVDXAk2yEkhyyA5RN162puqApx6b3+vcoYiGc2XpJsjVefGWYz
SSCeR6vtKUS3RfRq7m6y6SqXqyyvEUEI7u9A4xItq4M9EkaWIg3JnLmrgee6jH4A
O+TRNIx/dPY7D9Fd4E/j3xIThbOZ6qeeslFQ0ivDzs70DK0+Ulqv5V2Wrjr40qIn
3uWObcIEJNKeVgKOtXWbNcV/QdJ1TOWyPsSjfnvCYRH8qfgvE6lGAwASPhPS7lfN
`protect END_PROTECTED

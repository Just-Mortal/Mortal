`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/XksLTeZwdYIocy2CBd0Q+U2nSHfGY8GVmlJEYDp8bEEGNczVJ6CfnKYOx0ZxMG6
gdjbKEhAyL8Ac4V0eTZ5U30UjDyVA8dV6G65wmfYET1UOJhhw1n0Ef0FPagqSyZC
3NBem04kWBSZsCXBbytayYejx/B5qqW4fFvIYUDo7K11CVAWEUC6Mv/xPY4fkjUo
4KtUdijRkqNd4czLkpk9v0FSc9ivR6OGBGzV5fonv6lPG+5SjkfGpqIqGX7AhlHw
Qlc42lnHblycrTUrjXt95+P9qR5ysf+XA3izRtZiR2dZlHdAJD4fiNMvX7r/EQyQ
Jx1kULEjj/ejsB3qJtkKsaRqLqD7JBd7AqgZtAdr0sSiI/8jNkRRZF+szNkikkmb
sq57CnOVCrtMCj8hHVIRURxIvwmQUl+4237GQGd7KwqVT9riGT2ftt6gjPVBzjaK
zWPLgU0e7uTqbW3NPO8vDc7K7N0wg/LMAWFe5zCk9S/FrNIanhKuPUpOMPpYKvQz
ljwwqCI9HULzHtD3SeEQRtkKPwSG7w1eeg7nfNjNM1nVs/nDOqJLVe7TDAUZ3A9y
OxjLz0J7rkQ90rwDgeYTzn92qNOTg1+UaMUgJxoUt/eqSU9234i9tl+GIA6VO2x+
t3SFLVwZlY+v+L++eV282stfRp0h4artlgJi+IJjdiaHKHW5PyRfwHjSIBb9x4FR
rxka3PhbT2npf1Kc9sh4md7r3spZUxgh7DYwbGpJMRHhCck8CAb4gzXb1txTMWIz
UvjmpBpF+cr10Bf3Mfrlf+E6ogy0ZfnO+fkxfVTsUEvLB3HGkgrjquQ+u+2wPL19
dYdribhHfJou2qphAXjiKs4u85VGe/wpPwPOwRDZZaJ23x6ZEpwQx4/oNBfCqLRK
sL+RYjlM4aLJlJR306D3jtbHbCM26PVrY8btuS9Jdta+Wqfub+bFU7vnBj88qZvX
45C8dW4eqL3dR/QCTchYe/9KEpETGcMbYp2qR9vxSS8aw+VIjB9lBLqHsNcTQ9Vm
otkEfeNZjCV1rKSJfAFmEhPWLSnViRXgpFdG41fWmRenTcwY9yYYalqugO5R4j1N
vucGPgc7fw6uEOY2m835HqdgRbvMP7rI7elbWzv3/7+MPHBacEiOojRsGNH+L9tu
yfUc3FhTESX0R39A/NdTTH+Fnl+3rdR/1NNHyjX74C9GdMrzQHMdAqWkBh+wMG3w
D9Be2vB+NnIxDHr+U1sI8fMvZobmRSWM9AqMtSK1d2sOEj7Y9DyHMv5eySxK//3t
i5hwPTN7VOjizedwgF2UnJFVMOrMwi1ZMZ/vxYWwZwu7B4t4H7oauajrQ8bYdhxR
aYSfOhosMM6x3c1MBuzHQpscFfwuwL1XFGy10eIK0b1vu6IJjA/c3/ZmTDM03wwF
nd1IXoRPNK7V7qUn7x0bdccl+WAD1VbZh7BqVrXPCcPdaA7rKeg27rSuKwP7XZi6
2FBGNk4LccpvtE807fAVTT/a8UtVb71xiAIpOkU6WhATnC3aGOcgIDX1haapfEx4
6PeSGqXX6OaD0EzmMxAza9HlvBORFh8ojaWjjonhMDs5YCxauE7a10KjjL1ExUMS
6Jzxn/C5rIX397k7O6HWB2p3LamjJv3EBMklqoAxdtOEIgXYxo1zLY62zlwIKaOY
N3VTSmVSt6kyjHMc1ew5EInDnrHleLrQzHbCMTPu9H2vuyUREwIO8wnCuMTJQR9Z
CgKDeHo/LLr8FpNaI4Xs4FxmIGnNS9ehbnwnfBp75Gw+tYwKWaTpJtFcYkUz664t
7RK6SPuvvFIvlc/A2/MQYYVgGOv0k4yO6d95rnoPsOeacv5QTwKE5fehKRJircq0
rowb2sxlUWwd43Edwbq+Jx019Y67jb9c9xiYhTWEDysnvOj5WQe3KPVaxqDB9m8L
7SLlEGjQDmz/BFAiMZjf15uZz0SFpI9G/6I1uNjZ7vCKysmbTjdm6b4B8YgzVgQe
bvrAGlwU3k2Bg0WLqaotVlUr7nSevFovZf8L1O0UgLdgzbZxD9JTyyxvT4FWsyvU
zI06IkFH9dI5QUU9LEc2hsminf499CS4MNZTigNgjtzvYDe/KkNjwmn52fqQtzMB
ozDSwhIWWv0JxAFu447vUM37M5cCqP0Vc8tC6PDoWuA+CJF7XUan9EpX4KxGNwGP
90d1NQcgqZz2/4r1UJIRFBeG1FWRIi4DuXO99TB/8wWPximcR8+bvsEdXKAGPoHG
wYkZeZTPReZEh7EQfSKf/nXxAFUKG/L8djYAd550i3yVWm+Bs4IYNoC4k7CQFSlt
mKZQO1vNVJZVgaLdYPJyTsdjE9pk0XMZ3r7A+w8+04LOpaLldS5+R9m6GVCKaXcE
1A91Ta5tLNiahvj3y5MttTqK0EC7wUL/Y4vzMVpldfmbyB+iqz/qGiR7rkATbKiN
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kpr8YjbrjmW9uqZPzAL24HYitU+JVTQhku/C+KhtSaIjZ9tOGwPNxrkj/YbBJIKl
Vc8+Mqw0Es+2z4NSNSUWGexNMI084HbNPWWNHOnJBM9O8iNG8tirTxpTvP+QHOAV
nl5PPvu4DTuL4hmFM6iQ4BcpImXZ1yTCqJHER0zZWISNjBIQuwBbgKr6moAu57cQ
ol5vQXpJmNevri7ia55SfGkHfnggq4U9wrLZjHzh3scIVCeZ4B5q6t+zFJSCgEvD
bhwcZKLmDFoQRhhsIUMPKgYky5q08tBOjZ4SVMvMvfbUJvrG98WskAahg4gLsdEt
1/Z8Im+AD9OLOZqzRLEmk+mdRTJrXjeKTpZx/LOs33RIDBxce4Wgy7fKfMU3lLnB
QNWADh7Jdh18GAWvugYhQlOVvatan1tF5kzhRuhFsO1afZQAhaW3K8dpp9/1NOIZ
SoXdGz6opn5zCfyoZpmbEfSddXrIIgyx7EWLuKSu4S0nUh5YSYbq5RS8aHVhCsgn
mi7DIsrutHOpCaAbKzklWshOa2rBWpJNOZS/iTBnfm6tqqgN/TKzb3U7GMY6yz8i
fpBxOswzyjJrmK9QDMNyVw3kfahI6ktzFdSpcxnbdfnuO3Obv+tAuLO7odLssaUp
8YTnYj1AXxW6E84dBZ7UiPpUzvw45OmfuPB2Q8Kfta+TGf8fbEfFtl7BPstlajj+
dJVFmfFvP+kenEtrBk+YGopaV99FhYhWNTb276qpOVgjk4CaA1krB2rxq309MA0m
BmrIH4XgOMjqLeCryfGgBF1ghSdisS8sio8uEYEdvitoJdbc1xZmECe2lJoGv7jD
q5IfXCghhY8BkEvLioJ+sKsP/cCAXpOnBefQWptlLKfGIocD9Z7QylG3w8GzBfsh
fzWoqyKeThlhuxi4sXwdNbhlizz/HZDsik30VN0fQj7V/hHpYkWp0+fK1G5vFA9x
2FyPK2Qbbn0u8LM5o8UGBlV45QhwDxznSxol+6gNKd2ZrdhiFqwtiFx0uy6WGL9d
28njR47+CT0d9+tMYYEL9w==
`protect END_PROTECTED

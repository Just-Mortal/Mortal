`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6EIogq08rPgmNbXO4rK3Dylt+IZlv1YAnuJoTbQP9htyOUUG+YJPGUqosUqLvUak
ddSKVhew1a+XFt8Wwk8l4johDgX+/ITY13x7+ZcUi5MIOLWYvVjk7/X0hnA8yLC1
GQTqV4pjbNxFTTxle7zrIOEnmRjHwJD/DMcZbb8diVtG+cbyWcLUSDEHsBfKN8sw
xS8cPMEUNg1bzWvuOMo8tuRLihLsDHvMJSyB7CsjjDSrIZKjHD/GrpIDlo/B1l1C
cY1VbnCc/XbPbYXeSymIOCdFYUrY1lgYShM+GnIeQTea0lhnsclxldh8kuRN1Ytm
ssPAqT4qfNFh6rijEPHiwgGimQh9b+SFk6hege1WzebE0O78Rn7AajS+4ELyvgtM
xjEayYWmW5Ew5vBaDpPofkk4XSl7E70wbpkHN4zO1k8loDoHmp737ZULEHbRJ/Al
mUtGIPIObBNGHqSA1l27/Y+KGd9P+N5rUUspo8gSmWnszhcBxSRJ8dSbSOl9tHu/
JPRjfPupYp4ZXHCBdvI7I5tkYiz1z3B/wFth3/N+g1LkzRSKRdPj/1n0nd9Ctz0g
02Nrr/1f/YJaeLfDCYbZC1nrgHIkDRsY/mOpZVGFRnyDAecGNJLxXYtju/wmwWJ9
lg2xlMW3x6NM341jhXugS126+D6UqBU2PxWFolKBTumZx5D4ciYrhT2TzhO2eRyi
UNEy4JA52JT9ADmnSIWm0HVRPYIKO24Xf/wlIBaMrhHdiSgK8DGyzC7y0MeCyI92
gGKTNuBpdBIkJEKLuh+ETg8cIPcONoTsmLV/+dGMzHOf2FM158ZDn+6Q04u7RTOp
E7g41bToRh0UzZCGI7E8s2XdnTBxZBFDJuez1fchFgqoPNo+fogZ/zlS3hDzW2vo
QpXAd+rAN6hFgDllXv+aQmziEchYpvY15fJ0MYhcmV2b/p5qF2q5rSL28j9kEfyg
OP278xLScg+DJsZUaLu91eipXh7osR0YBCW4LAgQiV042GtaNA9aCZ3hwL0mQgep
vnkh0VtvBM5Ydo3rFRyPabtkK0ERqD6vWT7ejWtybjgTPFNqTPEsHa+/APgK2wHn
tUNJckKfbGOTWdxupCLYyELXsaY/dCyA3u3XPHc/ORAeNVlX0vYuyreG3iZxaqzV
1OK8VXVqb6w7jVSvvpfpo1ATxGxSNEs3Jr+BbLa+0fgxg5SlEtJNrXKcQeP7Tg7A
l0FDW/3HV8w9oL/4caSJb7IWoIpH0b1tBeq2Dj/8HOCYHIdZDsY0IYpq8RmsoW0M
GCrOoC9mTgBI2OcSbvAdeVCq8sD1pKBrZlq1WeCCgBpTXB8SloZ/3eGSZ5CN2P88
v1bOLleFuXrEfFGb3+YyWbsXa9+AJmNERRNFroJfCgWv2+KXbu8a3P53PStuw87G
I/kilD3olZYUP4ggo4pnLPCqJsmGBSCQcE3+mJ5XhRtDWCluppXnwcoXb4P/+SeX
/3N5FHU3QvGrMS3C4LOdfghBbfndeC9g9JpdOFYEwCSWi5aisezWevLcZKxUP921
8J+7DWiFi1tl+6oc5k7WvmtL9O7YjkLYTEF4G45zQYYs03LgoB2xYeXUUp12XgRw
UwHOE5r2y3iB0l0n0b1GlR7luTUdOFNYeYV1qaHjGpdUrfg3cWYn/PULkA323QJC
GB0cmXSF2qa9wLF2ZXC1sAYGer4wNiylNkPSboY7cUhA1GICMD5A1SoEHIN1fSCM
4RK0oiYCfw2GYnyGGy+q6rJncAW7GpOKiOosI69SZyTplQWjgKBVIW2KghH/rHzi
H5PgSxgjXbRnvCxTX8HQihA1qMXF5PD/dDAQXJkKzdpZB3CFiYSIxsDAauNV85r6
mcwarxURjn1wbfujTO2bi+cV0S3OorKTDcENwvoyyL2FLxDsN7jjOxtBaRkvWn3c
yvmGf2TnlnoUdFjycqVCtbhHtpBDcrlD/5yEIwFmS1t9BsK1S6IfYHNnqwouYIaL
u+pJRd3q2CYoZ0babueZUpOSfnhm6IqMYprAYNcGH2Bvcl5WGV9vJITD4GVWXWVi
8gicB17TnWe1Le9pK712vCpLa79PaooJ3QFbAhOn+ZPZkoA+Bgw+JLrqToz/J9jY
iT9axEhscefELf6eIok+svxiuLjtfogz+QhEuEVfY7XJ0yEOiN618t6Yt8NGYd/D
pNAkfSlHUZpsVzCYTqsUhm+bWNxcFi1cmkJvZPvyd1YK9e1ssZRyByTDxOpmsxrP
ZJnUhwvSyuumM9M5DC/V2tHn6vSn17pmuTdK2ChvfqgN2+iwBzsNnXfQNrfJiOEo
Mydm7yfbGWe4UvV3qGGkzntSYbXwloDJFndKAaCz5YsAJAPiORbyxU9VKHfq+N7h
Rrv2iNFoI04goQ9ifjXUvZL2OXEl7L0BByP6Sz8eKZen+ApPl2eSAV93ZS92MQEQ
QpIOCmAlahgFMLElc12tSm1v4zRaXj51Oxw+1R19pA+qJbqx5s3Wj4/HWObIcruT
BJfzb+6yIgx9q8u/yBiSv4fNz92gpd2F9mrG/WNHT+KcupHvp2alevd8W9Aq80Ti
nedQ0FoDFVcVQfHWHp5IgQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I1tfriVzNSjeCw9wrHl07EKWGkZfKyadB4tfwIXNvnZztzadXHS7oO0V+FZjtQ80
7zXxw6si56XVdue2A4o5p17xPmSh4VgF6cpgmiS3nD1Qic+YtELSL8KS836DelC7
DUasut5cOES/0ifhjnM0IHpyvTP9NGmFZzvJghikhFvQf7LPzyMc323Dgtj+77ih
vmlVKZXLbpk4y7i0dnBnpg0dO9oE6JE1I83aAiIBfMVfi20yh1et7BRxrd3/zAOZ
NtVQKqk+YbSSNwzWHr+Dbf96pImW0ZC4E22d4uRDDOTFg7WBE8tUtGUcrPRXc3hV
j5NJtLqKvdg8b1QbFG2aPDahgUhDzXd/CyD5ZQViwEFzS0JmqbiHEZ+URLMP9/0y
1+tPBy5sa/1v3VZ0vRhah8D3NXIrWV4Qk1JJEgZaUnyk9TM7cq1JL/0focol7JcW
SBFYo3zQ/EjMlgca2iCDEFtHjdSK2nUXAOvA88c0+dz2gepDV6F3c9NImCYMhkTE
bXmRtJP+uigcye6x+rpF8yNgTI0P8fChm0LrrhtpNWIAAoIHvZdjyOhleqwJl+4v
fJB8ThjdQZ/U+sbeY1sn01xQ9kNcPWzUV03L+4tW92X5Rz6ViuM1QpayEcJWGEjY
djJIMg7SXarI23CGy25igK8CdXenkQrZImJxkBVj/6Zxwctbd/yITqJd8M0HOnfO
fClz2cypS6Ye34XGBEPd2fTZDNt/ghzecc52VBMUOpbGh90Wjw6eXZyg6BxxdW+I
C92Q/NVgtWIcB9g7AQKSfQBUYfns5tB8sWTxLehDzXqb441CfOAIRuoai2MEskAU
yA7U1gLBWMc9AiC+RhCNUbcyM7fYMJ0zcxcLcQZx+uaucg4FRYyz0/rz0+HGg1z6
KLWROvRMzDoc3ZECyLJSgbxf3GnhYBVjfHSgNYYrgLep4ZQWQFFTq4Yt+KUmaNPy
q3fMk0QJ+f5mH7JC/Fgs0NDV/q6Fy8I7agCgNeKnkJR7WpL6gHWwwbCqeQIxENyx
+bpIsmP1q167mtvxKf/dOLzScycAyKf2NH+vxOYnVzjaJTcS/efBywQJfBuDZBbA
P2ExMvnnt/2wXXNHjzqe636P7SWWl9iwbzEjUiTIP8I7xRTCg/bJbIvMfF6ulvOh
ooggNYthFy8Ga+nfiBulVuRpoN916rjXMJKgCuEe/4hxWk6NQBRm5fkIVRZ06twh
2pFXv9ocXhngYe3NsyUi5E6ddxotwHfsA7QzMEYROGhen4eckgC6FSAIl7IU8jD8
+me/Id6DflabZD05DJSyCUUAtxGyyPoboi3+25LASsCJ4ftZug0wBTe6ZH/t7u8s
9ol8lDFNp4eyc2p1CRgBKSij/4nBG26IoKaym+qNvr7A1+5kmYzAzqkonfK5pmqL
N6voNPtc1QbiAaqAu7SMsAtZVRqMuzvfVO97uI7RcaPX+y3viVAkmCfZ+YYeXXpo
l4J7ZQ6Vfku7OJr2UOL5wJReuYuDKVsu/NXi4B4EKuZx/5KBj3/bpR45sf5naIsF
gq5V2Bs7kKkCzFyaHv3CuBaJusXHdL/iULrvVwY591H0WefFDTlC5vgxHvYcyDJc
zfMOch6XJhQGOAiCbb7zKhND8/cZSKhPtH4XiwMeZXPtMj+Ik72QM/Clx8eDByi8
4M4DYV0qODqZFCshDb7dSDNqGsx2AhEzj1dKwQ+L5Wek0ynTBWoH6FKJI2oFDVPt
UU8123U5FhsTm0ABVr4AvTvSk8wRwvkb7tm53ee3f8Ykb2qHhqRdXEwKen1dMiCS
Rl0cCMfY7ta6lZKepSPFfrbNDiknojfPF9EJWNJs2j9EeM36f9ot+9q4RS0Po4Sj
QP6R0ICDuwhKtApV7An26Y9XZ1+aIDce1Fd7Ef0M8XM9GYbI5a4baQSVq7jVL2KR
RJOteRDxYO4DYMpWuXmxr5T995PiayN0JPJXwlLC1+WSD4alR2NHJW0Gl2VmYf/s
JYf2zwnKy0XgEXuY+3owIvYSbkh0dIbYyfFv34HtoxVp3jLXUU7NSA/ONlDeqBp+
fPTJAkVCYmRWB0DIwKs9wo0gudDmSfMIilKMf1ZMHo4jMlGUKDV2NxOIpRETNKtH
+M/OYKu4q97dNh92D3N9vJ75njO6IuCJNg08CNLBOWD3bfoxFMbRxCYZd5OUS3+P
hY0FB0IllDIVuWpUkMoeDTaT7WHzP8uhx0U7BZ65JupaDl25/IS1/m5PlekUdMWo
6CjKqV6k/7YjcvrnXKL9nG+5UfsfSa1D+rWF/EnF0FwWCa0hBiCDAD9qzVpclGuV
N3EcU4XxES5MLqRvJcjUr6d+hOXkK0CzeFGY69Kpw3LwApvTSAkAcndakY5qtBM8
Eh2JS+h3x51QBM6wzy6DnJIH/YwlNp877c5A1p+oz0lpCTae9/C6l4GR7tkNOxv9
r/zb3+GmVmAxbYAyoOzoYcTomaFAfGOgU8/OiyFOIpp5OU9bGLKB3VQbadGqo+Sf
M6AFUqDIx62CDTjV23h/+v9vzvzKfMv+21RGn2Q80ejY7NU6TYLaVePqamhKru0O
mT7Wagq6bhIa92gHWhpd7SPptj/eeEoxY+sKBCCbDVEVTKroeFm0gIpwX4wnjtoe
taFXhWFH2g1/mq86MhPzGr8OR6QTZ3wthjRl8Ke0HoYS9iCFsSwDl0btmhV7lIVd
FcdeSgg1VwFOSN6iVKvSWTIGEe844HAhzehBzUDNnm41YOyu8Jh59ztzkXKFBC0W
XpRyZR+i2Ww1bo/xRtDy+UHm8Uyaul7v3lvCGQJ2MU+QdfUqXJZoRX2rMqixJbX+
oiYby5jydon37Y8KFv7OAgGuBrzUB0ayyi/khuBMS1s3VxLLQDdnqderFhF/E7J4
tapjwlkhoqLD9ULEcCGI5pWOQVN3NNTpxqn6JaS6EYasG0FLWZOP8D0BQUuJYiKO
Fiv9nM3ew+eOeYBX+y2RTZ4WOXW2GezZIBM6hbpgO7c9i5D6BlylNsYBsT6sp50b
heQOL9Jun7CFBKptctGGab36pXQwWgtl7V8Jz8Qo4osjv5+x7lTPY2Bn/DL65I0x
TSJ+sQUpZILVs821H3+nE48RrqFFg9q/OMNXeTEbq+4WWvtPD4a2CfyROlRGl0Z7
cAPCocAl80VnV7nEApNPO942kDX+itDJcBF6wpQhQtHVZyDCfAjLsubbvQ7j6Ldh
78BRrOJ1cIEPEMljPsJ2hGuIeCods7Po7l3IMIIu/6kfPemHpEfrKB1+aPs5GKYw
dCTVJDDC7sDyEB/u+8Qbl+MXf3dA4X0CK0MH1SDQ05U9CzsRtLwIdJ9qBBXPWWys
amTtv2iTRF3vMkJknR3NUgWKes1XhL8H61KLuOH3+1fOfcfZ2DSIqErU3xAG5QKw
CbDIGohdl/dGJZuoiAdmYtEAGsc29IDkpIJEhT3bE3xB+84teaoc20vMoOg0iz2i
WkNatmwk1MyIXbtRrioniEbirLDcz7byzccAeAEAiA3Rc298PD2HsR0EmkZxyCU1
wTfQDw1LoxQID+7ljSA8N0PAceqkbZ/113RX2ISJ6rcdDhJpsOeQdTWG2RvaC4CQ
uLv9+3g5TKFcHS2I7HOj0tCjYT6vyHIAZ3+eFVDHImts/92ciSQ3OYnl4VQtou1a
kDlkTvt/4Xgz4ia5zO3bzf8KsX7F/xSzN+en4uB+AV/5x+dSeBTNQAyRFWUXT9pU
iP8ZW3Lc76sI+XUtt+PDCM+1DfA0DMpf5WDOO00Tfj6enoTWvsocIQg6XvtzKaPY
c6/yrqBjrWrWXp1lZcImBjpp5nlBvbXvUPDDyGnax2MIguflL63EjQdGjbTIWi75
Wk6HZUUn6pL18HVlvV9uJ3lV7bZM68fcVc0EbeHOL2QBU0VaKd7VY/9YMjxFr2pz
YMIjH1JjU7/H8qgBE1ie61ldmRLo4M/ftzcTa9DQy25vNLLVZm3qzgeF2yGJBAV6
8EwqV7IVl4UVe627lzvHPWy6ztWkB8J2N4MVe6KYkY91KEUt72FFVP/9FbXzYP4z
XnrhXlG/w+YVgxzLQXrDiDA1wTuBDSy9HT0nEL0wAr4kMhqNcx+FGqHixbHWASIb
VpbQiapvAWpky6JXtfDuIR77WS3Bgu9HZAcSAKnFgGjw9thrbkHcLsBmbRfJFDvT
oGaYT8dy7Xbuesg6yYQdxEtVU8towaSyNHZtZ4pRDZZevMujbjPXaf+AXmtOox34
nfpEjhl16+NC5M02gCNKMgPYwhqnsuO0h6l8N6dQ0Ccr8ulVZF80mmx46OLpEaaQ
odyv3238OhJ0MaKHC0zwifX5C+RRNlegB1jqO/XgThmpPBWVLIBhTYgcYjS+JAUc
5th+9XFQSy2hiX5AHy1Oo5hlfWu/OcUnnrNbJmgNOMPnFA48Yxh+Qt3qQ05meaiU
65VQ6kbgzYz7YVtjgQ06pQudPromHTgU0vI1Fd5Rc6msnODohnnxPjS1uyf9mqgx
gYVnb8e9KlRUtvwhTuinGtArpIldgg8qe+noS45Ju6MaYoqwyThnQ3f8aCuzly4E
pmEahW20NbcKb2xlawwVms5+D64QWIpUa4mZhAAAM+om5lWLBaus71JcQSrEnfb2
F42Hq/jQkFTQjKFeJbc80ctLu6yxnBy/OrBnrGQ+r9MIwr7PzoL9OUkRhxZtennZ
dYfHQU0tm5nmnBifxpPABosMR/kK/MGCvKH/oIUYQLK3I+Ge3TqJZJlL9df1dpYS
gr2paSAnyQTYzIW2kQWWILGDMP6R7hY9IoLEJgUsTgjbZYwhCQmij2oB/eSf9j9K
ya5rFfGe4R5NNfc3RjFXoohyjrCqEqZOORA27Fg3gnkVT7TX0sBJvvYHeWN4E/lX
YxA98xX3JM2Fsp7MfgYgq2bF6ZVEK+V2uhmTCqWomcA8zW9V1Km5ySU6c9OFQJPB
yiLq9j2//bMKflaElmc6ysvfyeoGAAhBubaxoINetb4j1QlI6BM4Z85iDJH7Q+CT
XCbd/z4I0dFORZ2X6OGUh2a69hPMcgTecY/69SdAahsh7bvNfwIxpunvcXl5wN4S
QJ5a6Iscpoi7Et5SYznPSA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tmdIAJh792fHh6pen/TpyB07owlC565+0IfZ1BnYAngv0LfHCUI6cth43Xs4Bi15
dwKgjGF8wTYPpBqyL+M39qSwFKAqCfKg5fOR0RVqRRuu+MTJzx7YRDVnXw+gFYfR
r/KfsWDxTpV3biARnu13YRa0nIcpY6nzAq+CZIomvInXzUybTBX5CFVWpqlXvXhB
U8cOOv0559O72cU95Go/WjgtpwpGXOYj0o3kJTTLEjuqeJEv+c+u+kZIu+JkT8Jo
rSYbazC+3FaqCJlf2VMhypwHr0GcCat216itjgJH6UzRazc7qKoBmApte0c9SqBL
7bevKiB+neHEpLacWeD9/PY3ouKvaPZJj/308B8kaKNVH+05tMBi51yomoKIe9L+
iu0n6xy4Ti9vuOmYYBBnEWIC/it3qslFvG0OvucaGaIXhELQ6ABVo6LQTKvI97Em
rzitFTdNBHQ8/CLNYhk5khGr4UpGJAfq+ebMaCBLow2yClnu03BvLSFHLUuNrBe0
i3WpFxL77VxJtsvNwatUU2D5XRGGA7G7BYo7+c3yYEMRVs5PY6sZE0rqdDnofrjX
/BaU7zGs8zVlmHE+99qB79CAv9h3QuR154PKssO+ujU1YHEVj6O8xT4gQ3aH/UPh
not7w4ahOQ6J2uiY/42UTA/Cdn62LwvVd+T8IihyJ/rt2f/Cymg3Vwhs9VBwnS7X
sJGx4xNmkXtN1hm6Y/t2hiGCkP5QDyL6oI8dWhgvZhrtsH8quFfUgY/oBp/mnosQ
h+k9JYzWX8TfQTvpAotp6sBY/tUI7dieb+qPGRZNtIAckSLhSIk3GQ6HYuPFTQgz
qZ0z9qrAWWwNLjvn5KshHA==
`protect END_PROTECTED

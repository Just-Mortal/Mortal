`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asrNDXVTmaxtHoMGsEOcuAD0yDvYTuJvKP5KOdmkJabX7sTy27YbRvfi63y9tmTg
o1JaPuJAhDAnSgUJLNYK864nf1JAU8j/DfE1nvoYnWs5uK8OK2A8or/iCinF2ayy
VWFSiZ/WQUix2gfvcgJFTi3H7m9v1ROwhLtj/+H76dOQR5tyr/wI2M2UAxV3KeDw
Jc4b5ZklcbZlQmHdXmNrDmKUd4ZyzarhjkceDCvGIn+TCFQd3zIzeiJkiwuoMWVt
iN3m6j9IxiOefwwkvpmsLz5LSwTtdWSy2uGPU40fP/lx9ykwsFscOfZDXtCfDleQ
p+LImJVVjuYoinkkjdV4ItELRHsNnhnb7ad/+O1e4E4oUk5reiMWWDgfuQGoH0ob
NF1hM88X9pZSFVW+PMjEFzV84w9GmlvHqNkljcmNfuU6ArM5K6uQZxnaat0vHY4O
gTnE2F7BXyt5Kp190T48l824IZmJ3as0323GGdBaRXvm+4ypP4sFM2mATAspRaVO
3DAW7ICJdIjkDPbZH/K49uE6HKe0tcDhkyi2FWHFKsk=
`protect END_PROTECTED

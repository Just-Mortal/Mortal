`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/Px/LxtJNMdTM7306IBx3qayhh1vhAQfdFoGLvWQU1+QtkNeCVx5sYZU3tTtPzB
Jk51PWoKd0f1mwKw/9VnpIIWtaHTfz/p10SsrvwZSaQsOPyPlW/zRxT8dCGhkypf
0C1jLmvbn8Nc+gYWrNqBgVNUZdw1BZA2ja94Psb583MwAbmy5qaea/OY3MFAOGkq
FlXi4CqIMgXFgQ31NuVWVvLDr72YwFCPpmIZrDaVNZHNobxWceF4gyBJeInO2uNM
tt8f/iAS6o1dw28QVm9kM0tdhyjLGo4DcagZ5TPZ1iX32rxmPMhTJl/+/qqbiBEB
xleXQCr+fkYk+ZaE+lM/yeX8CTP+lXUIMYQmReqA/7PbIXHO/KVyIGyEakkpyY8K
8zW5sgyJKYK5m1RBwVSlvC5oCU0hzKJqJKfYMhGlLb8OR641GeNetO1sc3HxQdhC
gE35EFxObMt30zJFEvDmrI8y9pwo/+k5q5PrCp6i97ai84yguMUQ1whO/GSgqYXJ
AV3sfoCQr2Qw9rHgSIITZZS0jgo3SvLTY0nukskee6GIg8r894+r4X/tF3adIz0X
BmdawHYnPPl70PR63aGkLGf9BgLtJNzO4h8JThMws6JGTILu+mC8n6bG1QbxpctW
eV5idl9YDl7SQIS3E4YJkVS+YKIs9LiNsrx/Rce2ZWl2M0+nWfBnEdTa8aML2vyB
4BYUsa89gbRzMuCpMDHkRrm/rwd/ZSwBaeszHehAzB/hbM2CjRX+HiXKIsmWALim
cMgrvGPoJgJFHazPYkGfE8DIdn4JaiqdyTRkRxbbq1B3+SAVV/OohwUVvSSGhXOS
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rPGcah85PCU8UsOUSjFBMohXrjsWNtDV/4J7l//vaL5Kx6X73QooCWi1zJr9ExR5
/Ag+1RYCuufkp8f3dzBwprIPHrjkZepopOjxXWGAV42W1hXyksjevbaya2J+0lgj
IlalWlT1i4wuWhmnZoQvW4gfTV7TW3gYaQ9g8b8DHHV0O8NLZ8UuVerlkvale3nQ
svCmzy0H/1uFwq3Y2/2plmIGFsHo2mJjKQrK7gh63iQvvCZnRS4HYqgROHsqOq75
HeWT93iN/xS1Slx/anUfuhSwWCdJWockuM924ZlqXu85zcl+8NDnjZV6neDVvOWQ
9RH1tH+51brzVfdKVgiyFZmVNqCkY2o9v6QO6D9bkZxP0IyCDwSDoU3/J50hnHCh
qywYY8S2QxnKJ5DPZkuHBHI0ZqvI6I2E2X98+xJ5VtCPrCZMQrJ4BQFRSADjakgd
r3GqSeuTx3dvhBuZxaLnVjEc374fgBqVaRKzzMRGsf4VGZQ/ApDJLyjuY7a1HNDr
gQk4q2zZWfEgYS3OxXbpfpssFDDgNKbwksces7CEQatBcwRoAokFeck8WkxBgJYO
ol/mzR6hsywNySMt3GWBZH/hnA6suwLQuN9PztM0lT+KTAPuguWxBY95LsEdnuM9
XSgr54Difme53Uz6zwh2YKwBoTbsi9OzyAm3XaDyJq4QGHF0AXh/h2RkPL7BPQp5
Aqi89vVD6IwshefcewqzsPfdNxnAd3ZB5ppzHLDiiq7DswNdpdNuPl4pJtVU4U7t
o6FWKpIsPSzj9ekpKSChHiem5NB7L0t0qj1DoT9IZMXI3AZ4ckFsAf3XzrEOTjCH
OXQ+6ImekIsyJto3bjkgq9j0CA7Ko932iFOBIuvJHFIs7o+0Pd5tfOy/KXMbS8qS
EwoJY/JDlnIymVeXMIqwnyK9wDQrMzgEKfYESAlAd3xk4uwU7O+Uhctyu9J32VuV
HXg1MH6+1Ep7P7JHeUCKZ5dXpB3Ci7qYBfDhEZFj7VqMd7VN16oAQgg4AMtykbVQ
AxinUgqKr/E8M3ziC6hBoM4OEr4y06moEG0qsM9mU5lbJcNBYBo4GtiitewZU69J
vPxcXC7dXi/1nUCsu3ImSGsGiR6E7rslv9Y8z9+Si1FEFXNpM28lpPhoZOtUaHZT
2cCzoESPO9NbsFKD/NW5DnWbvkcUpbk2CmRUhtFuwpU1XGFELIkpyspc1KNJue4j
n50s7XkFDe3N97N0+NsifyKZbyM8TeIgPKrf+mR/pQh5WnDa/BJIal0ka9nmuPhW
ZxxCD3+hfaOMPf5xkvHp7ncwc+ig6a84LlT9molDmvMMeohpJzcefZBi6EO95KUq
lkQ/Msuj3jXhGKLTlcqBfUJqvyNAKD+No2m44Idfzffb/J97jzjwHHvcWWRTjzmC
uhE3rjsqqXJOOG6MwdIRfFhd2YSRwSaKPha0iBW1/D6qeo9jdvSIOKUeAjVjZEFf
xSSFIFqpQ1OxjOFLsHscuksPTGpo2jFrZBCmETVH5tpVHPLwYugsjQwUhYF6fR7h
2rcbdGHOYJDJ4jgV1KJEnZADmSGnBHu5OjDEH0i/ZQQUe5KtXD1+qYQHXFndVYeo
x7i1iXKoSKwS8/jhzP8B/6DSM5MPs2j3ynyAY7a/getr9/5JDM+0MPR+5q2VPmle
niupsdE85gRZc2dbjm6yo/HI0rrpXK1Q0E8iTF0HYbmAZl8FVTGsOt/CBhe8I2IZ
JzNpNP/aG6rnopzt0qm1JWShlG4XUv7Ix3LPp1z1UFnvxXmavD0lu5fTDkarxlfs
grv9AXq52zEUzQJ3Oc3g4PcmKeNzG1n3ci+cwAt1J0xBnmO2BZ+nDU2gXNxSq8od
BlBqRJYN3w2si7Z74ioz+nh6IHJp2us7WrtM53t7YBhz+xFoocQrpfNALhyTEguJ
tTB6a2ufleh1rN06JaBg3uLzUFqAcz6qOvPzDPpA9cautvQMFN/sfqdSGbS55Lvu
5oONMgVbd/p1VYmRufL6KSI3OAr95+W1FuTRBL8Gk3gc/hc2yoWk2y0SzyM0m8IH
2upE5VnhKR/BID7MaDGcsn5CWsll3Uz1BO9TeyPSk6NvfX1rUYQdPmRXsdnk1yzK
H/v5GKcYtD2LkNxc8xfpEll7Wc8g0CM0rvoscOPo104/d+R6r3zYdk75EGXvZU/a
Imr1bwjg3PYHP1VKBDSN0f1wGvttXqSRsDN1QoDl/7YsT7xCCjUw6NxU44I+4s5r
jINEejryq6T2eRUu6kLsYS0rBx9uDLMZS/lQJE8FXrZv7RlfRMFTf08sYTod7sT+
54uUnkzSGC+qqDbzpu5uF9HDt44DbkDQQNnGg0vPM88U7ovy1fcPmvF1xy6C97Og
DtK3uTmcJxhF9IvCEKDlHoD8nkWAJOslLiyCOaKt1C7QgdyX9pZ5qsCNenmpZ4tm
ZnUynShxXla19QUsl/C4jVF9Ymch3GCbo3a1CMVvIf4t3g6VmF+EUdcKlaoMLt0z
/yUtue8wb5rD0FGgZ2rSjj6w0eL6TKsSPZ7K93tyWqdSVbc5I6Bt0q7jmur2n/uq
QfaB//LNNfDCk1k3OOtmSlUd/NhI3OPIm8Qgdk92p+/SbfT7lCbLjg6wlIp9F3AU
49zcQ/9Gyh1eeP+rLPC/IvYSpVu0XOdUTenkildtK2J1s/7bC/x7CviAHPLc4WcL
/fgMMrbaCljhyKSV7IXP4Tp0EBOKIa2BVP3u0xJqT8GpZvzDGE0xjsoD2FBcpybQ
blucywafO+OXqCH9qmVVkNvm6gxEDgk+ucUSXDbE/h8PZ5IS+7aKIrIcMjOwfQ2S
bfnYESJGDdgLsgVrqwXE6vhNPq9oy4RjF9hwINOr56eCJsVg1ZMDsyhokXplgyy3
R+TNMopD1n0B7SuUayOcoN8uKLFcUKnOxHklR3SAfrqD9TDaJsNlubCM4PCcGqKS
3szc2BBw/wUKB/I342sYiAadHFe9kf1RwJ/bJXwM4mPUm3RiL9ICYMNNulEZ6IQs
Dc8esvjcgPb8S3G0OnRXEDnb79fE5ICHR2E/Qv/G/XF7BoCPBp+J8IC2tWQnQZnO
uQk8YGYXPnuWGDRZIHheUIs3SuwQwlwYFab1r2+u+6OugLn6aqHgRQ4irXECxOc4
JhbHgXB8UloL/ib9sAMbBMoOZUTJT0D7R6Lvn9msCtaUqAZhWp5tq80iZZFXAK1S
y2a6q3RKcHWl7wZa2oGGGvqK4FfgV0o2Ccgz5+YyHKCAc1MQpvp05EBoGcg6nLQv
SKIXcc9nD8ir2/iVWPufKT/q8NeSIIu+Bg+xh3aHe1w851NyaSebixj3mnuXaUzH
voq1nDRS2wI1WAV9ypn1x4ru9qcY8j5ax6EHqVTR+CRm3ylpJpnFaYAoJeCaTtzz
5i8aGHitx+i00mrsEKsoEFcvJXfBNHeT6CnczECRsgipoTZTXYNDuOg/vdlgQghi
Hmmek9kf+Zb+M8hVD6DkO2wudfI9iJqQJ/o6V//or1Q=
`protect END_PROTECTED

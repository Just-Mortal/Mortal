`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sPyRgPYxAoBQ6d9SxxkJyOQOLiPsML6clkq66au8s7SiHgnvBpjtqQg1SDhs6A4v
vTC4xv9N9pi2KuREbEpbIZXM7G5TtO2XlpA8dAkqtJgU8V4+wUF7TglmgvI7EYHb
bM8RbE+wBQ2YBEAwhh4AzKE4loOwau8g9xIwIM9/5/k07uNnLMCotcqVgwvqtf11
cDKYq2k+bMA+x2RVwwbMao2M9eh5SclpLRtAcY4aEw051z4Kz0ZS0Mb53iD2LCc+
4jlH7Rt0obWhekj3BPWq/EuKwhk02FO03Aln7fRyKbxE9ND2kVGVqwRwFXfcHwot
EGScBNOIaUe9SU1pY4hpWnkd3gqdbDbo2yp/t0Id5D36Qhs1sh+hUfUu5jSnVbyE
ThYlP8TgQ1FOYcHM2w/gYZ5CG2zvTrHCTMXO745AGjQoldoNnhzMKb++4HPVu7Yy
pjG34dM7aOl4DM1MS2aoaTw+18L6BGAeh5u3fS4zE29O7X1+Mhv8hEpYzwL8ZYEy
XOelSr1h3igG+jnnPVG/XA==
`protect END_PROTECTED

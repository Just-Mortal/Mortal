`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zoNTMk2+Pe2XzH0akOuXrniEUFyGwpWQrSF7Dnwseo1IfabR3fQ8cf8IRLYfow7a
85dAFO7XVRHZ10EGIboqEUYgX1/A5ZdFyDR8P0jHBokL5m86gGNLsqr2GZVLjmdL
0hL4nWGx2oINiKz+LSDH5hCThOvCFVqn9WTowkAxJi+CY7XTHWUoimaFDo1kpoc1
tRrAnmiboPZWcHQQUx8wKNgQIDGdXidOKH8Y6RGzJtvVeLl0h89NaGcU7j7rGkbl
41D+rEKUzZ0XkqNVc7N5YPfHW/4VH46lio7W2DChmT2PoUJRaIRIz2wmJXhOCV2l
R5wqPvS8MF4rxmca1gYsuFDAEGsCQagznPZbNVcce1qe939LauVsnhR7VXL7+/O7
OsumBfDNZp7zUHA7cmFxuB9tj7XallB4VDH6EwHO1gNzx1BAOf4LDGvH2K9Hyhi0
o5qRx8q4ECEJWLebo6nk6Roo5TpaO5I95KR3MW6K2kn3knekKjyU5gGJY7nOhVuN
jY781TZisvyD+tckZgs4Ip9gRvb0y2/ro75Bq/qhCzR8f5xgFE2mUwM3HWmYuYd1
tNrbuhZWkc0kp9kB741qisEsevOW8iiJQwqzWLfWhsDVvmJd9QuVBOW2daEA/XHs
vMcdlL/Hbg31utJYPrFbUw5MRj+lCkW1BROdmE2vcxC8zzTKoXX08gDvotbinilU
`protect END_PROTECTED

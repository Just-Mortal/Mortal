`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ES/6+c1tGoWbFtlMVjTiQBY93D83OI4LgGpVvWNiugD+Gf8YiII8BSRHQJqjew4P
KLiu1zniQdT5q4j/wVPhJo4uWWD8pUQuxs4jC+8LSPu9AQ0bhtPH0E7dfGl4b62C
RjJjTjsG3vgW9QzrTfzJ7qV4a7X3kZbJYEkT9MzvyO7gZa/eIlTKx5YwpJMUNx+/
ekxLqBQasrVl4Y0yHfDzu/vgrroYJQU7qshQkNvIAmlNUfvReVOeIP9ou4z8rHWX
g3daUQ2sJtdRriPONnIUlFt/XCqJE3pn3DMEb6hdo/U+K/34SBV4KU60j0cO7oGN
jzEIS9k9CHx6i8XKO3lzqWNXmaCnQavkclopUXnHX/3wgKF5qTchLtDUoRjK9P0v
3TjLI9s0+d33b/wXYgD76D+LGo+nStVOqUeCvCJLp11E61DH8Xn7Z+oTaF5L6yX7
ohqtl9XN53cFahOPYqVfFUXzYfaxlCttEA0KgSESrrzTW9G6AkW6qNn9eBjovuMn
V/9GtLtlW5zXBOBYlVgY1+B+Msv7qGqMGJ/6sFJTlX1xXjz3Ft5q+M/XFrv5uKfu
O7Ouw2/ZAyyiWrCA1h7usuY1GpQbxdQSnavVeaMuw9RQe6m4gTTKL8FHg0r4Uz4y
9pRWhtRARHOi8dG7+p6i9i+kcHBWFEzoMmDym5XITY8rUzTLLcZcwEz5JhAKrbNe
lE8DEVsiSgpRQkyxCgEBESHARROSM1lB7A8NjZ/4JigsQOvSQxUYAnRJVmYcW2UF
bp9Y13gW4V4deEwJH6tJs1q9uTNoYRbyIZJAPSwmppJCuWOrOlTYpzUojh0ONvsf
Np9eEM7Hw8jwqpFU755SaE2aEBukmZaoRFL9ErIARC8Qe/1D9ylzekFWRKB6ccKU
VBBd00Kg+pd483Xr6W7C9qiyZkCV9J0Tckpebd6892pmsbeNrt0FSPVJyxxxn81B
t+uXYemuc/Vn5ynLXhieWuEsgBHp6p1Cd4nX44QNTHTkEKnN3WY0idF4GXYcGD9i
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxuw62f1iUCAjndepwNV6nGpXdv2VndnzefKCyraZ9Oh/MCzDWuTtv/QnpLV5S27
lh75XcUfJVN2sHB36IjG+pFIRdddoN/K2lLx+Ls9uypGTrZkdOENGNOaqDssV3bY
SpXOqRifTG12o1c8BVFbR59Imd0OznGmZfesxf3N/+7PMqlYFxvqltoeQVfqkWEn
PBCKfKFgFDUv0QV6MFPzy8VjxRwVh76fKMdF//tt1u2oeZyZHinkcXcYszfqHhvX
twMEabUCB3JznnTQGX53qnYOw35gNhsjc6qg+mkNIw8Net4nSw2UdEQILLOAvGMn
ltYUiWQEgnBi21PylabCixJeh2XnrCc3aaEIU/j/DvBeCJo570kXY7FzpP6MpxTJ
pkOrmQlG0PLrNV44Mea7ibylB3DSik+JXWVlB86E2gpNyyzUATUJuJxirHRBjNpF
T3CpDJh5Ar4pVuFiKnYIam2QLvH0yCa5Ggjs75piQn8OHL/5ZjPfPxco6Tn9IrfJ
gQtDrIU/McW3HimQWI3+dB5FNKvQs290yL9lQjqoujdqRjsCHmPPjTqaXqwYuvvK
BbhrECeRIcDfA/AwppuKKlJ0/DhWyJBVe8C5emiUJoIgMOh8OiB9fHGRzPNAbPBJ
+eBLgkktne37KThOwBVTdbKNIgYKhUXHloCx6y+k8E5MPew1Fo1ICPKK2eQf9VyY
b8ljYhFWSYnRCdFBazIZhRYc0lTK+VjziZu75ZJktcIwfqtg6eYEiMkiOhrvOssh
0bPUFHAExQ6QcfO6xukullYjrb/laYfNZA5dnrLQHt+ffwXOMUGJnxzwdpYPliXx
X5xG1Pd122crBneIGN9PefaaLxpzHzbYbrDTuU2lUYxtGNSwB9G+eo/rWnlEu5NA
0edwkB/izRpq/FQf9kw3cDzz/o9IRgH5aAqs+vTKx4Slhhbeonyg3Hr6XH0YpMJ5
aP9k85o8nwdWMuQZxDzqXu5b86NhsH5pKyEDNFyUAV7sYyb1LIJ1UFIg3cgZAYqI
0Iqb5TrwVRb0nlgW8jMeNTcvRvSMW7yDQjOiJlOmqBeW/P4OCV3ldTzFEzPFJev1
vDIu5FWH4Hy09j+7NGDSTHXb9pjChsS8hbuF/Kg29zZWN6AqkMTF7H5YaOIVHgb4
+H2hz/LPnL51GqsKlaFbfo5L6+/3WNR7TP4SYK/Dp2bR+onUZzvR3vEyd3VGlNCl
MvxGFlqS8Lwj0YjXHuzz19pDeSYajOMGXJr90ai/d0Uv4fIsEh8aShMojUEXv4HI
b9XPjOdbUfPBpkSePF8aMPySiC4Qzg4H8iyokpYzKwYa8tGU5tkyFfFOCkVJ31Wt
3RcS81SoO/Hd1EQWXxbuY7io7bUfcYiW9+e7BzvwKIEMLATDIlMms7I13sI94wYD
rHGLoQW302wPFxuIAfH7Fyr9NiFDxQ+FQk7hj5rrmVyJcIjo+f/OcgSikcYyrw1Q
Gmvn1hqZ7iNqAzAaIMycD0J2l71uH2dKQb1KvhofEbQ1qbXyqNlvimflSFc5UVHF
fPM9Au8RtrmVCe4ZrLXABLHBRkoHPr+ztwMGg10BH6JVYXMtuVh70NDUS5OzjQEx
V5HXwU1+4Njk6tpzPdYgS0qzIINhN+cn6AW7ks7AT9Ea7ux7PeX8xRBxrQPZBBWE
i7Bl3Rq1AusWTPL6wR/PAAkXzO3TMLUQolLkb6VhoypfSxduAjKtDrXwrgZZ0Ptm
nhsUIHQwCfCMVr8HxRUTOwitAWNyhLKaEbmAuyFQM2qaiMvFjHgxOPdAgxPzxW8y
56sFmZJv0XUF6YodrnSMJEoUUWT+lI+avlNogb8rVFLaSsi1rGQm7uuD0wOjD9zP
TsRxALnB2Jbw+v3Rx4c64igiJ8tZtenLUUzhetgb4Kvd7E/IrlQxaD8nZ5OH7j7a
cbtrPE0WiBQq2oVgEDlSyKV2ytCgEP6XcUssMEydSnnvJNicJE2MwObTuKtrCPy7
NERw2YmMeqGXUoR3EFVtk2uYYinYMvPII+9Q7eJlHzhVCMyX9wjkCDZTsLJxh4Zf
1D9LMwUf0Jexry7pXPt2qpe+a5zf12voraUEyI6yBhyeKuhmoGmT/EaDSfrY+EdH
AxI82DWYAXfM6HCCuMP7jl2j/Gig+T8uc4WV38IFPKzrN5ODbEibGBOCDizIjgPn
WyJLmg/sMSDFnbwNYBIwAo0B1gWcqcjbg8zIVEiR8TvI1eKQPnRMIkQYV2Uxkz1V
QDXeQBhVV+eB+VxkPRUKSPRHNLwG32QtR2S+mlI473FdcYheeo9N1ylUl2e/As02
OmLt8iIyZ/XZY0iwVPcuLmoYQ1w0+1riGl1Rqr+43WTv4mzeHbYe6qAUEUL1aKbX
u6AbLMZUskbyXhaeQ3vLOuoYk+niTotVQSQx8syjVsYnF0k484H1n2cnyf3EuIZe
t95krN36SS46DbYV5QRoLnbm80O9DqhXL1UbYPteJc0Wk1+Ktn1pTrFJjP31nD3e
u3NEzxWuQbxrZIsvWuMs3DH2Pyuj17fwlnvKVAPmHocItNBWGGApdTOoQYqxruNN
ypzQNwlpIC1XBtwaf8XKbOhWjvmwFUGvAiudf+jdv4hW10F88y8okOvu+PdxJmZ5
CP/SwOhi0PeKB8LWhgR8ueF1s7NhcTIEY8fZ7q0zA2SGzj0AIcknePqYriRM88aq
jncOtnOH9rGoAnjR+lR8SZD/sOHDe5Jpnqfr+6NpyPMKx0JF+g/ZuhIqCa2gYgSF
qQpuS3tLe+3r4uLcdgU4MNALz3Ik9g8w+cSD0KEbUo0auVL5Lq2F50CbP0OtO0lj
6kuOQt7rahWLmgDGSLTTAQfyZFy0fdHs9KJgTOxSM0sf0Cvhd4lWB4HHNQqZpSKM
coAdjpsR3pSq+OrfIJQt6B/XiNEGOJS2+nXyTi9W9dSA2inVHVFwfd5WrTqqXQgy
U9V5nazrUCFhLGk/1dkbBEF2SV6nHcZtQxMWq1zqQRD27m0DSVZEJweN0me3lp+o
FCGSAmQYVtqDhH1OsvUkaeuZgr2UI6amqI9mc5xQx8HCnBETAZxxTrc/jfwNHcXq
K4xvCX+oSrMnq7vVmYawyMW/xK3iGtEWJ1UHGzEhNG06W4e+OGFKzrQy9YdG3OGN
EeYfRB4VrB2YnJ8QKlF6cBAT58xUjUEFN+XV8h/DDwArthAuEIIEKMv1MRShXGu8
wWtIdaproqERKOR7byEu2YX3buzHjbF2VqYAubtD4w5rDaoJc/pdmu7KWh2qYsHM
B5GSMFeunUyJ8YQIdRIVftNbaQzA1ZZl5RSiWWXOHyHH2sOCaRN0/X+l6Qs54OSr
nQgNwo4t3EAwvpccizNJhe8s5xnGcIDT43/TIIfWIvFUNfpOzOB1w1pUESGxVdUB
deDnZSiwKIHyscupyyuVQGnOnbg275HOS5N3DEuz2MxU4bDtkRQg7ewmVdkuvZvi
xURgxpTrwNoQ4O3UgjfnyDMGcECilH2MBQoWpGUzkGv0gSXalMBemG2DEYSYC5xA
RpTTAdyuyKtHH45PbfIzdZMk85zQ6R0Ugp2C0y+VFmo6lIDDhI5W2D45rq+1aZaZ
6eoZioJGKO53/+voT2vyl7Sr4ie0uwSS+zW9rr+L5Ll83UC6R0/Y7/omYTUyYZCW
KNfzvCYbcvSlOPu4pJwHhWiPksLRij9OB8cA5q4EsW/LwollbpEAE4e6Hp3hv7sm
MAw3XvkKhI2R0WigYTuFi9RsU9eip/zUOrldndC8rFytVoiQVHmh/PxwDicmNY0l
vpzwckRN8CPo1fPDMubZ1Mm7keEyI5GKsHyzzaV8rJ0bh3UnRpYbJJOfU+MP6Y+M
2kBMwnebCWo3bVALwEIrg2oy5PqCqVZaP7I/7AXjo3VVKv5AMjEtRbxyzY6eaSHj
32PmxJIcU5zHbmBBkz9kEoR/iNmJL9umB13g6+jK0h3dd+gmDiU96fl7Aanp2nZi
gvRnEl4AETNXuWrGIdHfoJ4uX7wiiX8kA6etxp9s3hu9hpHaZdZn41lbY3g2RQXF
wgPef85PDB0liow2S6uA6/colusSl2QWJBhvHWEyKvgs/QK8aTgIXeUenuoXI3n6
QqQxgQurfQXzUU/p6kwxTL7wIn1tGrGz7mXbqVzOrLW9FFOYzqp31xev/G2KJqlu
1R9w3i3FVFJRbvd5rKSwDPUgmO7RppOAPymcOvMuZ2SYFOb9uRGJYEIwQzMe71eo
PGMJoVVE4Azx14mq/y8LmHuMIC3c/zmG/wElyEJDFQavwYA7SrwKWE0m4geT11BM
83wZzIo31GD+Qi9IjklTSBojcxveZM8uIwo4STdcs5cj6Wy8cJQgs30coUhvsaYT
okENlSMkTvUiGaZ9ts6o2Z977WA/vRbdAIVdYWSaJLrOZTRW3lWrLpEvEUotTAv6
5xfld4vRwA2m1952f2L+bBHn/31bVEcNKoWk++3LZMt/1RlXIiOy43aBmVCRAuJR
Bv0MIZNrqjvJrczfPxP/3HankgTbVFdAVNE9pL2ueN4Q6X9Xr+V+7aSBpf0N33HV
0e83yGb4xNOlrVJrmo8W9pBt9RznOYbGqjvyjQIrOM22Ri9Z0xVV5qh/h5iTISYf
/K4OYQ/DdeXd9mO4Sbq8ZrqOLYsMKW+3wJNWBSQKBiTXCXGHbRRU3rtWeLomgTQq
ZJGEnWgB4GpKLNF8l3x4uxqMSf2vZTGfy6Vonhua5gAaoTaG8SoKRyjHpxJlByIG
3jZYIoT+8Isdm7DxPg1JIIayH6lzAQd1FupIkGjUL5xJIV4w1pmjgsbM6sA8ac9n
RFDtMxV0HhGATOpLv3KcCan3ZUVppcAPH5oa575jGuF/r/VKpp7NzqhAzDCQ7oaW
OgMPxojV/FGg9odgYOGMxB+Mp2U2vdqxmx0xaskGYOy1HNlffpujtb/N0XoeiFxY
d5DxwrGj2LupqzfY2+t2Z+OxYYrA0nn/ECjK8NKDh1GjqqriRHhvPvZvTMDUcsx1
sfNzMxu9WipvIUyw8Edq0Kmd91jOapJ6kEFPiFyh2R1vpMtrbuZMi52fGara/kAC
cAjNtdGejiyScPpjaIapivL/vL/BEDSJ50LUaSYC07a2yfcrzKoeLHKRPkdOytZ4
OMPgqABV1QR2n8WBhcYD+wJuWApAD6Gmc0d8Jxgm3AZfYXBfxTyNDLHnk6Eayby4
TiUa7SyY++WE+zrS2UjD7EVymzMf3e4f5lGJyjk9Uj/iGLXitu6LuItanIIPKyXh
nGEFx61mjiFpI4c/AVjzddtIJ5SapK9k2kuEK72jNFe6Cuz04LLnaKCNhvvs8YpS
rk5OPzu6B37NLt/iuy90gfiOJkkymhghEtfoEnknbjwYjyCFWeE/+MNy/WEzrNzC
xrR9HmNEHsm3GHJMGuK08qPmCn/QJk8jGQ5yeAatvFlyXRKpH4q/8eyciF+O7OIi
3LNp32Q6dOu3AN8FEQvjO+/87qgGfEZ4TdIB3MYpBKy1FnLX03ueF9RzTVr79B3B
zM5IAdTgX3oNPa5q172Fi+awO0hHaote/up6wV0+HogDPQy+e+Rb0IYmokTedMJ6
wCXZmO0dEEE77cmZqs+HItWZMHzopiqTh0o2br8f5wb6KXc0pJCnpwEe49S9xqfW
NtJcA8+Hahll+fQHD6hezDPnrru4X2T8ht8Gn8zW0stepjI8QaGyRHpNW6f9JZwu
/6emgkKmgkSbCfzgG9g3N0SV3TAzX8G0XQhEw+s4Kfglq4nge2ZFzWIecHkJhNmY
yBUD6s4v4yf5FkILltN4u/Z03Zu6t0lBh051FoNPLYGwwRW70SrcD7mIxQQpNhqG
AsALr12ENOsydFeUVXLJJSOUHSQ5hVD9FXvkHQdpRuVy3tL1XdnzHmfHMsoGqIp/
aPsmW8hclo4q3HjpqDrJmm0b3QvVi4K85/ggnYksrMpWwc2i5nYWB6C2DMoIWW1n
YdEmdBOPtFZ3FgsUxU2jBIR8YUctjQc2bhtGOpjMWu/XgLz+CRJYaYsL1rFFSdmL
uxpmi0s2lflzMjD/aY99qGPXMyOSb7054l01H0qdEyb49UCILd8HSUQijRab2snN
rwSOfFA1aFOSqBGp91AQPx/B/iKf8W9o23Z/VOOozcRLeDlYKMIeKgY5QIS/nzdJ
9dQQ3AhD4iIzUzaIANzooHRiDyNCq0Hubvye08+A0AySSe1iAB+Pi5E0iR6nOquY
Ao+TRd0RHpgGYJy5fMRZQVMppSFpswx/lJa4I7t+ABswc2euiw3fDvXT/NZgsrEH
GkhlJW1E7L48RG/uEaKbBeiaKaOzytJ8CSX459MC4Ud4GwHdc9yHDDgDf8RPYi67
D7JdxtxR8qjCaWMd4Oo5tfnLkxkhGqOMKPSuI0Von7N1s3Tl986u9J2mJ/gSwLoy
8t6SesBTbqimFYutv81ehUPHuyQcjP1UtnNwOSshM/h0CfReiPVBi7snyED3f+/T
BHm9rEF60AH6kEHuhGxtwmQrjUjLWJF8N15dZYvoKQwLBz1u85WveiqXnLy1VNmr
hfwEUMF4DMjADIAqyvANuiAFPY+tkXoxFYSpmGTWv4JlwvjQjbUZ+bkqgyc9REOa
Z5F091kle5wvNrFBaMdlGFjv0xxYTfR5EvVdJ5OLevB6KsEe4PQZPPIaWKpTh5i4
JmRw3TcfZJkXwvbigHgcSd5FmfzoofHAb3+6dMneMbuftuxWw/+mXBdIM1JA0oFc
l1CssRQCTXz+mIPhcw0HEo/lWr4KFbaMxXmcadvbvjx8qa33HKAl8RVQb1AN9gld
QN87KkgU62UITo5E6PL3ZlUIiQFqZDBagXS6XhZt+qkksN/Deh69wKr4vC/h7w8b
E4TsqLYDzIpWeG3oDFGsY+LwFsbwI0CK+RAGYvPx569fWoa055UZFiQBNN5ptJbW
YtaOv5xOdq9FYLqGm80it3oWUPwH63vhCwVyjYVUZyVbvokEp7eENhFJUTdNAmri
P7q6mu3vSKjkqshNNv5tokgpD78NetzLFOGPvMB66HlcKuIbknsBVQLFwh4KEd5h
hbZvvcPYxm1wrSuuGeR5QIIs1GFnlshG6T/OzOCdQCwAcM/WoosGtsLJ9RruE5X3
LdHdlOXjGmcF7VDftO8384jhzg5urZ3YGGiCRBU0w2yfZGSyhPP5Grfj5rHPxDbZ
JYCOnWAJnW26il0tgjfP5kvmbu2gZq6voVxs+9+2W4qP7Xn1PL2bVMRQEaqv92f+
P5FgAG0U+e2KsusZB36/EfsR0TpYt1tzIhlOexcnZCZAKDTbWJ1i4WsL9j5e20gP
L8WDHy2w9DH2yDa6/DZyKW1paXahSXE7oPIxjRSQhpzb0twk5D7xP+qeFinAeBKE
SZJybCwQWhWMaIXx2e1H3TCgTO2zmOEb2SUPXeePLDOVGnhUwsFKehwEClprZV0I
maJPBla2tCFkPjdRKMGjE16lqf0FXe4/wwuG6VSfbU0FvGIky6y7KMZeOP3DCx1z
Uw9W/MgeHRH8QPp6w/U3ZnJslxJs9koXsElqfbKS82OapRVga06/7W+ovmrxQ+cY
e09yv0eLxOqXNDOmnacdFBpeHq77gz7IHeXFCpvM67+STuwXSr/LNYkySPxleFrJ
2luD807iyet8XEP4ln2TRkWW72rp6wT43cNvwNfHMCd+vToQ98MWczNIBBdQmDxf
G/NaCcrfRE7yU+6pH+590v39Cp5knBYw3/O5KxvyHsocCeZptGAARe5oxnvrJ/Ck
SX+LY/NSlww8SGOLVg3U2zE/7aSrbhv6hXYTQ7BuQO55qCXmspBuGLbfJMSxa9xd
XdgwkiHzjdAAbk5rtP/P4d+XE7J7bq14af/TyjeozcBkFW0yfHv80KrQCvvdvjs9
AGLwlVuV47NezR/mjMndtG2Qwq8n0ufNoY58lWRAFzslFXVRj6NvD/JhNx7Yyrp5
i9lgVIr7AW3l6jneWvcVAab7ULPBdJ3dP6jye8tgcpBjhcp1OZW5UasTwnqHH1Jn
armvA7OxgQlU6XGMPcONIxFWzKr8jdE7QxGub/gFSQk1rMhpD0lHMZH6mG7KkA5w
QCMnl/x328jKY8xRpQ7X/YQGY8Jb8QfKYE721iJA3SSkGXXJy8AWesb4u1W0ysij
eCykErlA8TpG/vJp3Zq70TCRiHfsISjNxZz5XzozVTfmjRKMHmgjHqyrC2IxafFW
+4Y3RJzfkYrgULgnqLqGMK2mtMQozcwVYckWy5UBw7BtqQF9UFEkmR/UCNcGbnN0
7wnxlEXB6sXey2HvW0rUWH4nj7S6tIEiXvhdBzvRyG6vXdoKTCThMaTeGpRNZTLX
7XCi4reP1j0YwKIwx+uZsf0Qc13Fg7xvtVwJ11PMl6O+rruT8rYr8bj/P8BFGPDH
Zzb3/r3P9KC2LqNKEIfeWiU7c3aYxLhBDNRyTOUpsusLQIXwKCqY6nRpfVp+wwCd
5o30DheQhPFmLyGxnud+GCaxg5fxlyYolLKSPXvcvrhPScRfh9WcjiY0NIUrzAVd
zWu/PhDWLWA5+r7Gme9vSWzEHQWbNcPqXguV9y/jNlgg5Znts3kU2Y4JmPkGIv+Q
zNVfBytGRwxrnI8WzXQFFSIPyQigJy06BZE1Xlgbz+aWy/ozCwZwEKbZX3dqjIAr
5CgKpMuyYIKZbn8hH56gMqhk5exYdkfjTiLpUVOXJzQChEvsdJ+D2hZTYbS9FPG7
QsSZImclLMbpGQbrWbu8fbL5oDrc+g5eRKDgwSdQT/ENS97IsGHUQKlBj0ifahNt
Qgn7z2hGC2jZTlY7f3VeFUc+eD3uEsM00L/EDNOk6dGUV7z8S1QNehok0IxywikJ
c1u4T9vD4t3FugpHjFVn54WWqXdA0iHqx2xLgrhbIRmimrHwtDLITOSXVXJ/fwxi
sDzZ9KZDwduZxaLE3jE0P+h+7vSFRBYrvZgBEIUD8tssC6CX/DY2XFikqS3dcs2h
1AYU95i1BoTZ+0GjBTg43BUWM7eztZhMgc4wch/ylJnqgw6+10uTwfUUrMnjM1rf
5+9FOFHuzg/ejub5ajxYdjMVoXFFDB1byheBCi3JsWRnaBdc+j/sE86WpOwW9KdL
50ezasDG/xE71WBncZCXi5vNeIxJqT5EF+Oatna4BKc/X4X2FXAtNt1BCKHLM5nr
RLeKpZDOLC4RUkg4i/kuIibS5+WnxCbtlHD9V14HzBL6fYdhUIogXrZeOLqI8+OT
bPMpJRBZ/mVqT0Mv/+E02B8IZs9odRsu6woM80+9PcIUl36bUriTzeBVq1z15DE7
erlPhp/lJwqi5HhLGmOAwzFKWhQJ9HmM+vTe8nQnNFet6rfhd1PpU9K55SkyQTiM
AKOZ2w8zvRhwlSTCN9JcicYhIImsBacbYN/R9DZq+/0W/RDxOPFz53NSp3q49fji
GI/5kv5K8mk7bXqmNRw3Wg91muhwbUKA7WXuUichOl6NgWBy6VyyPwohm0Tdv9iJ
t5XdRZFnEbsHTwYtl8M7AbKcep5mU6fgq644xPEC15rHG2k+tZ2Fyc2wV9Fus6fK
iUC1HYqnGW54w88bwelG249AhPP2U3y9QE3EjZoaBOw8abjD31cq+Tj4BSMN72zN
sXw5P0UJOS5m/xDeo3Ff0OiX8fh5wM8MW1C9I3oLKOC7S0M7ca0kMRDlqOwErh9X
BEwXWFWwfSXDUJTjWrqsztJ3CWuP0ASqE8KBfgdNzjcRPPOPrpXVlwj6BLYNGay7
owXVRN3hzLHcRPWvpiwgunO2fxpFF3O4t3pJGBF24X+wbIl8OIIZHxnU4o0UNPb9
t4Wne1SrYBilgEW4/cVwrzXk81Z7jOyiGyKtp3mha1218rbi0Nb7f2Kw7huau7eY
csmvZRn1zKUlHYAVRtysrlSIh3ReZU4v3l3tNFD3qyHEf6JhcWNC/LsKX/Ri8aCk
yoQ+LFzbdo1II8pzwjye4ExHkQHwb3bG/RqpOG5b07ju4Xew3Mt5u8hnM6rfDf4+
sz3esHrPBpIwVSUFtrRk4G6dbfsxyWFgXFSVimz2SRchQC/gs8MSBeSX3Uyd5QrP
yFE6ITQfQ3rd3qWA7Q7V781z22lZPcxN2QEIpcBBGv4FI1AIvl3LOjhMZIPR28fT
jSYYY56+OHJla8vkhsRbGxwgVUVqnHrqYJCJ5iktOqQ7HOJQGHDflQaFDj56KhPx
txBOWH6pOUnBw/ydY7O5jiK7Sx+O54R1f8sd+Qn96dWHWARpd20MK/Hk68XcLA77
dvXbFPce508V2JgfpxQ0Y/1UapytT5m3l4E5hiXVWnombXus6j1yp2BcOoH3/zqd
KEUdz0gzHufc8t0adsH8SG5YQd9NMta4kDK+Wu6hLSkp/Yz/D7bP5xYuIhItJdwz
FGte4uOA95YpHir2d5MqhCRj8T0dMYzSKeCdsjadZv78TBEiFAs2vXnvxn6gCRHP
/KIKo7eyM021k6f3NOc067yoO46R+emAkk6K9GIsl5uhFzPtUW3YSLu4tV5gpWan
4KRCtl+Ii34WJY4+UPducrQgNDc+kLxgxssncNl48BxyDJL8NnOqYA2ChY1Yir3i
VH/d+eSHsiCoOlKSOr7rM50HHivE/xMwsPR/+95K50Sa3LJyJcKQt/nzeQth+/Xu
dV4V5N/cV2/+HgiPPKrubqshbXOTWGFu+bmb4tMYXW/D+hDBx3Aq/H+oAtOMEV98
7yZPJlq6/NV/sfdUace2N/0S9CUo2piB0V6Y65J5byFkT2aIf1h3AsZUB0HSOKSV
Eyqz8jyiuXi53cngfVR+GvydLz1rq+Zzgrp3Hm4rad3eZVRd/S1W9Enm5E1DQULZ
DPVVXwzCmAm6v0skdWyCDePAnMWMilCgnOJoDmdxD/dH22ZG8VGnO+Ou4JwjEkb9
qANG6BcjtajAEJyNiHn6pbJcVlZwfu97SpOzYUPSqyitfxAU2dI0mfooZ7GsjMPI
SQhqdIwZ0xKheqIfXnjLnIywfJIdt6p8vx9BzVeHi9jvtCH3qajJWv2iF7W7Suws
/ZmB7HTKDzrIZ+OIM6s6J4HrzUZsph/65bmWbNdXYLwEnALg9aZhYCTNaRVqUdfk
PyO6DKjhHdjMKSg3MhdXsarFRb+Su3r0J/01sGtn+oE7JSzPC/Zc9/2lrF8rGON0
xDnX3CVhk7iNPJE5P3zS4vqYdn3LyO6ATI1oUizZSFFbwU9nhqwVm/WLwxjBZr6W
ZqnUHGswPRoOwr/dVqM0BXi1zWf/u78aVjE9HX6l73sw5ryoYqw2EaIJIcUGKqIv
oPuWDdvkds+mFfcrLk9jzPx/xO0MDM+7omQ2ORL3HM9Ad75K8z7xYr2s1gas4rpz
Zl3A07corg5UrJcMpr59MRvE3G5ki0i+uuwrwDj8zKFCFt1qs/49qmK0ZAFusswv
oKBVyaOWXU3NiUHsKyxY6B1z3khY/CAaq7s/BiL/qQSeXcPEEfSkEkBVdxUbUjZj
UigtUYcENQ9hP99hlZUSkt+OF0NODZoD5H9277pXX8tcDPu59h4xPNeWAF7GRvhU
OK+5sWKhEDGtE1MMVOImDuWkVS+g5/YZZrn+y5kqHcMNIQgbRG57iqKQmgWo3W8w
UzET6cKVGzqYqaX+FpPVMTQ7T+cY/RFwOQvjtsW3J6AC3pC/jcXx6h5P9c6LGrSs
7MCIQfQqk4USZhpLIMWa/cJ8GwHFK/v9EDXL3cyhUzVA5zVZzWiUFFFvolJ2Phe6
IlzNaDE0+5Uzs5Nd1WMcE7bETmuQKABnSVA+Cz64Yxa23Nqym4OYkxFgXv2sXGBB
uqjW6e5XqySAYC6/vZ8OMtrW0tEMixCYsTwaS6tJHQHOTwwcdQQMeQ2KzHxPAv1h
faDnTI8lTrZTqMc88CNQM28nFMQ35kwBEpxvqkBXFLkPpxLYe9zsf5VVdgtqa5cN
AwKyUeWP1pZQO0n5Ink6OAzL4MSnCH5V33SbDHNfJ7BuQ0kijfPhTjOECLXP0UdT
3C40bEDX5uSl5HLXzYCIgCUKVCa2iBBrM7EB43muMZhpD5Vl9UHovLTGF6Rp7tvn
NKWbRP2sOD+eZZuMp+7cH3r8Yz5SxlZw7LQkscOH+dhnQwkAOkTvUSMFJV3k6FyP
hR2PdoMTdTLYZcS+Q6feVBgQtGOOwt5cUtK/9JDUKc8X1WyWBS1ZJJ/IxoKb0euN
a17iWJLVvNrZ5KloiHO6oTlYSmP365FdeihcE+vGRYMCbw7dR5xY2oCexTsc7mw3
rHUyKvHKxSDTe4XUkI4aLRYeZD1ioED+FerYdkwOizY6MsQrcY0L2fAqAbdmI/oW
E/veIqdSkFjNKSjqe0oE8/nuq+jq/2oWrc3Qh5tXfllKGEV/y6CWclRcqksoUYjN
IO833kPiJRtIud1cJ3OXcSNG5EWSRulnhH2QUOQ4yutDnR4ce08gAWNx2kehtFFY
7F9M75WmSbtxPLPT1nJU/iE8PoEWGPwxUHwwHBqtXR8L9YtaqCoEpcRw4v0v7+E9
pY8ALEoddBaX0iSVpOAIvL9QEo0j/ehBpVCCGL9DeMDvNoMbAsnbbUeJN6HL8nUu
LsV0k70EUisD5USlchDezhsmOswz/UmOPTtITL91jzwbXlaEuy/YBoqC6Rtdr35B
H5GoDS65tKk4ozGLKEJymq1RPB2q3F5CIRN5epyhMt5GMzHwfrFxTDWBAZjSbMa/
gtVttmzNL9pT+deAjayXmivyORJK4liewpL6NgytfJP3+zudu3QcZ/iLYWWutJKH
vPvrV0QlmDjy3zHBHFBVI2AXwuVWme6DJneptacYizRC1hUDOfXvhJqDU/zv9+Px
52W4XqACOAbzGnB8oeYWRdtIomw22j1Wr4+43Ga7L+YZor1gVBGE+lcVqywAsjQ2
SDZqJkRqBkhn0RbkWUkHqiDixTRbIz7edqjMoIut1BUKHToAUULinp9B7vs+Oqec
FTtow3M0u5m0maW/HSvlLXLhgo0uOuOqN2htwB5jcexcN6ZnWFESxpNpgc2/eH7x
T15/TX8CnZcRB+ajuNfW+HqCMu693IKraKQm5Hx53Dy+ShBmk38y3Km+5Hir7gAa
T/GtrMeAHbHf7iKfRikrpiUl7q4rR3EchkHfwYx870XIhJ5aVfDL54u1q97k96Wj
1g/M3bIeraY8vKUIoHKPXRcp4fUZ0G4UIrvEz+4hP6tfaDX5Q/hu3ITPHnsl8DBY
SZXe+iCK4RypRsXmsQ13eWLUHsamQJL+sbDQVKXPltSK7TzdwVse975oBKRPSSmy
/KSNQcxJGLj2Y6Hz6gwrzDSYMdcIcfqHJM60MeMY0MzRqP98uw7BGyfXYgWwghDe
d9mf2tKYE1Qf9il0eR6rSJWQ/nye35U7UwYgtzcnWhUb5X3T3ZCnth8aXj5d3llu
aCXoGMd5khrRQTJI7PNy9yVKMffVsJVrDoedtBpPJMIUiFKHnrNY5SiY0LbdL8r7
T+bBS7yYjFI9p6BnrNzsVlKcdO8fg6KUy0EWMjNp+hla9MVGuPRPtZZhGZp7SGB1
P9HS3Df3HlY0+NN3JYNrw8mHozAt5aY5wTOxMjBhUh4eIH+5viiflnFd56Bj566i
hoFWpjNH70EjVB3Fa1zbYf96dSlxh4YUcCQhieuJLq4Qji27hgKXhA4mXNpDOdAw
xC+z35V9cl1X4IaaHmFpCQ8kDpCWreF1Vtqpwhg7rONM2QB5SLgWl7JAoMl4kTpT
IGrXbaI1D9TPqiSVeVq8ZrrXHrEQ7+Na4dNi/nrzSKdNPBQZV60/a42UOIV9fvuD
ZLs02n+dM9l76ZoylH2/JcKkOG3UDv8rACbItzg3LuFQCn/+rz+voM0xK4nOVCEk
+5Hwc6fwj7GZpbk1rt8r3SREoERBH2JmTirIal6ONcupom4MOpy78Xfp3e93iZxb
N7i1+VLQ+Bon56KtW3nxdoNS3XVLRPxmwC6CYWdU/9ft6w89sNwydMuZHP5la5mX
l4Iu4p3M/RVBP70TrRfSC41A8G1wOONa2kHhOY+Oejiaq9AATtAzL8bgFYK8TGi/
aTezxa8paeafINTZLsStbCcxvB4HvnXfOQ2IHMgZW0v/Ehr3rtkqSifSotszRcB8
CnBL6QybtPTaQVB+q0Mxszod69DuCNs8+HRY/jEHEYD4DIlVLUvvNE9O9EPExz09
f1TxC3pzv80T9f9fsEN1DGwdPlW7kZwrZo0N15Azqk2PIla2lfIy+INpLpE/98RU
IDgluJZ36776Anp7425osR1befzdyI/guR2KzdkMEHxipJqFG0F8P8g5MsM7gTaB
MBvgsHZskWERf16XCRYgWxu65Dj7JbQ18Kfx39buJRl6QJy1bIHjnhfsGik6isDS
kh0fJ8DVdDbO7dSA8COE82UfwUqYF8zeSkh5TBQZje6j7+dDzAn/LpwL581jyxfl
tTLvJ+vCc1TxgacIfJpVAg18xDzDB/vKn+yBKS8LLRcRejXt3khiJdCGEzWw8kyd
GKZ8qBbC0Ci2slNYfLq506y0+WWD8Gkt4iCQmaj+xk32fcYKIGtzmWK8wvl37asA
dS0eoAEixGkBNMCJmDJDpP2g1hxTeP7dDikr1eXPvolm/W/jvD1MO4kTIC2ccB61
XML0F50SaIoCdleWZV2iSeDtokgi2oe5gHy6YAhiJGwZT06jn5E+lKOS16adKeeb
KOimQMukPkcx2ghhKCNF5hQWOda7HteoDZs0umU8Cu5w8zZtInQEVmwjUNuLabS+
MUEbdigqRjWDY12QHp9J7EVGDdEKzG7DBNRH1ymJgn061OhRScqRcmNhYP1DjiA3
BvgdwcpHUtZi45fgJweMB3uF+fWB8HpgDHniG+RYHNhbhW1sfccLwaDNRMS+qqHU
36/w8Ioo9UyWGA/OltiY1w==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7DQZNHA0r+OTug2+mnkn3cVNZ6+R79gJKzD4iJaFb0TfLIS0ban3kB28cGmf3tCU
dqW9cXM0bsL7nvzKm+MoZDC2bY3Hslc0pYSiR2bHM3U8d/3jv0WBepYWVjdAWIhr
l65zmbL2JGQNaHN5Ne/AcBF0x6ILmIYOHKInDiEwLIDW8JlyVZRlaxCKjnyX+nX4
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lurqeyYH4RVvlOhX2sWUFLeECiYtc0f48jtYTmSwF2UUgi6XVAnITKcyvbL7pJ5L
QdzaOZlcQc54BDNsh5MnbWVnifBwWlaL4N5XGrbXVkkJpfpIqINUZ6itf4z+Rdgy
NjtGuQrbg+JbuAiQRQHLBTmluuG57qA6Mdt+vn/2b/ld72oMbl2NKQ9VQ6V5xA28
GAdMR+6NGD1YtHZmw2To/NWW2HydJ37jt2UrKgFmXQ6umOJCPC0w2k4vep9shtNN
l5RClqquglNrCbfTDZV6hClSO1veFvokSYNQx3JA92lWoE3YNMr/qiOp8mWywQDZ
dhtfUBUjQA9bbNM72F9MWHqEFyM3yKjrerzHvcvz1Vmhr2iubO8nwAsS+HEqMCqj
P1VxNShmPTZydRUiK8lkwEjNvHh/AbNGgMSCazgcvfcgSX8/rz7lEbEM2CLQ2YFQ
p0N08n7FsrtNYJb3oJwRidLpsK5g7SMCUWhR3nOrHong03TzqA2L3R/sJBn6TdNF
+PvQvIR3dLXo7Krut5KCAcCALVhoaYw43Ke5R8QNKgSmgu2hLGlf/GrRCL8eD9ZS
lL+RVBFrHaAaqDKMXN/EsFjF1kGCBVR2lk4G16PMH00ACmLRdHFmr2FnkdHVKk9k
mc7wFgm0XVIiaK5dvs14TfweogmuLPy0/PC27Wudrmka5DZ3AvQlZAhSBfBrR/ts
lUGkSt0tbnT9SoJPf7LWhQFwx1V7lZiI9qk1L9yye89NiShH0iEbw0EuhlRN3a7d
d84YNCEBB20EfCtRSdauaL4/f6gFDswFwZDf3KqqIL/6+xngtk4CcV9gqnjFiVI/
oAlXxbj02fxYyDxwBbXJxGjU0CTIIKl1Pf3rFxXeyl9U0HDQTWvXwaqbESf0v29a
YlYK7303Yok9svcRwugMwGYGU5CbCK85IU048/qDsWLYsN56FH03mpoUNF9AkqyW
tsTgv1YGFqk11ib7TCz1VDbTqw3LydTJKnZT3y1nhHOKoan03fsHt+rwlckyM2S1
xcv/3XxyBCFfnl8r+I3U9+GYdNaD11ATtfeNtB3s3CwYSUecLM7uMTC1D1I/1arv
lMpjcKIvNDR3mdG5J1p9z/dmw2XKr3a97Ir3RqNoaW6sE9V6aO7dUQUANIA060mS
K/9Zs6PWsnfsZutbf5rON4rAAhiAqCA79BX/FWHxnQjN/qTS/5PP9+gONqm9tenQ
qAsWc1ER6eX7ehiFaO5P4kRHwv2Ps4AVt0vMQO6a2UMBCwFZFJwPd1Gg2/9KwQjM
+61UWeRWnu/mded2VYxTsYi0zek/UasnT1J0ah94KoEioeain9lEUoCWyCLdov8k
rkVO9RsI3F1roJ1VTPf5n3H95mMhvvaHwyvuSUx1t6hsmM++oq4v2DSapv35lmSl
ftriY3hINkyoJe3aZNNhfiLO6B3bJunnlzUFMxK4IBk=
`protect END_PROTECTED

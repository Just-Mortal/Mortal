`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c4gz2QT2OrMYWACn4TkFGZKIXGao/aEviP+iDv3EOOlJNNugPL1aEKJK+LTl8DU+
NDUN+GhdmRrE9DN8f04o1RnuYJV+Iswl307z0mEeWNubIsdRtkfrORJuRdquVzn0
5B46wLky0e1wrEFd23T74HuP2+g2DoY2tm/PVWQyplnJkVIkbKy6tgzeDXchbPMj
hSjV5E+ir5DHh7KvaQNHQAb5/0ntNKP6TzzjghRBLXhei2DwWXP3kNW7sfy7SZ8E
hb/OcKbXOSwbJX0yTSQ/UJPFN9BuxMmWSl5CO/Wv/WuLgnLoJ6q2RbYulWOI8Eb1
4XBo6ZyxQbKDvYTLs323RRgQuQ1/16vGwQyYHDZPj4kPZ5527+PZnanZs4JYqK6n
zjAvXIc6Nf2vxhuJ36yBqg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0Nzcuaf3vg638159LDlWHVDA3dtsG11ICDT1MofXsbvbOItPFjkf3/I+dDZp3UP
1f2JEoFOW9X/EJmI0fwxSbz1vQsMah9kkGYjjC2lrV5d5jBhSGgZZs0VF59ZRtsW
aDeujuofgQ6fpEzlCzyzPRK/2ZdZBisAa45AXfpR0CYMTN/G3whYAULwvMFS9Qk1
JyJhtWLlqVWL+ptZ+Ig/SIOMCPChPJTIaoP5WctPCBQJXluekTVCkeUCFuYGHkvW
+0X8i5Noe/zP3TJpV1kLLCSdPf1WQe5N0SgTaoGeoqRmqSGZBuF9m/tQ0pQnq5CX
YeZChlsmlRwS0rQLyNZ78nbr2Fsk7ilEctU2sff/HgKqagqjQN02EfCtZb6O1aOz
FytR+K1i0XBvoQm7QLhxKvixYRf8Bm51KHjm43mEdGSh44VQv6D7adaWeorDTYid
ins0CHI/cDIaXuGT7fDj0odelwrICfyyHbdTVOXWi7g=
`protect END_PROTECTED

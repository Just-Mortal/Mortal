`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HUb6Km9uRj3k2bzIgxbQAmjeeBbfnXYP0zKV3DPB6zXo476rit4oP7UmkkMBkPxK
rDlCv/51GjcreJiefm1H7cGST1VEb7646i8H36AFvMCul9vlpWI06/vrPrJ0KsTt
2CdFf4dM6G6gBbFouM14qV0fV26htitmqvZk1Zy6HkY8Sqi2nI88unzpmM8g8N1k
bN4iihbmHILmi1VSVGh41TKHyP7cWZEom+sqMEUikZGrjfgkkK3J8uyuXjOriTa/
72IUrDcd2Kir8nHs1pVuP2cku1oaJ+aeGXQW/LG2JM7/xDZEp5TqOO1RQ/D6H6z+
tVrTOfVlOT9BRFfWf3HqZ2l95I/n5BHoT1HLOKvc11gPWgeYAljITiufFVmff4oa
f18ajjKMvekykGa8o0yGGZXiJE82ZSZfy9RC/+ZbmRDs2IR6IczG0XW7wQBAVqfn
r97GkpL9ATWBnYwItgxZQHbzqAVjg5Ec2mLWakor6VzAYsX71HRUN9mz3Q+cZSmt
xCs6kvhPRR86lML+gSTg1lumkkqhk8LG+sVk1XNU6z3Dd61Q0CnNAyhhl0EGaPlK
WuBNYxV+gUCukhJpDfk6PjxjwRYn7siLCbJOj3oGV/PhhSuS46wRCdpUZqRyusOG
r4GaExoIpqmfwegr8Ek+SjOxWiTdHVG+Ga2nZkkXYNoQf96i0aGXa+Ws4eEp5B0S
C7123Dh+Tcxxn6M62WoKppch4absSEBt9V3u84tQNUsW4IpwjBgW7QdzGezbMY8i
jJKx3togvxTxQcUdwlRneCc1v6JmoXmBNqbKc4lzOs2UqLEnYYgA59H1lR99gL6f
Use8S4bSFOh72C8CzNMhKHbjRjHN0jEs+ySeIw+Trpfh0r22ecynsL//dYYRki4N
MBpNUXqQc2z8ZmonH8+6kn8O5SA39M+iTLpOo3/az8phAuZrwxhhy2dTD+M8Lrvh
xGQNOSHDBH1cul0d0q7AA7mnHnQ3yuEXkxunpYZEYxV+Ca93GJo3abyaeG/U1hqq
kS0m9UhSiZ1hr5Y0q7dbZTI2nOFUDPEebRYWm2e8B1tM5wdxQLmjEn+Zkdjl5qK9
3yCH8LHT/5gn25z6NEeBhB7ZxyVf7u7hlHx5fsM/3GP4kwpt8QSuPwfybAZOtnJc
5t+nfN6hRS8KPu3KBkruB1hWncQOZ0RJfUGGlwF/aHE08gy+/f/YikqJPsZmUBrx
i/PvWfznLUMMsIfnrWXASoA8CBi4iMKd8ahE47r4plwI5pAJNKmaFGtpvnip3uiy
B7vWoMX2C4clnFIMRg3v4Ng8QIAfOZN+l4G4PMVkoMK1AkTXrR33wCILnUx4L7FQ
pmA1g3K1UMHJnsSNTxpqirERGOa7Ka7D85nBvPLneBbtgmxd/2w1pEs7O4gUDWEc
o2hYCFEc4oUSZXLUkSe7tY3YX5QkBkfHUl0Cgqlssp7x7lHk9evvGawpJCGvzZ0V
i1mFISWoF7/PUAVgW6nVD/mPITTPewXaqfl3mV3m/je7qtV8maii4EIGXfFIfQor
wRUo0SawCZRlmm9LTx5zSxE1luGZ940tVjswopz+Ie4gcHk0/elzDDM+Mzor4cVT
ZPsw8ZZDfnfuQc3nGEREd3EcYoA9CUEauQo45q6WKdnbGf+wgj9xa6rHaXQJyIke
Q1ANaSI/Q5jCJmkx/37Xl0t32XqmGkcSiq/gzLCoYvl6U24MwBg6oFtvsS4gdhG4
kiXvzdLLBRAWF/+JGX1g9qaV8CP/tT8k0pmC3rHvj2Egyq3eVqEEOhzWfnZ5V2mt
gtlNYK59/+tW8d4S/NCBDt5il24U5ohXZ27Vg7nsWTZRDGX42qTaj4AoYuURtO68
WUMkFEWdieWM3O4zMJ1p9tdEkRX94pkIdueq17QKFqLHl0OhaCkVGE8a2VuW+QOg
aQ9QrGRvPlXeS3WlyeD0LL8fBpb8T/Ir5erWNNvs3DUnLWQboRuWCKhP3t/AONws
h3RvtgJfIoh+12MBHAWdGfO+PHDHta09JZkQyK6H38mA5aUSVSkyB5DuJPLtVgov
Rskw1e6XxvEGWcsTjg1XaNJipDpkCBeAGRzjSyLINgKPpnmo2mUBnT2dshMPiUGK
mDiRhp+aPjoseyBk8iqGtuwtdAmWzH8EYMy1vw7pxvUI9f2NpV2rAw25tKZ4PbC3
kuteZP48NJtrCmSVYD3d33uevGBwkLSUsrslk47ZUJ44c34XZkmnZAuQ+JjT4K9P
CO2ekVacO8ZlDKBaIFqQONkaBOLhOHk4nZFoEVZ0K4xQ9BPnh0A33xOhZriZIrXt
cD4D9tqzu/AHPZXJ+u3gkGRiDsOScwKxgKoEhYMpphMm4FaJrOwCssCATl74bpIy
0P/5VBX8j2H4koSvTtXnfGBE2JDL4n7t4cUDyrSoJKM0jnfx1LN3fSYALjXy4+Nd
qqurJdYLnpUyu4V4BdHNnQ==
`protect END_PROTECTED

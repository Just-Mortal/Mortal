`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8HKaG9LPPqnUoy9RI92ph46TfMKwN+ySe+VI/pYCTB7McUOvPmq0owIsLAaua5AJ
gKFYF4dUSDMa/ZkePakdSWga8myxJABRLhUXsJ+We6pgoZbe8eBvWAysyNtHoKk+
HdJQq4ZqqXiykbxe3XIwjM+teKe/USTvnTNTZbjgk0RL73uOAeQxdBQHstGxJKXR
gjUk//Z83a2NRrAORIXcVWuuYHWGqiU9QCr3xQHZnV5neSr81CNaG/9t6/Dwwmea
9nrSJ5YRMDPktXPyxVtQO2RVCLT3fCF3ve9QA7LfaWgZZYrV2xEQQTBJz+TrAhGX
P5HYYHd27OoqgCHVz4uzhYu/GoJVuM7JjagDUL2z08/WApzuvD7byQgdHAqhIumk
aXAoS+GxY0WRj+Hz49GaSTi0nF/LxvDixrrj/cTGZ6jddkDxflDRKc9H74e90iol
1W44zNlOTwZtiMF3dHja3hWTTE6YP5pO8DEGN44128Y/3z7Rn8fDnnVnTpiiWFqL
SWCZlxdqzeizTh8gZ4qapBq1Lqh7IKlOw1MwX/byiA5E4GByf0Xj+l2TpKIYiqWF
NbrAjDdt5yd64tT49n17fizjYJ0rFNAkCD1dNeWTVbDcx7pdkiB/ct/RVjHCzwqq
Sr6StZ5Oz3hH5SzMWUAE5TYtQkWnUDLwq+DuBOvvcAUyCnMBoBZlsQN1UTGi7tC+
cZCC7qBQQCY3ETF8jqZzOswgStgB4fIVBD3SFiQ9lhnhkyUYbLOcixm3roFkFSCZ
fFpyMAN3v/lZyxoqARZFWIaUOXjSnDz3Tlo9MDMG05lXKNOj/J7zFTsaoz9H6GMU
QYyF2tfccE3kT+GitsKXBon7Vm5uN0Q69XD/OQQvYkA0wmLd6/kvmlZcbbt/+lFm
G1WrFqGnZwy35Q4bdbF3qh7MYLc1TOZejpE2qY3rzfoVd/Sb6HOljhX2pOEahIgi
Lcu5AfAHJ5ISF8aW8+VfL7IqPCmVvmAYMnbE/zejkLkMqEZqK02AQT+ANTXMvRz+
lUSkIWM1q9hFDpduSuLewNSpIKP/Qf5VPswuWh/Q4S/s1yGZTL5GUxQ98mkXG3pY
pTC6CxlTMedQhylO/4t6SeW28GzH/vd35pJ/tX8OlzMk89ZaEXd0NOqD9GJsa+9z
g6cQ7EsWak2WFPtepdCw/SiyPnQb1n1dnidwgxk8tz4wSvMY+G8Cp4MtYbjpaWDw
CjKMJlBI0RUxSe1V6Cvs11vrXSjEzBls7KETVp4V9CXTTZEXiFeXKKfikHF0vKLx
n0Z26AsgxVNMXcIsn1J2GW8R61WXSeR9NGs9EReI9W8/jvaF+ZxkF/LrKSAoTpEs
kes9YZU44NG+s6fMS4rj7K/R3qybzdbFemq0NJR4skYF9c6eiNtkvzLH2vkBQALF
+3q/7CVGi7//SIL6Dn7D0S70NTL4gLByE47LlaPD+qP82SX2+4GEdteJGZ7adTEK
Pefhdc5BTQLAbNtGmPENKCqjERzVjYkfHzLaYnJMbC8xqiC3uKe04y0MSlGzbq3+
UoSikv1c+3ytB1obOIFvMdVdprX6/JXhoFzM/VucjsA8O+0OXI9ZWlC8oGX26nWG
iQK6pAOYN5Rg+thPIe6qYIUHLRDE13Ap31WifCvtfd6g0hZjzGNerbE4VUockI5w
3s7z7MPr9wsJme0KZoaBZe0rU/jcZW5PE3XpCK1M7zmIP4xBrz2Uke0Px9DIEVZR
oUpjf9Y83mURlVpJJChAdzNVjvolNQ+HfCXvSXVI6lPdvllk0f4v1UtdGIqis7Vg
FXSmn2C+ItRbWzsV/rmnZDLFWkLNLnkd+fPGmbmnp4uKx2hJOcZk0yUQHySXVnxS
H+bqUKTIE9kLOtmqZfwZz//lvJu4TUd3ewq2N+sb1bLSkhxLjH84Gnpj/PA9TsL8
XfOPUiXet3b1ONFiWakJbJsnOd+R38VcsAYrb8QkaWHNIyaTiUiVPQd8Evut051o
rVMVNqFHrla9lbRvobebUfVm8j7SnMd1CIJB+GTZ6PTNBd2fNXwYt3i5f6a2HUr+
r+6L6ZX5mriZSHofra3z4ikFdSR6HJSdvNmg+6koGpamgVKUDS4xv8kGq7OuPz/9
ulm+UKWH0qjR1QUxKZFlZ78DYo+Ylq5FnObRVWARLRqbAqBAwogJkq8/o+kgxV8I
SfkvXgFfjRdM2za36unCeuBj05YtgBeOMutvLehJjI2Qm3+/MICAnNmSgmCQB2yS
0IFhiP39AB/p38Q4pjReIPl+Kxd3D1VWTgSGVWK3+Sm+wn16NOaTfSR75dZck5S0
aGZJ3DIyKAkfLZ6qenWSPtCOOd2WD/Yt1d4NE+HM+NCxP2a4D6i3ZMNzYLx9mCjz
38Dr98tqmjUnKEArz5FkJs1/DjvlSy8WThPdZapQtHRIXqUYzfP5V7vbxsLruB2m
6isVO95MKZKrbhLv6oK3pyrC7WPirKBGSVkUGHBb4lFpi/BF5QJgbKipUMPMq+7a
QsGxUAblBNTQFpu13e1VNzBKVLA6jeUoTbSZWaCjrHim/HIdkerIcv22ABojX9Vb
hfaX3MBjSwPo8mI7ZPyHOeViy79cOmHD+xFOEF1B3GfY+l1qau/96VZaeAHDIpOa
RwCu1nJuxqwM1cZNiK/EpM7PriEShhoIhP5FxF+K+QMQG+W7qMo4pv9lgHj8rI5M
yE4qEUbC9lQPABIw+vftY1gshCM8xkp4CSua9jCK9NB7rxFoJEGksrMDMZVWd1W1
`protect END_PROTECTED

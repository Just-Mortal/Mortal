`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
stOnCdB7gxRU+xq/LK9tCApjbOv8R63vMqkZ8MTVAT+5JbiC05vauBwXcudEr0Lw
5OKnP2P2gAffwM+3/qkFdxN4Y286lCYyFUeYOqTRDxZzSX/xsqsVeIRUBxNm83lw
MBTAaEPJk7RMCjxI7YeoCFQlCFQz72BKdpV6uEpaMFMNMYMySLZZU4GRiv/KXcW+
xzX3rXRQyAwhMaCkIXnLdxoJ9R/l/Fl59y2NNyT4Ij7jBfD2h7Dv9S9EYtQjcpqi
So9fxuYoz6NJQe6rTqtYGGa74hCQUf741zBCarQJUcTkBVzuZtB29nvdhLad85nW
rx/riZrI/ZTVJq3F9Z6v8Sfp8BxVtmv5oXqY5w+YybUNgQMeJcg7/GWGmt5LcHVH
GlOTwVASh63eEu4U2vnXtPWSxUm6QCgbesDsuqUWAfsdbeTxRzoxXn8xPZS0F5d7
zwp2XUpOh/JADBCEWTgxz2XHonspHV6z8dgtUXzWHEcRRnYEIKs0Whbovr9KBG8d
tbxbluMDQ6SeMDbUZV2aXX1qsY4SI/A8g0TW5Xzdo37Gd87A4AovzNd/hYiDi8zi
8z8Wt9zb1I/tdfvfnUoTPMdcZi8/pBqbLzz1sq/uYDpTw54bkVOniaReKKNkKm7O
vzDoxGmj0V+dhjixSwmt3wp4M+k+JBNf0VG/QtD+8aN/B6kxHCpRrya7I0I3UStT
mByY+J2CpRcA6/iz+XjshnRXg53BxaKWo6nu5oG/nRRyzEp9yMt0Vl79gxNceZxa
T0JGa4ZkIToimzfJBPb+tw5bbqLlU5U6yHbwVZF8IfX/liADei9JPeJPhr3GXt5H
`protect END_PROTECTED

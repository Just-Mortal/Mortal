`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zMVPpApPvOWW0Z3I5HUF8pt9sySbkCTySUVQgRZet4uJwO/mhbfTKB49mPsXXJZ1
2o+N6B/QdNfungXrpsVFALjU6lROPuUim2yu+HM+hGIbo1Z9d4dzPmjyOHYx7LEd
SVcJQ6/FvYMmyxAhGibpOt20EihK/v5eZALuq1mTBKkuSl+uuaY7RCmN1yvS8bv2
f8BWyTQLLPFyiQNf6tSrHvll6QFdLH9U8JCzbwyHPOtifsHI2V6EVcUQWpz4PflH
DjokOnSFFfbLYMpa/HO1HdsryEbjA2gt5V/qyd+A2gWImWEG9Peu5wD211qfEtBH
UXbvh59jbkXREPGzInOTeSibIGAvOGKaweKgrzgnoqeN8x7osxyMjG1RxUVXxfE8
FSh9/mCevTCGfwNLAcM09fZM4FWuan+Q4ZPQxsJinrU9ukk53TzrBRHl86PrhKhx
GJVfoUUDX3SMQn3Tgdhxut9ISgKttuFVJDDJF93+SzMGlpyx94Hz5UkrpUkkB4JG
7w9GZ0PcSujKvKnYtzHBOw==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DoekbEs3fc/7p/YChzXEIKQuvbSVGa3TLA1KmaNT4eoQDPB2lfkTJxu6sDSJXSQB
mRRUPFMPTbCkOpcUk6/Qs27SbiP56SxjPkl5k+gx+bIgrO7H8uJkMYdPjvVF/cWz
BQWuFH6fL6XDtpRJfCCJPcSrvluYSyCC7xNXaMQxaLCjjDjx6PWmvYugGbtOzuNl
5hgZftxZu157p9/7rVIV1rjNhRkm11El6IFovZaCZ8iXanqEsiwvK8Gj+b9wyWId
4NwlPKTnPJFp0Jg5hsvrNRhYtct4VgqwicFbDe4NtPty/zLvgR0nYlhLGX/MMsxT
nQN8/jN98qhb2e+RW68pF4NTeGh/oGl3VAQMbV73fodvwHKTHB+azw/RVssCPx1d
wl+9I939B9f7vUkXnSvMXvPw6NPTzWzMjZztw/Oa+TpCgEiL6AlF3ChOsmf04hcL
fk4eSGYeH7U7n71gc1gk0RMbvCB+cpgBAe69caKid6Y/QWIwZsHL4dm2eO1B1KPq
ZPj9OLIsiWYyybusoLq8hf40Yn9K+jcYWBfzdfrs1VHf+EIvcUDPIV184C4G0+Cl
6cNtr0BkZ9Hp/oNs1kfNwI+QzLzszSF3BN0cc3B1NIqfS3Imlv+T/uB97IL065Pp
j1Hg30BlxAB5/e3+Xtkd0KUTK3EEx+8J34/P1Ds18iP0yK2wiG5oMLh0F7aIaa9W
7OenHi4DGIML1Nf2mETabiORpABR/M8T4mXt+NrMCIOpFoweYlWwBTuIdDmfH/jo
J7plMQor5lBw/8ijhKXSo+dnWGD2p+vDWnaGJHsMgHm86syUqKeqJMRcDu7NoCHv
h7bzt5+ABDW+SzymcoiqtWzOo3Q4Ld6y/84jTruPCFnH1Kgp7uD+oQa6hhj0CHDq
kXs7mPbkjuD0UUkx22OegO1uSP3OG5ZT1eEZXnwArWM2xUuPPU+GEsRG7jP4AoHo
UkH6XGzWVLUfkRyrF2L0SIRrdfkr5Dvyh/mu6obCaaDbdkpJpQPomEPnDCc5ycop
Qc7LsS6cb9l851eP1id8+6En38iChKxwNt/Mv3oROOA9RuIgFBhNc4tdFgxOQ4KI
QsWeEBS4RRCoq64GTdwkGIiJ3H575rwA3idAG9OZjaW8LuaGL//8LWk2t47k4+oD
OhNaBgtv7FN1E/Vb/BOPbLJGUWOA8EsGeFtx/ZHw2O9J5ndFYO2Y7iN8CrBky2ew
PBbTt0bES3yvIpDPM0Sh1rKtYNuPiGP6OtITaIGea/nbr8j72HhZndfDVD8eefz9
b4cEQN0dS15NKbfffD7Y46+Rl+bBhzcZ/pwEnzxUHJGAUCSEXj1q6P+SAUAMt0L3
Uv/yrUqeEatXff8JOALmt6WYvTwQr4f8ZzwEqMXsHa/fQzTVyDEqMua763/9Mdff
0FnAoEI9xcuz5N8vFYIcpypM7m8Ey4s2cR6uVFbPekSF9kJld/1cbi5yAnsu1GCy
o0gWWsIWIm/FqUaT95kPT1Oblh67cL0sa8k6ObiqviwV51cxSDmDbN2CWas7kOG1
f3US74NYTFl7Sqp1XSCcsyiivKwh+4dDtj4Q+8nv0xPh8GDGH5t3T6zAke0refdM
HggKhR7qwljWwN8D7ZEkqxrHrR1yfKmCrkqprVRjQzkuTwlXRG03y3DdrSny49at
xBFQrCQXsLght80tpUBxHKsE+R8nnxBXfeg4UwbFbnRtyqcPlJzOZFCX26FsAy+m
kLKH8rKW1SD5in5FnrrqhBoDahychfanzIqD0pnbtQzvDGougqwHT650/4RI2tUv
0mA42L/8+wlKn3+rqbks7fS1EjnU1gaU3lGGVBQ3DliT5DcTHQkMVNY092eYc3ER
HpPillPjI+fmtXkuHTqrdnfMvrFL41VNe7odmjScSFUqg7lkj2ZWGZazCDQvmvmc
OWClXxDWWQryOG64aIcWDs7EV8tF6Ki8uQF5JCKJkDOztTUb6iSjqMTgI+D+cN0G
bcpYvXzpzYEpbVa5g7Y+IQraNkjAdttAU17eA92fkCJ2DnR/rzdCNt9LLxcrsPNC
6OyKkhCoRrgACWOJNaFY1ljlBuSy4B8Q8YipSri4in6i7AYIuH1Xf1gfmban5KI6
dxSCmIrGEQuo11dsG8FJUpe4nDjAOfUK02v8WZBthrMNvP5oaYT+wFJe7mFCpBbo
uufGmjXxS7da2btGBBWT2sIXTL/wPF0fsQ27PpXsNxYLo84kpPUojjZglJayAVal
V51zChceH05d0H7iTo6xYyemhZ6iE6hRNtbkrvQ0Tm6TrJQGv3Ues4YKDPNlVmXU
BP06PBEP7VOtI9Vjfq8k7DbRtwYiagBcb/slcg7673qg1TFWSqdYQCiLTP44qfCF
/4p3tfXL8hnBK/IV+zSjICj4HtomLFCvF9j7USwrIX5wfdheY/dCefZb79RW5JyA
lYk9r4yNcRy9xQL76MAC6uHNAPciorsXIsExEDw6KbAcdk6OH0QpD+bMdIQjGXux
RDhiB56lloJz+Y6LcSp1HqzbFSKcqAR05jXDOwLbdv7WVMbpDra07uspxlncSe6l
k73yWRkBekZtB6o6Y4qZeCviDwAy3nuO6kXuw3W4+nDlfWoY7k/xGwOTqZvVYgPy
fbFL5kB90u9tZ5OuwPC90YykY1ouev+/z1BoXdoShRV1IVFM1LhVJQ09acHxw0si
lGbbNwEW5CdeHTScNCNnTA7nXiRVFN5pT4Ito7UiK4gO0HqrXrL7BGxLXv9tnWx5
zBp3RBX7Jc4xP1BHbjHcqEpb+h2EzxMFJc4M3rx8pE5wUe1Ch0W5yjoDkZPi83cK
9YdO2xp1o3ps6CSpsy3fFCduCRYw+SKBGGgiaQ/zcxbw7Bjp4IonoQeOpbp/l9n5
kUYG8+o8eClBzt6yuEg7s3I35Lj9yjQyf7WdmvfEQUaR0OcpvGR5gA0+2LMkWoT7
73zwpHfjAhvWgczBgivaUnqbOHVC7alocDE7Ob+AVQ+e1lQL8y5OdPrLvFFwNES2
mJvN7vdTfPBELkWpEuprx4yTnOLDppcHcRXH9pgr9oFOpvP5OApZv5BmUe+dsT2w
9ayMQbe8yCOnBU7ErVxFgiR2IIcnqhRNu7F0iB339hxBVlzQvoIo6D4uTceq8pt5
t+vLf1R+NMGeuNtzXHhygvNhEDwS7XThhMOPRGBCUGBjwNEkqpWWRLMRVycRj1fC
wMIE/Z5Anu7vC+chDdIxErcnusD0fXuiaxTev5+c3n9ASDQhzcel0oywjGmBqdE9
H7kbUAdfYaggPdTYvn0EdeaGAhYk6VXiSAVmgA4vnjYlRYgk9YuO8l7PA6X5Ogth
lZgdARRaK85nqJWrVUp82lnkh3BUO9inTEwz5y6aFQM=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8A3O7T3APdZYzQI6Uic8g3xMr5ENqvakxFEDIz+cRIwpivBKUXIRWhvmlu7L57pL
4rWJ+NzOciHVWILLxusGL1vNx9BNuGtiUQS2czj91xLC7ttcKN2Bcukvv0oDzSx8
jhIO933ajAF5SxkRMAGRUYoJwOWJ4BtT4s519tE0byhaKBaZiaH/bexPKYvrrb6C
ZACbA2EUMjeJuCOHQ+I2dvGOP+miihADuY89IGcoDf/12yhD+Mnhf6wZ8NMrmL3U
j9icaxrxge6PZSUFzfkFT8+vP0tWXZNh3pGw58gEuklxmL5P/lLmUFjGYlnLJthi
wOw8IUHwPorNTrf5LyrBdeaAyDJ/Y/RY2eR99AKMmVq95YHkNk5Hx2k2xGRys8V9
eEh4hrHm0nY3XUcn0C0P/VtX1k8JDTVUJ6rtqBmqm25+hrH4TwC2LvR7qLuoWOCi
lTTXXHg+vEGvRItYqzwROnXXPhq3YSXoJa4nocGObuU=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qPi9inNl9BBr42VmafBnjjCOHlYWQfOjhyNVmGSLkhTO8lH+PrtMh9LiTXp+eEGj
c86c+QPjZ+MgaYznzjXBZpyGoyG0wK9mfejqTheBr3O020EKCcqwjS8MbCDfaiE5
jpARzHrmu7XsCwGr2S0hSJJQ779igH/2kN7JprcgLAxMwgvxTBw6nvlI4yZKv6fg
DiayxNtbY48TBiCVi0vwuBafrQ+TuOgIt8tWo5jYvgEVIaZBL2l+rF+dHY++j5nR
tHU5aqJUqujqeuIU2oGm5IDEP/+bDzYV9L1bfULr3nG5jPCKkH+Xkg7IuoQgk/hz
X9odPHsjEnEcbFiFThpdwOYyh/1Dy2pbQhfML7Rtko7qYMZIAXZO/8F/Wive9pEg
/bOOCKIEjrGWcdb/xamf0sQytqsxXtVCCzr8Ug02bcQ/9VVkkL5wIkKOiZipcKCW
azXqXfhaktUcv8vLuSwTotVWuD0CAOH2xA0/mYt9ti48WYogXgWLhFuNPdMiRHK8
ucBIj4ZjEz8jxJBLMlA2vn+cAVsWubkiTDr++9ISN5GC1QFnNtPS76ovEOJECkXU
QIgR0qK1dPUtwXKxnKM2L0q0+BCdnpo5Kjp25HB00LylkyXxMYEINLqEcZLcHHnJ
BQ4rUcF7DwU28f/o1LIrctDIFQicdZ1ra4sRF8QNjgo9V08jVx6pNOzT/t32Tcyf
Ow7WprRFydX8jDsJ6fJTPGA/HF7FBpKxB2EiFXm+aBWhQPLZYZQ987xaE104SkQb
B/mRlu+XuZ9n5/ZM/L7EsjAkZ6O/8IvwjN+AfOZOuMjIyqnbnqxiSi1XzmZE170U
E0I3JSXbyxRkwm2Map90Rdopx5aaxZWmoHgO5H56X3JWN/oYE3zOt3EOc3JgGT9c
qh85foVzGRbclSneKJVM+4mrCcMKpWd7PGKnwqgGRm4Cy283QR+WRrN4x1dA5Ehf
tahx69t93ku5PiDP2sYEbJUM7ob53cvo2fzpl6z0LFkBmLaPkPng76TWu9X7Ntlv
6TWZ6q1tYzHdwVt9pQ0JTZQGfWnfn0aniw7P1vhgWoN6RBJUbhpdbOi9loT3qoSO
1aSYcZE91FbDXaJvFoEDvd6kR+Rp0vLSNtWXmxythcYtW5SU8tRlXIx+6y1GvRTd
ucd+qk4DvjM/mZiK9xOK7nzLPGB9t9E9qodjBaMIECu8h8Wb5XGl60F4EKa22KDh
9uRnFhvpNzNoilQ6LzYI8EMAjLg5d36WZ8Wuh4Wkeu7FD7iMKqP7/Hg6Y7pm8O6K
eBFM/qig/3B79twonfE9KgACxSBoHWt93KhuUjU4D7GKoRN7u8bot7PHsU5bJNUt
O+Z+GZcOWrH4AT1LcYjqp1y7MnMLgmLKb7Dt8I+K4fatMkZug89JWAkfG5cvuuOA
erQbh7DCJFKViL8BhOLZc9lLXKim1iQIyWu/lL7ZGflVYJJL3EpBiJG56j0y961N
k1COT885zKHXC2r84U5nGlvXOPriIzK5GnevN5Wc2u8N50G1p9GIa1Wl8LZy2LIf
6KsUrDqyJLwSbzrGf6LkR8dQp66cV3RwhYqQyCCPSGencTnDFCP2JawM/ozeMjCF
JwYrYJz2njIYLus0QWBhdfV0H1tz/bi9Rnpwn+/GP+TQvar/r3gnhxBf9eEBpbfx
54fSMIpv47So0GYl/VLBsDfImtd03T1U0CfY/LZa8q3NEu4qpfSXrIQsQI7lGkew
Fg9GpdQvTy/uVFP/HdgQ+ItFsIosBcc1qW1e9qdkowAxz6wOEqgXmmJ8AEzgUCsP
AMQaov+z2CxMmK+4y44iNTi4pCNMALYV6+0xKI2AdZ7riMOOt6wziUYb8MyVjmRz
bzJy9Tg98EMLT4e7tcP8dtT9u/fnFI39HjBbdSxO45RBtDOSFF7cWyM5F2XweTTp
f2dwFYcQi0Zr817RDwkOTE8B4VkBjR6T1YzWczqx3oWJzG4mdtxBv5My5uBPnX/0
bGUaeUn3Uak+G7S9LZqxhuHUHHfS1/Pycnf3xEgimPv8aI65FWfoHBvMhdR17EYI
+V1RYR04EgFfolowduDW28JhnLsUEScs1f1ZCwbCpVyz0fdgpHFGLg+ljfGl79sd
yNqOG+J7hNAxsXbu+mWK6nvRn8bQV7KkwlHHqklEiVDROK13o3v3ojumhQqLYffh
DHgszhshfpVqxynicU/47gxJaovdlBrF/Y75WNApbD3y9+iXyKRVIvv28bixclPk
9agldmJ0bEKmT/zGW4PizPlfWx/eHUyssFpmCD8DoOelDIDy+YNDa8uwuzZ3Mo+W
p8JDU6Eu+15p2BOLFbLo7LoZTn1NmNikE2sbHV0MUDQsrLLQzfhmVEZ3pDn1ngFX
+rvKfxvnWy6uYCtblixky33W4bYWvwpq3trpsPBwUswnE9K7Xlt+NaqSsRkwYUMv
auUOpuB8sD58YnO4z6ussSv/CWU/Ty1aMNscRwtPmyhAcipGSN2MCelwJavCi0RH
GntB1VwpqZPkh9HpmoZbnF7uHfMWpkwIoKoKR83wbdKdx9y/uTVjIMvFq1gUxndI
I435sTp9HYtymEqQLELFffHhhGMpvEr1DFj/ssUCujzJvMpPQ6s/csjbDnv/wtFF
863vy/5+pDaQEh3+FMNSyRZPeCnte38ELiZoUNQKcDwEaBQtpzEjW59ehMkS/46f
+YKxIUAavUUoVkr5dWHIXW7gZnmkDMTj4Wk1nBf7295uV6BNGsqYwRhgIzoJX29i
k1Sd6cPzVd39OlQOHnsI+GceZ0MhngoOFyFYlwzktB+OE3lGaH1p5MbHxTXMBMtW
TbgGQSy/j0nc1q1zp9gV8wtgkSyhIuvALu+qlWXai+YrwkCTc9y4OXw5/zQaz88K
0vDWRdK4onn8OUln6GiU432IDF5nsw6yaFtCWTdpkICcpyH+pBBD89nP4GLGrNEa
nPf9aAqup25UkCKQccg9+X+cuQ1HlRrsZhF9CY+R64E=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p9w1BRRp3KGCAc8jbtTgxWVI50+CwGH13swPIsSc7kvBGmQCwk2zpVGhWHm0dWyJ
D5y6bpcMgFupiwdO7uQExxOXzVemcPkYdABExGoU2B85iETiOLgtTN+Kv9vlNcqo
Qch6uD19Yshw5pu3h1lifQDUfe6TwDl9gYRRCSEbpfrQdtHy1KDTvLlLjjf/6nmf
8EvOQb2+jKVxM9eYJ4RkSyVoZV4RJOOhINm3jJrkuUiM49R4WZrmMChmFslZGGkj
5OJ8J8uwulvtXlXb5ySDsi0WcdWH0urwMekiLFaeWImocgbta7xBkZ9RDQwLvgsB
A4F2G/Hz9B/PBLIwexYFose03RL4k8iEktQfBFmltIcyRerkcCB712w1H7kikLbg
BOb6o3cQLCBq6hePz5aBYm8gdIxK46w1HJlgIy2m3q5n2A8RhmCTSyGjPzw6uxGE
NX3EPXyRfHk+ay45mQgs39PqOhsvGK/ix673icaa5Nr0H33pM4hiET2NWd3TOHyw
S0DZmqKyDTYFjq8jnLzaD07Lvndel1dMmdVpnBGpaLte02aPQHRP/QmRrCG0m2Go
rA9Qgh7kOqePoEWpt9Ry8Ek25lolQB5S0vork8J9plE52N7ut2jyOHhxTZtDeFdO
DP6F9aC1F9LyfidAlGDiWQoe/bwHJFOZB9k/mmpC61HjSB6AaoOrFBmiOSxOR8b6
CWKcPsJsyWY2wFXY/yewH1x8VO/l6UjkupRlo67ABEgfzms/jPOGr/fRLmA7b2jC
82/HkxZgzQAjOKzIZxtwMygCYUds2R3ykkAp91D7IZNockma5lxNUzsGCGA4UeAT
SuBM4Vspwq4kGny8GcyOhr9waBpKBTQ+vgdtXtfPTp8rrfLjRLZT2YniZlH20BDH
QsiPLbWRgEltsuWszYzDySkAWhJ7A0cZ1ihkzTa+fjglPNAUd2BgykpEigpfsyxz
7RIrXCQHhDwW8BnW7e1KJGOIICluOKkg2PJ1HWZ1bYtFqsJgMDr6iIZC1zbbG8ow
QK8sUPio32JPZSNQisw+4kHJrtL0JBxizvV2XYYRNA2sp9v3MSiI2/uh2jPomaxw
gWdiTm+FQstV23lpHX1GI3sTJwUBRSd5Gne8UgGfC1gSNgtL+AnvQhB4EJMhm692
xg0WAGl7Km3JkQDkotADrNz6GcpA3nxR4hHkZ0yhMRUFp4HGx29HYICsAvRBBpWA
ISquRQvq+9uZqH7++KVabqCJfnf9Q5Sgf8glKWYOgXE2B1zdvZTy1P/XDIj9ImXY
D7GVoynuS6nkRU3ViyJdElI2G0Sx0OgeafEeSdjLfeFN++9xl6Dm+bXw+K4pidJ1
AITukZaIllDtBXbX/CdUSN3j+tNhfAL3l8v60Wn23YVqVtgs/LPPNHj/kQtd4jj+
54lDiZeQu+25omm8+LoSfrwv8JViR3gAv/jhD1xZ5d/Z7ZzbO+n+y5Cr9djdYWtK
xA8b628bp6IJLQa9kXt1t+a+1jFKznk1zevRrM8GvBwjXdVg1nCz4FTnMlli4LUR
KmJ6SCUrEYBnX80UZsPnZbytqoz7jC0eHypmurhs2Asjz3nH+4rZfSlRtePpdi4l
JouV9CRGes+oPwVrB/PyNc6qU7gX2PD1KggGvdYEUqXpsiCSYfE3wPn32OzPkk6K
bFuWiKii0Duk740Nbp3VS8qSNtjAfjIp4VHXvk4n/Vmv6Aqqt1YWngJgP0zy7Xz7
JVzAULlWNeM1J2kisiwh7YM8PUfF/33DvJxJOztuhE7/z5/jYMYfnaDZacHRD484
E8wmRKl7euzUVUuSaoLchcWE4EpNDjqKu8IgufUUP2HZbyID8durp288IkvpUhGz
8HopK0d7igXbUo69hKGKKoRwf0NGEAmmPhiULqr+rIgA3YlK1qq1IIHWCrQWFGBt
ZxvmV3s0EbqAiQ87yEFKAOgVI0uysQGyoe5yQCIxGLS0QH86J1rwg4ris12dMO4T
J+zbhuAcX9ZnEhNa/IHaZ32b9rYVsmFItQTdRc0kWztD1HvmAjhXEFwHoghsQg61
2In5oNg7faSIFcKG428fT8LkBZ1qR4/AJrN+YKgIwOm957Ts8DZAittbfgaUFxnf
MqJhtEb7o2ejg+ddmu+lGKH04Qt1aGZP+QTwbiaVv9ISoiCudnkLo0DMCYyvZlnj
RlPMVPOfL+b3vRtniqHzKRKAKnqefvNWb6BemLhsm99rFJGhueCWDGUnORKNRFbd
zKsvbiyt36BPdLdMkY7on4qjDnRfL0Dr0i/c5Azf4HLF7YKMm10JLs2O3CEiHG08
t5ncUUuLPqm8xBwsgch6HDKaAvlsC3mQ9JOlpe4JgVxp6ttzr9lFAYMW1WFp2X1w
kz1fACsT3rVtxDC07J3E1C4JuHpocGWdcAGo4mAdSuaoha5UwGOqfb0QH56OPy+Q
areJJRPjs5KXcr3OAz65Qsr6UcbZru7/LKcvXzDROdySDQoMbl0vy54eCYWfUH3t
Eu84Tcy7qa3lO/+xVbtpz8vNZ7SwMgyCsbAkVlSl9ZzVqPQtQZRDTOQm3sRRmVGg
61vVJWig3L/KpQWsRf26z+zlh0rhlx+1x9hnpfBBI+3GSS9+PremtcC41HoM2HdA
fRivDUQgdxC9ogspQ56mIqWSCn+sBF3r8Bm5rn64DHQ1jNFGbc3Cu985cp3Fs8DU
glUHjbPfq+cRViBXVYs56N9nOeljJY8sdAv8sstQPG5zonxQaPh4qt1QAzfhPEeM
FTrnWgJzHa0mzlEpJH/5t5pCbKscRXDxF87HHZMvtIjZ9m0fJOBIB9an5sq9DhKb
bXZVrWcAgnXD5hlAAPzvxJsMsJxNwbGw54DqN9ZPDTjpyPb5o29wxtPOYrMvgpaF
46W9S1P6NYknsVxaCx6DD7HPFCvdrCIUrReStDvAGkYQPvVyfZAGhw928lnz3YH5
OVq31oCOwbnz26BRTGO2ZwpATFva4hJMlc+5CwPXOmMmcYhr9uLtUEDcMQPuGVKz
DRGNl9UMXLm5LDZdPlmoN9CySutRv8xc1yc/rrz40g3Yz2Lus6bOzq5qpebyafQu
GgfJJt+tKw7CO77WJmzZRlvCkAKMvCpK8qxq7QleMYk5GY3XMl1edkYXxPC+THO7
mv0pOkiq2XvwXBMXkvOZDSaj/SjxRHFWaGkiJbGkbzqQLnHQUs6CMJPRbrW+b50a
m7WqQnQ0O2ZIBR5Amz9dlUcohDWcMsZcW2odksQ7HXLsKcqcM9nm/8IZAc7mmkwW
ygTmHya7TTtUn1e23WSJwo5NKvuLG6RmURwRsRxqPjTo4En1iPrLl6NwL5Ix3LrC
oZR7ht8Fb/dsUZz/+WI/iB7Ykrns8pSuHHCsVsuVVjvA1OrgdSDP3XseWvSK6xIk
Qt8iDG/fcX8VG+4zpjQDCYgvabLq/x5/JSazj+JZJPO92PvDP/YVASfzFONgAkBI
lPJYuPL95IKP6sWQQ2AZveVzTzBMUZs1vtMl4UPy3k93V0iMKui1gQaJli1ZW+sl
SKgLfFn1vuH9MYNCL7QwMwQSoc28AcyVzuADzrGsy3b81SMS1bySd86v9FpXbQRx
eZOe29GcvIdacnNwOEs0dQVKJyHLID/SAL90r/b3TR2dvPpVK0ma6YMWjV0MX95+
2KTjnaEbzj9xqsvXFCnknDLQSz0V/WuW7uNSPXh1CkwgNlwYR4d5EGwG+v410FaX
jTwHYvthZSseLQPJLngQLMvG0w1gLsnV82mQepV5De0ZVAOb4mW9Gsf+gMNfYFzr
in0Pz8QZ9ajAwwnrOo7L6kmn97P0Kyydv8/DvnANaIYyQFK+E9UneubKISgvYLJW
Bul4h5DP2JpAv8UHIGQGuhZvKDCuKukvqfWAVhTjvEgDh+mgpc8izyf9b7zeoUS6
kchELqlfiKeGvUNFi15aFRCKvGBLHqkFO7cqqk+lDzM+q74lGdvGmOsMSG06FrGH
VQl2FmoX0KoZoCm4MfM4eIl69nWM3oXeXrMa7FUEdTOj3mpa7w+fSRrtc7uLNTWt
8uaNmhBs9CIMtLmFSmuy7wY1e0sB3wL1cILwMyrUNiUMBRzlBRfqHceIPPvrCtOo
zd5leQMvcxdbcykDPxLHUhGmOTwxJBBtaIIWh6NLdVELme/s7O2UvD/HLIGH2hKB
NnFf3i2cE3f7W46u1U+aTkeICYPAKAlRXfm4yEoHQESU9HuFjQcihJdBwbG27HaM
x8i8RhHvBAT9m3xMPoaQYokunl80gWl08EtU/+yZZJDVpOJqltibT1qHKdX6ZTil
BgkBWIwLmVhh0PIGgv4F/p9+Ks6OVrjumpRMslfVT3xta+Sc4nlerpUdvRkKCagL
B5o9fARdkPkOcVPRO2FhEvlfaeGVCSD8ZOj+vS0HMPI3CU64lJW3xaKImeiZ7iBm
qGS6h+GDgd4xDEP3Ar1LG//4yGhr5nlpdmW68HmzIkqbwCo66NmVPZPGkOvDsQ0W
7JLwVmbH8rb9t8Vc6GFx1x6LYhcmpkwKxPAdy4QCmKRaF7eGVai+AqP1xJIiXe2t
yjTLhQ6ir5WWQ29riG+mBmCXSrNpfVxf5U9LNUls8FmkgQCy/sRF7/MXZ3PsAwEo
lk6y+pVuWJCy5qd3/sltIBqNjwjiXzMJRbmXsUvcyce3WBuPz/lBFgeTKrczBcDf
7AnnowRgMO84ZLXpqLrQMg0nD4BoTAGfU6vMPyfLxAUGIUaE4WYioo+Xh+eOEjkB
sYGmR27QM6QF8o72OACFUrJMhjKjbr50j0mbTBi7Vjd5pUM9loz5dn39PYLqNhjF
FpsGeyg8z923Xbah4e7Jkistg6FJHrA4sFLVxydbovmDqcNdXI7GyYsbYVcDqCbg
6UrJtaSvqm4tW35hEdL3sJPjzE47iCeyxX4m9fm/0aBrqC9uVSYyizUGAbffiEnw
6qyLJ22+WWA/oGYPCjb7iZ21UuXlPDjuezmkcZKynMqwDB1J4gvRbiqmH7YZNWx6
7tqzAk0GAxf5h7O62KWPTqksX1ytBEtW7c7Ej9Qi+jh1xbQSwushq3nu2Far0PkK
oTHnj7nQorIj6wtp/Zczvxovb+fGQwDyKiSQpg/ijOJgdtgym51EyeqdKef6CL5T
r34XEeLEhc3tiXITcd10WCkB2jC5RN4aaO6/EW9bpu55mtIW3+tY+mxPwGIWsbPc
0RYegTxKrP55nAPYIUjzpc9b0JhgEfpEM0ZIDAQF6rb3GcbRrdoXK7mTS0PBzOXr
C4lVa2hSliilm208RY97gdCwl/xZ0XqUPOY5e7onsIBgxkhU/dhqTk8u7r3dTOMc
ElHmTYMUA30z0uCINxffN0YDRuqU5ivdDilJ4d+32T3EzUC8YzPq+awSVo+xQ4wW
r6RhkbV0JDsEFjEvPJCaPK+DahD4cucDk7xXPDevSuz2xdURcnyhuk9KJTw6+fud
hbedzmBlMMSCn8hnK5RCCkTi7vH+91sukTEv+67wyVNlBUBhbz/gPcIiUh7JJg7t
nMNctFtdudEPdcsHuf6R1eTzDqPAi0xvRJNZIi0aM+a/ebVT9tPDus3uQA++Zpmt
rOgx9Oudnqgm0UwGIoIhNpFZM7jLDQDHeOZ/qM6nqw+Tw801ftxeDy0v0yvZzpe2
v8uRqG9wd0Z7LLJ8uYM4LCisfb1rHoUEDsViQFK5YEipHxT/FBr1w/Bp2IOGYT13
hc53urA6d5btwLSjtFMI9Ff6SjvHwJsL8bl0TWyi8iQfBzg0g1fJj4uV0Q8/TSnR
pUizTpNtMn45KezqXThudxaxLZsyHMfmnmalp+Wz/bwSiD6jg4B/Y/4wVXuO4blk
rGjZ5UkiuzNe/j/LhYwivznS1R/zMXJw0ue9XJZwejAv8ni/cMgUz43XxIk9LjFe
Zx60+yPAGtusZQrsa9rzElqNwJw4rPqJE/O7r6F7amwTu/rJvHyUUlxoTRYZZizE
U8zUSL5iYY8KTN2cGurl1k4cehOJTJIdiXd+SQ+gFCIWUzD0b6L7ZgO1atji+CqG
mVkAYFy6jDJ90ZdjkWtTpAAKMh8NgZ9syrTmASCHEjwbAczXtIX27uSLSTaGmHo4
XahwCTL1RkVlWd21IPLZDfNAdGPj0rECmNmqnEL6csKFmcWRvrhl6OEq/r7/dPoH
SyQmO2Z7kp15UBvFtA2xcVGDDR1pDIn7KrBvVf3yTI2z2+aTookcT+TmLprWPHnj
U92NPK3Lzs1fl5YAN8xKCzKVKVpx2pajhdv9vbv9KM1V467F8WwDPbmk6O00gcNe
TijGQnzM3H+oWjSIgkDiNDmPvP+smXFwWr0cOVGWJJ7q0lx2mQAMYBEpy+C8hT3B
kZxPphuXf2ZKLY5T7lMgFPJ/d1ExBMnm5586ybC1CfCPXwRm0yoTKyKDDtqYDOrq
asdkkvSqcQ1zjQRYqvcQyyLUQACH/mcDA46+TRLy0e0Xx6LBfDeltExgaoo4prPm
U+Kv5ywMyljjlKKBvXrbOTBMOdRPp56sdYOpw9xnaJ3/nAsKrVr21ARTVOtS85n5
gfzyPA6YmlvYsSe39EEPhcyhQwDT64BF6ZR978n+FgiWLTkcGDd3oPIu/l1bnPvL
WU9NZcqgrZYjv53jQp60Aqh4ZBz10dIcQC3FYmMq+p5GcG47w8ViHZMNw+AKQpSm
0S+QY5YbMoNYMkOI/J6e7KHSFrDMWLiQpmoUbuI7OomveMWNsgj+3BGwteLrsBBh
bjBT4lsGPccfxV7y+ethGiWp+sNR8uPpNd8tOUoCl++VQ0sP4jnerWPsVCkNHQaX
kADR5RWxKd7A5WfBfox3iUqWeTRg+YlWDad8Jg0MBgSw5HF3Jh+l85Egl9TTeUzZ
GHkFDlmXmFYg/G9TBSBRbUh882e9RFPmiOE9Shf9+7EBn3TODGgKa7b4ado+hccL
q1WQF1Yd+hVUhde4pF+/UFWP9Gmf1JyJn7LqJS2N63sBDzvrpzY+/8fT4rcX+1Se
dovGTvOlOTKDvarwwvvaiLtPA47MhQ8NnpB1EftZG5WtQTLs/AKMjhtm8APzudoo
9wyM3Lqm+UWOcas4kvbikrNo/El4lhTkUwEm5j3i//0MuA6MmCFvvQjheP3/O7mI
67WXtShfLqYI+7yh5qo1FqDYoBPj7lewKERkTNUiU1okRuec4Ei4Joe8CmBcXKk6
K1GcvsZ16rwBKfLIlNveJC4m2tOiCFO/ITe7Qc5u/6nVXx6z+AjVvJwlCUBaKD+n
XQjo3kwe6QXTx3TABmo6AJ35ORVFrAWZp6goVTTF0GGt7x0tB+O6kpTuUQn3K/L2
6XBsrMN0O09paDo22hyJlVA1vFSgsgeeTyPKVvL/eUf00CxH31707FKtkRoyx739
sayoouUfA03RyKDKXUhirVWyg+9CRGN+16zmks07h2M5oTwtEutjYVOCsIy+1Zlo
d9IY5WEhSUYk9TcloCXwKHHi3J/8DHDQR5LoSk/3GtlMl+DnGJ65m7/ZoKVo1wZm
lolUoT0o9/qxMgtMDjDXmalP1cAqU5SgZirdFwA8qvu05yuGnMQNP+KysJDdOdwX
rGPoKS5fmXCQrIsY0x37JATwS/Rz1sW2mdKrnfE1HKQLJu8PfOBeoY63xobnZrhk
O9k1y3tY0aLaVDeX4ftivH+ApIiwtQTu2OD7PLWt74lXFephHJQLVHxRY1RGo/u0
498z/6sMNxqGTLDljgconouDvrIz3VBb2sRARCK/ZOOH/HuFAi7IWxrr+uWTji/r
hCPT+cfBEZsE3F3AZVhix8Ok8eaU7MrBuAabg/do/yDuUTR9mty3IOCrRwJpQnmi
Z8mt7jD+qaTsLU0RBFA4ojhWtFS/wFCbmwKU0AOYGHlOvUl4WPZvBnH7QA/Uiiso
0B3OIZKULZXgDmUq6V0MN+u7CU6OXf+2L75RaeNzMfC7BJa3z3TNJaIGmJ787Czt
r6qDiUF66i915og/atnU6MuxAywOSaj9rrsJsMbGGG9x1VRWm+JOdjfhGoTjUxRv
6bwlMfb6kHkgFnAOlU1z1POc2VUJCgZmScojszz3nZ2pqlh0Qre6B46eqlRzUBeb
sIQAQHKqJspnhj53t2GaYR6sjYSa3Y+geww3DxDv7w082L3tAdbI5Kbwza7i8kZK
Lra6mUhCb5em1DXmMkSNK0qcb8vBqC1p2d33Y9Ftas9SmIgzyhVJIN2rvladdTwx
zA+YW0qyjfKxUBOroAT9RNhujnKnGJ6dfkgviV2rotTHCvcGm+qWocT0FYiGhaxB
uard54YX1K+FXiZloxVrujovkfdZKalUOkNF7S1eyps6O2osahOKrjJ7CdXvh/s+
dsz4rcsvzNBlPWuuH2D1YSzHGrIhwial2nDXFXLnxrZ5WotaMpclAjNSoIZu0DRo
Wq23L80p2DdDmcmKTUc6BMr4QNXZQTB7TUlQToVNyQQ+LbNalki3yhjC8RFBsPtM
e9XTedC0aKtuKTRBXXWk79ufsTTYK4J5K5s7wwWLHJ1hzq8A+FVkhgcklLTZAfRC
01FnHjIP/NBAaN0UXYv8mgqf4D0+Ja7HoehLlLdMMdLVNzrF/RoE63NePoBdgYSm
CR2p5ESlUJbuHqnSjvTBcVZvdn2Q9UqygEeG8BypuzEBSpozw+Wa1pmRdIk1iibC
3G8AgTp7GL0roAZerzrBx+gVwgzaB+5kiQI9fUAwX102DipBJNxwoSbBtNfd5Mvm
1aG2DqINuX6Hhpr28buRcHDkjgcfMf4Jlt+MrEhJQGLhSloMK7I/vKGXvdeg+qF5
QmVvjIsEXcUzQIW9mRkK8xRydtuytRhDasQcHliD2qw+W9OaxFGgWvVK3ePXXubO
NihapBDZ74yk2KVr0r4zlHLFBytblJUqEuX0DWihxPxfXg1ClPz2cEzE2L9lbzz4
eczBb3v6OGN0eC97458qifMTgLZ5xZMIvAhwKHB5l6snxruGaTzB/Qu+lAyEe0f7
YQSTxXKUDBb6huRgULujVGIhJWiiRF45j/k1KG9dRWRRfi1H57QP18SrKgqIIXPx
8RENLzntnq81Ier5+bA6Ag2AXNuck9/seVGIWvI0Kv61dC+a8qWzQkcm59KdPZtD
ZiUItMKTsQCSo3GZN3LYjuBMASGI3XMaMyFoTIz1yD0NJFV7MZhXSUg0YrZeRN77
i6iOfGYVMC85TUbm0HwybI9wJx8/TqTDM74crGzO8A5MVLat5XKEpYje0jzxTx5A
0SG+vD2l8Xm8jzH1WjtToeOunkRq0tBuCGVVyqVGRqKYeVRSLH6UpuSBpreP6Q6Z
sLvznHap4lfa2wnuMMHxt7PBwWPGDGxtSQyJJWiL4xWRaOjpGX5AdeIiZXvc1APP
vcTCHmwcq8a9FxwWu2mJ2F4dAQPA86omjpBVV9aYY9aS4u7/S9qaQNW16vXtwnkY
nAzpklQDaGHfuomgv0hiDpFJzhyOt4lZ8JgpwPUxG1N6qvCGDF12K3iaeE7JCpV1
Hn9dyAlu2hAb2/fHlcwlr28GOGymzuO0A7X+8IxGGq3HEGYj7oF5a5iYmh2NV459
lyb3QmSCEY5eUZFpnTldNI5zeqSsKs9wKtsCfaeKphuzPdo4E01TKvZNQqHl2V1Y
1SnQ5uW1XblJrY/qBYk6to3UiOoBEAQDteGM+e6u/b9jUi3v04eC9ZtHB3UXy3nl
e6M5KaYOwnrVQLMRgHRraBE3oYn6wUFmaZgqfBm4f0fEtE7YriNOpLdyOtrEDGlg
vkkmbljJGrBT6Bwrzq8w0tz5b4QLy8R7fCenP708H7+bX81aic+suzjg5SnJ9URq
kHdR0euKz3urnhV76axYSTm6/iEfRSrYIpoJCBtcnifY+V9UINXMTmKdno2xKCgI
rKRjDFvG8Rt97kyo+db4bZzrr/Dt0vjGez3W0U7jamrRwHTtKk5SL9HHMrL60uLc
dQjKOQSR2wChKB87VlTQMjiGmF5ijklIfJffc7GlX0xDQuUSNmP0ZfyW1gCYpWx1
n9GpJrEHBgI9yHb0kKB/bRznRuQjrjM1mnSJjY+4zUuq4V/+P3emnCs0Sxj0q183
cIHvBXJWlTtyCjiVQWH5LfQStjzc/EueB5TrByK6pWG0pjnPBhVEYn4GZPH9dbaX
XlsgK52Ij2MHBoYG2VBmOr7N1Ms88IESBcICThysposDPbr7r7yL8ZwG5Y4dp896
QvoAjgnmgpaXQy38jQ45+1Ts28Y/J3zJNDd0PaV6EgQvUnMc2giNHbMEMsJ1YvU5
WtDZ2mnObVxqxv3rBLOWsNNEnBMMrsLMRTMg+6lARZ2mIM5J2X65UOHJIt7/GmS5
kNi9PJwwvAmBJusKnvfVVFyo8yR5aaGuJ3RveZfq9hgVIqZV+GEJZjO6/2NvxbTf
TZtqMbcSjK1oCgdOpsRi3SE11+e5Cmjo0pCxkiAThSiMZfcoqxy+PPXLfe2a4szE
IUbaC3xow06SDOcQwwroACgF75gwIK20CnDbFz4g5ZFqnG8rDYleT3mVBOkOr33U
Yg/Eho8johE3j0HNZOgsHb4bwjRQE1pQTeLr37pYgCOnwwgfAcoTkpSKOd1mi3Jx
HBoN1HhLp13/hYz0vXhpEOPbQN8D42wFpRprI16O+KRaVQizu2MTEsRhAfaQKIML
F2wkXVVtw6g1oSNrEdEeCVDlSStUx/exo62sRgeDOQSJ6wTvDcu3zVWflIM1d7pN
IfMV+VYLE0F+ztirq7oVNN3Fhz4bFjski9WA4XSKgJJA4X2qdqfsuJYFLL9A4Z42
Nxqa8Qoh/bDlG5SbtqWC995v3VHxgLhrlTjJwA9bscpBNq2/Z629l2JaX3l+jwMh
jQnbeQjn23IyMob0RCrQU63oQeRLvrmKsvBp9mVekHt4Bwa8FkabdgJF8smrVjDh
Sk0nT+psC+wksVz3LM9L4X2czx8FJ3Z5LJdkuic3lOeT4fmgiS1zz5Qsdwamt9vz
/qZjGRuX8fGEdRoHp6uRT1t3GJ3WJuVQJg830vOMv2f/JllL3KF3H5y3a04mnvXM
+tKmCyhqX2DTD/vJO6UxDL51ghYbZrwQDWAu3mqvOFr8tHJgsPZQvpLKfc5FXu/d
ZSjxojq6/yJQGb6BHTIqw7OC6qYHCRz0c8XSnLCjSUrJZ/YDt7mSNzYhPnfkdsNH
w8tN+EygcH/u315+74NkHy8Y5t7B8lzXGyHGYgQVp7GQItqEN86hD0gQipPe8rNq
IRDyb8iMK6j3ULdL9WPqPOXO3xTxOjIyIcopVKwHP+tNnljbHVm7XyqVi2MecjTF
F/YwQaRkfkvfbjJS6pQJ+hXtY62+/cqksryXbYBIg2gR38wiYAQEjQBTsXqRxMTA
F4WG0CA9Cdp7j2fvIWkRXNaCx6UYVuN9e9U9rJpuVW8U1oM0KTwijQu9CvIXqJp4
sAEASwji27tWobgic/HiytkZL7+Ifxc7Oqqy3EdFaY7VaGum4JWBsvoi8qKVMznS
7j6C+/Ahurbv4zLLEjwWEcPn7cCRhJYrc7YDdvKUTZgIV8c1CAMLqW3RosxPcabq
icwXhsNyNSOBAredC9+JXH1fIW6dKHnZ/alr3PDQL/+IgjorxhO09AZv0ppd3/Tf
jiROhGBMzF+GnTvcCCKavlpInTr65Mm8ViNN8PC+zhWRxxM14B8VtkikCREJ/KDL
xQVuuC3RsQckh17wY1HZVffOJFRs3WoWsaPSVlN1gd1eJxoWF0eKvnaGJ+zxsYEX
NzB2rsSazavthYVDyfbpLt2MzlJFmLLizgAVwcXJgbA/6Hn/ghrSNTwD8UwCBY+j
rd57VLqrg7Oo2sI3qk43ZRUXufLNF1z2BWK3Tg3OZHrl2EQmC4g556PC8mrOeM7w
4U227JENcpdswK6fic1kVcnTxc8qa3W6BGG0XH0Zuj/f6sPeyQrVUdQ96Vd3XWUL
9m3MhuQJ10/3TCfDJ85v7lJCmMGe0sAnmI6NWU66jiUKVZJG1qpEPjzMeqv+XhAT
zStlq0n2Y+DhEGs6MKSpDNOBoM8gElRSpQvvMqSLFxyUAW+GVwqZ/L8bI+33Nsi/
B5wn3OEQSEyvfpdA6OStIH7Pqhg5uE2uEzHizszqvg8ncqe1nN87QcoZDYgrItDn
Nu2d/rNy6zEbjc1bKYCDRtNWaVNdCJUpN3n/LzaJmxNW7kKuF1GC4v7bQ8m5dh47
9sOD5QtYZdC2YJL7+KP62HfADJ6iap7mxXXroQ6Qcnn8N4hGTKXAN4D6+0P+3NCO
XvFnAxllSs4cXElOts7028Zmt/p+82qpUA1c14VXc9ssI1PeEp0SbCoIRSiJ5aD5
Z8miFcvkGZDq00u1hKiuGxNkImBQ0bCCy1FapfoD75/eGeVqmWzV3pfrvJBLXido
BI9dCeoJdC+O9lzRNw0xcmie3s/lubDQF9QsMGv+WSbC6iZq93TP83yAFTxU6U9p
9uwHIbuEVv/aXOPnYfYH200qLqVujI3TwuGy2RYp6hCeuAlsK//gYTPxxiFNYdCf
1/7oxIC4EK7IBJZmkvM8sYnJbRcbAKYlzTj30VimQWBCmy62zrnJcBPViOhdiX6y
dMgL2l6FbaJ9xqG9+MOXFjRj6mq/GBtjICxv/2DFtuTUwr3D/SDnsD4sBaY4We/a
pBizavBWMZn18yRIjtPI4i+aOyJ3buc9lPLld42IT7jHAwqwMDMuvcJ30zEZyS1b
2AHqEzbikw3mTfJ9p1MCBKlhR6p/plphpxPZznDTdgMz+7a23Cm2EhT7ue5qIzbA
d+PZx2RiX4eanf2eNNmcBafuDioIEesvpO2NofW2Uotn9VMhtwqXeoS+rUQdF2dL
JJ5vrQwqJMIkpzlKjYPZnI3RDtKfEqlge2QFuLSWAg0BxODlqCMQwMFf9ti+s5dr
5A+uzl2FX6ka72npDem3jgCaQrGzCki0PtiFX0eCZ2gjKDc0569ZJmPHnlWLDkCJ
MjwCuya2kgrlF8ayR1Zscw7kYekLJq3isbDbYOtf5BKUbwRcT+J9dM3KUbytZZ9h
00S4IZG/z2w6D5LJz0dCSjP1UaYb4vXaVWOSov5eSyjfItHWOdAY8QsgWg8l8hXN
K0rVJj78GUWIrH3zveJkn1TLn+m2Ng3+XkxXoIJeeeTUmaqyHYUQ3z5Iyr1refKw
GyUpjDf3OXNATXs64ujdWSQorcFcQXethlz8yciyBYXnUTojO3aq4SE5aVzX6Mqt
+1LH41RXmWCp2UiI/9a3GGDJX0wXtDatBgOxuYDtQMJPzp8gL3o7nxt74RNtN7Bb
o7e9Q4Z3bMNBqcpkVFA8j/V8YVVE8LGVUjy1CZ5J/YNmZZLfShe1HopsZN5Uzy63
0q95pVhiPsdw349YbNCu1Huf3LaoxEuznPCXTmeHQtmvgndUDMJ0MaqlNdgCdQun
4+qrjcaj6NKFKjvoCydtVrB2PFFhcLRYYOtydGaMgLNyWFhyvXcjmCDyfw5QHopu
WcBzkqYCOhXyV/OD7wA7CF4Av00KuQIO/EtD4Rzk3BJCotbtj5CnEJoseECUS+nc
mYcOHNBM/BW7F2tJ+sMAtETSxruaEhpXfCpQWz06IL0pH0vWfpN9WoEWkbBBDl7f
u+qQR28UvvwHAbFz11CXjpFcWK8MxxxlWlBf+e4+1POvgvSbSz0/wzS1mpTEfEZz
R+YM7qxFGMHkx9KDOdhMcTVEpSRkViMyyD3Ii4k5vlRASX9Nl4UbbzB+NohkBE2m
U+GCtxPSm7QwLmniFt5NOCsMuyu1mjWolNhFszvEhpjvQjKpX1fFlF9nL/ZSyMjz
JuaUgqqifHzZ+PiLP0yatKs37GTJs9CjKJvMh0y0CVo=
`protect END_PROTECTED

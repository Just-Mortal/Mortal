`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nm66gyGCILdZrXKSNUouwpWbOl+M2kGPZ8dMM5o/0k6XqCJGEEaIqAM5d6mx2dIl
twipASi+yi7d4y8zS4TojcGeTl9Rl/i/sUwc/NkKbjvB20dTbc3epJZ/DJMCSlDt
K8/HReecF4Xe/j200+MkIb8YIL2rBBKLzJ+5mY5LRKXK39ngRVeXhktZaB3aoqje
/Z01SzvpaCZj19mWjsqZGw5pw1Znnv70bzaST44QgUDjO/ub5jVdTZiihAtbfOcX
5ICWXhh+JKDZAiyyfrGjg6ynpRqguG6vWHMuRp1kG1/L5untIsU4CTCaU8UBY7Hb
yw0SdkCy1+TZ7haOZo3jeobZfvDeJM5KQ/VHWsJZrmBbj92nHlGle163ZVoBV/Ue
Og8iG9Vev2Kzde+pdRDgP4XHbHu/Hit6ku+GK1jfiQUyX4fmfzLmCRumYqbxySZ6
6VHnEUDpBlNHbT1eiwzaNs9Cmz9gADNjDxTMvXSJ/XXi1qvmRafD/3+cd6flmDeX
9KP7KSALgOHJ7gDNlRSMpjHudyeX2e48KkP8K0nEIOIA33pDqtSAVLH5ADNxa/q1
V4tJ+Ta3XGF4x32j+/7HCFPuo2+048Iz1sNljGi0OjF3fZJuvEmUZbPHqzi38vpY
YyVdetWHle5oVYqocFwDDbHIte6ruhcx9mBzO9qeLPgw9BL0sP91PTN+L8XSOqAm
z3Rd4HE5J7fCopTK6jVt/F8S0laD8NIP7iLgDNzR21GODp7OGbqva/HGd93RwPJQ
amJFZn0RQ9F0wozsrbIM86Xz8fTV9/XPgJj7Y5xRAkzscfox1iKibos2fU+JB7T4
wo0cww4bnMt9GRPOLzurjxmopG/hmQ0rEwOgmICnsfJkSqi8iEr9g3amJx1plqhH
GD9jpCsgYHTICKJCpk2tNcXpB+p3WrGnlCkxjwp3/SF++1/Dd3eSV7insl5OyODG
WUgwTkmqDl/0rGJYSXpkLFVjzlKkgNWMQlekDZVvIRb//gqX9zCZI3VwI1XICT9c
PNfHPaxkup4BzKattcYUdOvCWyfSWxIKaZ/FoeKvrWscvtNazAj5Glj9azzObQM/
Nst8d2my87m6Anxh5fajRIfGCI0wj5O17DAe2HlqeHZrZ61BSEyV+Evr8cVHvIiv
/VSu0WydN1VKlAOdKTA5YQxiW1oKcn9bu+OFmoAdZIOCgb+vWOT8d6z/jnOowaeO
tlWNVSff44jlkdCTHrVYTJoIcGdjTEdhb7RETYZCouZiX9dAGl2z2CQm8x4+n2ib
cfIHdK0ycfVfQbIaTkDO/9CZVmk9dqtzoTxTG/B4zrBWK3DtykRsFgXruehCJRVj
+pfrvX1vBVy8aBhloI8dBF3qDTNQ0YhXQ6N371FCUhDqkGP+ejGlw72M1IcMcAsO
ZzGVmmVa6kFgww1FYLEUYU5HorF0WZgLge2gQl+pAL6m7b23VldXziRgL/pYMZ9f
Gk1dEw60/MuxizZ2Dij20cUTqidgQC00pppAu/HeqR6H8sy+eV89u7jCcTOw6hQq
m7MubZ1kSA5nKLlLQnGzo4MbKeYImM2LiMh6hSh2bGGpsqBBx2L1gg8ablTAd6SP
h74tWstfQXZl9G5h6/7x54z95Gw6o6uLhBpCEYCbqNQYlHxrWGiHaAHW3Ct1a8XI
T/dmIHDR33/kT1I4NERlC/n5HT2n1l8Ppo+3Uqq0a4HDR/35DHU+4rl2lQMXULEa
M0bXEbu2HtMxgG+7rLDpsG04gK2kEKqVRA6AMwOhseeA8kc3ES7bdRncjr284AUB
eCjXU+4EqAhgu/IXXUelQZnAhAKkqjmGlTwxjpadGrL/uc4GcQg5Dv1QrnOUrlAU
NKXXamoHJ4j2zzWSx5q9QhwwVSeauVheTmYMv8gYgYQJQx7OTBEXJXtrxbCyQ/8H
j5iaTuxMmiqynnMgrxZEAhMw3wK9lP0X6aS9A1LWpd9qRcZtVOI4fKupB+r/Us+8
haK0NwO94V7hlmaLeQCbn+0NB+jETgeYuqsE6AYJoIiBac2qNTISFLPEZut3Ucvc
NCeRki+gvsIDtYiOTcHNYG/ha4daaiTbVEO30PbCC2fpA162Q4uof+OVvVLCG+20
A0Gj0EzbP9AhzF/RWAcX7qTyjS+ibn4HctzCx0KbvhxhDMoxbK7fnASHpOOxpzD9
emYt8V18rN7OulchA+35gwUoivwBf55leFliikJ/AR5LPNnXRQGYreiaKmh79sBb
4D04VGSEdIn5z10gNKDYWmljGtoIaUzcoC6QkVYaLbKpTlN337FisPILIzyWLRtf
TVZ6LwHYffgIEr/oNn/oe9Nb4K+P7s/oSOcOVVMJgBzjb86idat3kkuE86CJHA12
zH/m58qua49sY1WN/edt7JwjMmm9WHqxleo9Pko0RpHWMNvsxcUFpqkRFBAF8u2/
/VlbkX1fr3pdjrkb26vQ/YaPLoqRuBvJJeldyznoTNdw4y4sjf5WNwaW2M59riOp
qPVS+dI0H0zgu/kaJTKiwKAM3W5fiFJqDsf3MXblVUC6BWbvbEENQ/q52943nGM7
96r9M3c3don459P/DNVbJZ6hrQQapBYycNcOX++OG6HRuUrU8SOHWJcwi1kpIzdL
phhMqGP6M6IC6ub3ls8QHZM5SvIRvQ1g9XWKA9WfY9vSTrJj2cGEi5Pe7Pc+oWhb
67eYir2gsBlg57hA2cCo8XbnmPJRYOdFOkVMDBlwIFLXr3vHYeoX4Z192u73oS2+
pu+zk8s/hxpGGYTqr1Ke2K2dMLviqyW9HHq7LB9hYIOPvtw/d4v5PNrvUSppDVxd
SKqsBRHvFFZPBXJzRdbr1d4VpjLqUquf9HnMy2SpN1UU2MqxiWSeEy7bkWWAanxC
Puh6TBJathlenTp43mIl46ini6yH5Luba2JoS/dIa7VCN4QHNDVDJKJ3vplb7A0j
qMyftaQDaXEC4fYjtn2styG/2yG8jr2K369JFXmPUjKZohnpugElZCrr8D6SGkn2
C9nYIka+xVbeGdAj7P5mE8ICkKa5D5wzHC01YHCuGPsQ0rZzgDOWgoDQW7V7Pzws
oJZdgPe5sQod74l19PxCLds7Prfl2fLBxIkImGM1OW9+UFRtezBv4y0OUC7N7RUZ
Np50J60oO+DIMAeE8wZWAJeb8AMHOtaPyfjbzeNlTDRyEny4ifactsAOLWeVowEy
5ZXPUNqvRssD0AM3OIG3Fg==
`protect END_PROTECTED

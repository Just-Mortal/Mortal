`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ba4YxUmZy0kpC49ZtVbpjmxz6oyxuLCzp7zU9bqOCg9iwchKgkfDQ/auQPOAQNKp
3SA0DtC9KC09MoyP/dc00Ps2edKCHX8k5yPAHRqJRkEimgucdaGfCp5RqrkbE+kb
zDd1g3iZSwrCiAA4QEO1pAgb8LYKJAeRspPAJ44B3dJeXh5atVBWozT9AEgsOxRE
+ut1u9WbiFWW64Y93leyYUWUzgjWdYMpaz+5CNTMzIftqUyZwce9xD785Y0YFfmr
RcBQJoV0tNVUar1Kzk2NtHPmfjaSVqiYjXIWI6MedbDB0My5ciiEZYE47XTuCsUX
HWgdvYQwMreE3lY8RWLP3JeM49SKLYYKQJUgeCWa5NDqSBtSsQ0iCMjqLXTNLPEj
bTK6MdOfyTnjSKdyg31oQzElvyJ8eWPL2w/wo+cG+IrHO0xdXyR0OU0aUHNC+jDv
QVTBRWcRkKsazHJpV9WN4B5+eKtdAFsuboobRk7mJuumgTnc50kzMw0C2lhmX7lh
sqrJRw2JsOUZwAw/MEw+4Q+fD/8PDxLJTkhHyyWD30qXptGtUmjjNS23AkBttOfE
o75jZs5SRns04lYGIK6aoepdx1dkfi/gv0SShWMzazgniyp8saKXvlCXqdwaIumJ
HPI6ktzDRvAOTuy8ns1qmQ40TBCF7q/IuyfjTvL+c6CW5h3Hb/JLKdOu9ocLjQOu
SxVS4DzHI0ycuRhZYpEyXqbVKSjD8tXCNA7qjifWvRYS+E6yZoF4b67kmt3CxzE5
sq/l1fc43qnHGdTlk4DUIbrECRSqUN+BAUKuz6tiduQg4jDTDBrTV55Gi0eWCLmM
2mr21XRYcvQqDyQ2mBlyDMFfqP5GHCkr/lOqb6zC1uAhwWeczzi9LwU/vfaY6vXp
KKz3ydtLeQ1qx4Z9hzdMRdKapdNOs/Qr/9y6apgrcaGp15GsPyfhA6gdVOygcTBH
5vgwWUT6Jh0h5YZeDNj+p7h9shPG/ZNdp8PBJUJFLhwTkmZMcAqG+WUwrOMAt+it
vLr+zhNcFCFcZE7BhKt466TfleL6zq4lr2DW3QkFXbTmfO+cMj7VpBfSyHAcl47m
5KBEBv5HMDSswFONVDVQCyLDazCPgrHk8x6SfT24jKBoq+YfQfn8L9hQTRLJVLX7
q1EoCzNApYiVUO6qGtuKHa0BT98V4/F77AX1EsjmQmSTXmibw1hq+Je6WgZT97QQ
MvqI6Z9beKIQpd3oKZVyXqOuFMyfBwBoDpE1spoPzgUqbsvdwkeR/SujniWuqfvf
LLJUzP7D/+tW19NdkYVNyyLCX5rS/87xBpSHiyNyUkGWa3Nh/G8DdjqY0xSdXsY2
Sjx5IuizTZ8x+vAqSsI42rflUFxm0pnfBsEwnqWMvM4v5a2I7r0K0Ti5H20jzHsg
r+NjrPYGXl+DFsuXEFdIY9uTGr4vXfCaBUgQ8AgYuMz77YKICevU7ipwNrvcRd2w
TVdwQJvytsr99ABjm/N0547dbXxq3OMbSZt7ACEOqc4uBLhtcaFvdyaD5TOYNcy9
WbBHuQJmV18wf7wuxy3jcoBRY1tLzIQ5mjsV0NYgnM0bbCp2pbrW89UcnhH81tsg
hE7KAy/qDV8X5/AFvv6dg3QGC4ZeUCwe0Hcc3P+tuC2K+qlCvCni4Ef1YoRlOyLx
pu9mv3OGF+HNgPM7QKtxSNteC+IwixdaTLczyPLcn3P/oWH/GxAtpHBLNe0RtjCK
3QXxoY94nYojHsDz2M9KZojPGnNgHtvkPuu9XUY0xMpATvA3OwwKdhbDZr5ELBmD
FY5cDhmuaxuiM7K5h4hvIA0u0giqB9Bn3oLrF74cWwymwpVTPnpbVjTQ55e3HJCT
TFFaEU6C4Pz/IRblj99ybTua/ugOhw20UfKr7/n8DLkLmZHbek/JLu7j4oKnLq7x
0X+83SvIVQJiObZuGPGnEHvMZJ/CihF+Gy75XdHU780WxxVhl3swANHe1i6ell3P
cnR+HjGvkApcfQEr7V11CpNRIpSQ8/6dhPVZ/nSwCKZKysZ0Kx64dUNXkIiIPZ91
99fTN1JFyIR8iWIp9S8OjkE+4L6JFMneufmZE//JLtc7avlzo53sJKYdWW2VUzsF
c7il9dKwCpvD2Y5jGeIkcn658eyUhzpYnJ1kviGjkxkRSMpQQCjQ/+0aDE6hoyR6
odQLiIiQIkPHA3wrHojfTJnQ4Tytske0Cf5Ol2l9xqFSU5XInfpG0Pvj2FtztrNT
e9U296AvktnxXC5n2PqEhxrvDrAHmW9UleNAVeTBihKSyajF4p9/d4A2dM2BODbD
BmRWSZzWY3TnrbZmz2FpGCK+OTjA0P5X7DXQFJn4WbYd2fyl9TWedaQ2NaynngW4
+9soZEkjogs3M9ZSl6xN3fToR980wyllASpulvVsQuyjZ0ehXh7/y/8gJL72Qro4
WUuCeKJKuMxB/bpCNCKxrVQ+ybyKbjesDMdV5Rq9kGyToaSdAjic6q6n9BIgZhJ2
VGp+S85XeICJtrrFdc1gLw0i2i/WbevvXuH59Tp8qWTKcnSxGN3KQ+g7tM4ztPgO
o5xNB4UJp8s+R2HD0SJscT3rKUptaOHuB2S/kGf1vqbNvyyKsLl62TuQ8Cm+CH42
SfPCW3M4WiKIX8GsaXh81B4Dy2PldqPjFi05Mm59o83uvAg+mBFu4KwhLWnWXX24
ai56670jK4LfBGRs1Tttq0AXh1uSEeptael2v5B3LQYm0Pru6CZRFOBN0Gurej30
CyK/oSllWN5v1GorpcdvZE3pbefx8ULm7A/PbqzFT/cZdTlSq1Jq7Yj3yCY0+28o
qGeIbWkGKQf8GlNABMhSpFvTqQLVn67XIcp95l8oHmv1BFxEIV+ECnTs0H6x9UKi
8/Cq1wZ1PRWONHNbp7qh2XVbvEsIIwFA6+BujLrnk1wFSyGtb2yEmAGtPTXgk4h1
PsII7IRtWTNBtYeoZ1isPjuy0xakjGaiRI2ThL3Fd0T8qZs8a7bq1ADiODVp9EfW
nLDYD/Amfs1u4oLXBOCh/penzz9ZHY/REJDpoKFrWnk0Uc7/BeLTEGCoy96U06xp
xW7reqckRPU9/OuwrbPdObOLUskRRUZxfO3FmOiWlgkfDE46dNIDjaHM14q9c6ge
DJU/ao2prVuRbZc8WV3D4NXDR/g9Vjbub+pVwdJTKgq7sdO3/D3uKSBWdr/NKcAl
dwWCANyA5mTaIVGaZET5l200HqsMM+WtlJgZEJgXcx/uYXmYC23cn5ZnCr1rHBdw
aTvRgJBQpVHGH4AqPm6Hn+aZqUe7zTVXfLdLv77X0eDQ/Esxm+Gt8o2hqNfkOoSW
cAkTkHoqQ19M4KO0TPtiXerQQX152/k6mQCF3hi95BsdDbrxtZT4K2DnUvXNyubC
mLJsIlFV4F3gYm+Xe8Hx4CRQeDBtwqA/taE+5rfTmNIfBDWAaYmWd2BqO3I64BT+
VrkMVjIlcDg8R1pW4Klo/C+wgrR+Gu0iXQO7+WeqedibZOoi87VVOk+2zvD+mjGF
`protect END_PROTECTED

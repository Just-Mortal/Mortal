`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+evh9cDWar3r8Bdp8a2NB/ubcP8X/fKX3ct7wVw4N126psUZPwCtUQ+Nuuuul52u
95+pFuv/BOKtE8wuk7xdeDinM3NzAZ3oneywCeGQ6McJ6snyGBTjbuAfcw2YnbQ7
Wk7/H5AnSk9gquHhiDxSybvv2q84L3Gzbww2Xi2LTvYayhT4TwdDfxgnV4HmqK1v
banZy7FtpCTvvRpgEkfKlq/QlN2x9nWazkCU9vZ/6esCpTeye+8ZZfLohv5OKtB8
qqSY7+Qydl0ihLC2HKIfqCDQiWX26XhCphb9aK8sc2TxGVPvlFtBm3xIqOxvSPc1
eEnLTHfFcf9zcg2lmFdjSCm+vvYal1XjjZsA3FZTuCNfKchTNqA/TFTG1VrtRpRf
XCQN1tAlLizvT8vPtToTh6lz9Jxg50ig6HkVzcPBnNMC3V7KyQqh+9yOlb6V6RKL
BmDcbkPmpVaaZLz35aoYjuT7ETvsmjw0EiM6oHiXIPSwgKVhuIzM/r9oKuRoTkaV
cGlDy/GMPLjacQypvBcNo/kSHoBGgECwlrdG+iYkpfUwKQGjQrgT/hqqB5mktMId
IAaPsRT90TQ2FDRNaqAoxgnt0s7Lx02tX0SlDeaP5N8y01hKadxIPnVqr8swLn46
mqGA07GlizumnC4GBOFo8seNtwjg+0H20Ht+ZObVigRnlfYCh7zU2eLB9qW18cHz
iuaMQ5YrUcfu9LmyNjtLCgwDsv7iymLFjddcRp9c/yFpOy/5sRx4OZKdzD/WryDe
wldE/yUMvctHSHYezplHtSFxwci1E7Fj5IHIbCLd6dRFh95Jk8CmIbgNKA5soz7D
zykfQd/TYL8aWC79dKCgrsSnwb1tRGsHy/9kPviqBkJtD8WbFN4/46Tgiy+t/1tI
/BV+6wBGe8SHRjxBPNBDZqL1z4i+o4LJgVO+HTKKY9cpzQwKFwgWWPsh1U7yeMwO
N4US7FQx672SasBgoBWKW6CT2vpPxHc5cxZxdUuPU73c0OuUVjO6zW9WDRSOJ0bs
/HUGy6OyqoW55RecfMCZNufyDxjKx3ER4bWkkG6Oyo5RKoapR8pWRi5fL8/EMXFm
yzAFgaYUl7Bdc9+c3Ef1IqOPblYagEhOdreTMNnIRyB3VzS9NwMdG+VE1gOPujpE
PfvMCNNpJj5ophPhSRqXbTJsCJXTVoFyLLJ0P2eZO++pRgcIVVxP5j43UC/TulJ6
IgZiotsR8AiibvnbdK6AfbxPY+en5p3ugcE6Z5ElnekCPy7/r5EGShqoTV7Nb9qn
cjio0ek3BebWHkGpG3u3DGGG6DhlCuZapWbtBh3RMk3S7q1Zdb8aN01xmh59o5ML
Nxtaa/uGMYNlfJFiGCHYOx9GXQ2nCTRU8ckja+r98qNNmB90QdEzbhOrA/ne1fVW
uP0q5Mdu/PMmWzjao8VTy+G4687EgI+CKnWj74j4iuOEdYvJVeKxTV68gYBG2SmO
XEw51sKK6OVhGsutyXwMQd4WZDfIua19raEY2Kl6yxHw8pKBzFwNJ3b3ttARzCyU
aUxdPmWmfJ59D91IEoC1RNuJIXak93mYtBAouaNErJSb19yKjWmL2p/8TVwgL7dO
oFJh3l+YAHTy9rxw2PYhbXAqrQ84xSDf6sl19GO/QGOYY7NIs6Xp5ZSC4gMeh484
zXModw2VlGLWFpVTjYiiqyFwo7FW5JEteX6uc5ExKTKTFBWDLY9B6MKjOmD/rGOz
Q/Mi1pIwISFcOMNrX802RE/MkxWJJ0PsbVo43Cg9XBQSDJKRt5VKSOpC4DfB8QrB
z2UnPrv4NU+9nUaXxGztxl1jGh/53/p2guTRk7sj0Dxhi/QY9CcRNWUwfycNt7FH
+6UclgQheebGh3NvWD+UCq0l1rpAYy+j8z5XdwPNPKkd0SwmFkbaxteyGKKMMBHR
JY5IXtckoJd72FYOxBLI86Vbb0oqfJ51lfxFdHkv81OjycSvU0ToINrSsTKSaNnv
ptE803F2bGY0HKemOdP/yMT8nTES7idP0NWJs5IIibVBjmpVo1rU+tqcZDA4tqa6
OX7aZ1ib1YuSRjiJjxyW5xKejDef2v+GhY7Ia5eanZ2PaO6FkaVHA2Dm3leyfKwg
VKpTH9iIVxfsM1U3wpe5v7TiBcch4/S7lJh4Y06pwJwsF/d2Z1Oo4Pvhc6EKmQSw
aJzFhRAKCnnxpwaWL5slkjIzEagLFDkC9p9J8FlR3Jo4phifyTxJCbsyu4ViWZhJ
sQq5tDBTP9YoQOt5+HxoPMSTGP54FhEippwzRwwbVta3ZIPFotomhFQm3i586bqh
iaTp+UwBTCtgom5xrKmSPBbvDRI1CVD98I/fqgZQDCvwamr6UkHV3MV7vO7OhCv9
qyRrYyUGrH/2+LBML/fmPeBTWO0FcK90UcjBnuDG9bxh+U0SzALU350+8aij1t7E
njVkebOsDXot1SA2GkKsPshfZj7oSNtO9idhejMdG3wWA+1bb5bwiCJYHD15mlu8
W/psyO5gz1Yx7A0FHgCYGwW2WbYky2rxax3RR+IS3eVmkwGtcgvKRKXtzLcNuZcp
+IbsavZsihMHWqNmONOcpNPJlPctFJERF7zriAmaVJwNH8KrIOGS8nhFNVxuZmjW
v50QjaXR1rFeUAidMk+KZ6cEGVe0JccnW5j8Q7+ir3Pavy4E2u5O+4lveI2C30D6
ThpicZ4w/ZdG0WT3otxQF6uTGct9t6moBv8/TuyU3btfEtO2D77y2m9y++bPhF6Y
QA8uzERFF1sjpm6FDq3SxsJwmLvrEdnwLfb1t18K0uHmzDLWknwfiTVJ8AkhDM62
Q6h1ErPoUuSv/Vd/ppVTmmhR62pDv6tA07HZcmGhG/E1Tsxy79uuCEkClCvBXf/M
CUVKUFIBefuFVS3BJBoynHlzYsWPHt0vN1UrTSEORyjtDxmjtQiFLJgy0A0oB0SD
Yu+Au+HG+lfJy4gn0BXKXzxXYmoj6erT1qDO0nshEiQnRVdCZpgnDSUzNoU4EiEM
`protect END_PROTECTED

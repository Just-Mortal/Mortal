`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSV8ZmSOTs6Ha/7QV7D1XCg4fsiWSjbAwWMHEfgElDjICzXNkoOl2K95t/IDC3cP
QLbSdjZuRRcXts1q3DbCBrze3cT+2ZIq3qBbmn2qhqHOzaNMaj/P1B+YPkvwf0uc
FoqOhr4lGdlf4dCKAYIWeJPa1aYDZWZlYHHMTymjDHowwSN5h8gaq1nm/FiQM5js
hOvVz94uHNR32/Gv0RTxuHonvV5lzPGnFaPgblHx5+9XZDOFIVzmqg3opDWQ0GOr
ACB+WtPtPHmuKGbSJFeLlXm2iBCsIXZe0mJP7yDUiu2VlqKTtxCosUPzepm+vctZ
SKlfF7gbNqPSXN6uy1ydn/48RmYDxJoTtu3Z8BSauw3+yfZlseUZTFJLCyrsCMJt
XXetHZplZ3kjZ3QB6TF64FY1VIYrafLSuHI1x37AuBejiUGS4KJeAemkIc1+b6c2
RAeNYepKzTiHycx/295mpAiDPmruLwZG+dO6fKY/zjbLCj3vvHQCxFc3B7YkWKYt
XnrenxLlzI/fAsi65jb246fOn7ZlzAqhWYNf9f2bE4S2PmvgutRYmuwZpaH23J5N
KkJZ1fKZ9MdztawXPWf7LR2UhLl3HFBUIr8A+kb5wdTELxvdVtEHEy5Om57/KEXH
pa3vR8knezen6coJuGMusptNJB7v5pBc3h3KTUfl4Ad+uO9MXIWKTbp3mZZaJbgL
yjxYz0++dDKz3V7TkBAG03LPU9y1nlnDGhlyFYGgZvstIDcCQcBSFo522O570Tzg
8oPR1phjBotNuovWq77JkO1+Hix9PwHpvmGO5h5urQwftZFVOCYAx1EaFYaW9KmC
NDOu7vv+8snzHhXnumA6hcpHeWEEM8WizQBPfCEntajgE9vAqHrlxGStTN3bKPZP
nw6Qb1HExBHE6FHdFaO1sOfVaaqs1Q7YokTyCOp5Cj35xsYAwnhaHBbdTxL7/ZIV
bVeEHL6vlQ30uOUijUTcTyHAbHyIcOUFYDyDdMVKghekYTFkyLb1L4FzuZJNZ6Sq
mgFyvV4oJxpyZSxhH9hhw/0UbgKJTSTy521STKkoPiIqOBB45Wtyb3nGG6tn0oXk
vekp/F3JEACb+FlyvfbGHg==
`protect END_PROTECTED

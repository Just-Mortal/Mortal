`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UDbxnxZxF/4ByMfQtrQmNuA44nwHvmBj07t7Pe7muLvvm1+rZvQ7LhMxMyusX7ah
vPmpQffhs/Fp+cV28l1GHXbSfOTXreQhAjG78wmnik3NE1nyuaj8rOB9//1Y3IXt
C+RZHQRDnvpNNpgKPCDCHaWU0lazv7b79Ub7QU3gBquEOq3mypDMp4Ka74ixj5H5
EwrEVvSScW+UGWENPvPMNXdFng2cR2BvtYw2Xd2z9KtXbkLUxVzru4A3PRheybMs
43Q7+emduMIyZnaAhJH/hOe7z1DZJBvQY+e1k3xFxokt540IIGBeLX1Su5d9e7dt
BoW6GTLUw5RZ6DkWnn1GfEqk+2MBmJjocJaEkhsjJiuBV9dvWAaV8o3N73hxUvZA
8w7aRRzdi8mFSB4UxOhepz7CdsrHuH7v/VA2oBrDsXr9c2E9L5/+KtHM/icepCt/
TCGeBg0BruNcFSP9xOoXY15nwwnOUnLYyjD973B22digjIzSMjInVRHaI3IPV/SW
REngMZKd9wPQw1IlTiJeJAgGpbNAHjQeu3jzOM7xNkaYlInjBSeVV5aiFj73FreC
zBUDqkqdfRUqinLiiDpKVQ==
`protect END_PROTECTED

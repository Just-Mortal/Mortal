`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aI8l17zgWZPDToTyB9/NzHE3QUl3+bbYGtlFIYpuKvdlYTppvhJ9K//5JAilTIkZ
Wd4SloBDJudUzOQyPMQwSoKQtaFeYBoUsZjMHPf0LWR+8Rzf2uwVdq4HvKzC9tTw
+xK26YYnhGsFSWVASpEZt7p79K2d844nsEara4JvH7e0QQcuhTGdSMzj3MV1KJhi
6jbVoSMdvkFXoUetVVdVzTNpojjWq4TRm+z5PTtOuLwW/ohT5QzYsPkdnSiz3/4J
tWmbWF2bG4pqcAgrwiMj/dIAP9j5RIJk1NXvVLKQxuquFRndsvgDNnccA6h88TgU
Q3N54SLxgfi/KJT5/SeS6dA7byk7L7MIwiWL4Pg1Y6eRWwX4Ec5xmkD3JDvrl9gH
AjKSAuJy/TZIk9LiD3LHcSYlunTRWGXYy8EDxBzI4TLBOc2ftLSrpRL/5GxKUvHA
LdTpGcxQtBjzei/V+ovbAJH1M9dqi2Gpe/6z2v6C1VzO4m3/H1Y77vo4j5aILAO1
pVbe3PuMAOXe/NpA5W7FgIAAnCf9WViVJfVai5yghACEuPdDq2NQ/Op7OTCSSHGo
PKHGTzwWtG7wc17nVgqi1RTj448tW52BFwebDieeMvLdMmBw3YidWqsWMpUS0DLM
Sw18n0j7YxtU+ZZKnwuZvMZTczPEGF8JAjia6XDv+wsSa0MdsH0QzV+UivGz9A6j
ommXVI+x0gSkqRXKRl6K9pkXVE6lmVzCzFYidVzAc17e4f021Jmt4cZX8g/Mv1QY
pmrD5I3c4rPgJw0f630M9g83mRJlQsB+U0m1D8R/U1XKhtAM8TWBsjLWp6Fb/PtS
dtVV4gt4bh/f9wI7e2XnCfF2o56HQeXQ/kWZaUlZjs2/PIgCYr6nuQh4YYsP0KD4
aDK2XCkR+nJnQQGY/IaGYsQs/OKnftt0zAl9Ws26MCVFE2CRYPuy7m9vlXlgM7ts
c6iW2WAtSjxoJVnPeCkTjD0u8C6Ze/sfFuKx/vkpiV3lH11fW0YstvlAgCw/Cd36
XpGnGlutrDYD6XcJb8dVWz98TyrEBNIJ+KdpKypxuimmjRIeuHZ0EdVokLZES0hz
qIdFqLgVm3aa4grJgc42Os6ht/KdcnoMOZt/VQZvDsH+q/FEeigPpoZiUCLnD0Gh
o6aE6rFJTbgP+CkghJPNUOaKqjgBoTZcsRbqSQVB/9n2j+TepIUI2ZMDUaBgU/bi
LjPqLdkYQaY6AGU8c5cOY7dGZY5iOsaE6U2wb0ne/vPQsLObvpxuuXkSAl68k2LA
8uu/B5FLcOgtgq5lHeYAQPTxbpN/7NwBNN37pONQLGiO+Esz4/LVqwnX/C1xuRwH
KP5n4v5ZwKENZocxk6VUmU3tibIog12F0+KT0tbLLMTixelWwgTqRoTsnOg4NHVQ
aVzvGO48JzSnRpKYuTGK8i2SeUfN+TUr8RtU6m9Zvk7P8rI21bnFNjytgmIiHarJ
6tvDJhLYuDO475POmkGWi+HplkFotFAqMUw1uw85FNIF5HtQ8FKbUozJqWWTTMxc
RbNYIOdlvdAalJehwRAe3GT6bkxbfG+3z34dVPEc3AC/954idQI18s1NROpBhqaA
SxahnPnPzOCqnH0KLX7ZTD3jNZJ6a+FgvYcG/DLR0H+HOHNXWaDf5E4EMIiDPm/7
ZSUtzKvwAtnScfVGUmqopy6PBuT/oW26npBL8QSAtrbrFtaPrnLw0RUKSwKH/3YA
n11ZO8yqWVkqNMUaUMQJaAwsAIAinPoHitJ/BtW2x5zi/32BNYPqjB0Y6zgjPHei
u0lmb17htLBkOPJN0vA2oc+FZ7ezqX3GNM665FBYpMbqhKTwZu2W7GKtLdwzNT2R
gTqAvgzyuTgXLDdUAigDspCl5vNShoZyzuBpezlJglkuj6Exilpo1eYQyRPJ6Mf7
PEdjdgohfd3MUlGMc4Az7TU3CgW0NIbIkCrxejuTqCXa95pUi7W/hqetSkvNLgum
76HzTxQzXslZX1VaQ0rlislWZRUUO7qfzoZ+Ski5SebTLJFG5AyGZTe4pYQRJveR
yFiOjxAwasUwrK/U+uJ1+61zKB05eIdYTOrzl0MxK1h++jOP6k2hev1pypZeFBhL
LMXZIfggh3QPOUtzd4ImqTuWI4Aj64iOzqCCPUjeE4PC9JzN6euMzwRp4EAowEnN
agkASN+Bp83nXeUqJZ4AzagdkwCjuZAQdtUEc/ktsVv3rCPPdW0DG8f1i6uAV5mq
gd09pmwJY8SAkM8TMicGKu3z8T8KAdIL+6JGDX54Mgc9eaoLVbuSEeN2mePjzalO
tc+e2woHwoMUD6N50hGULdUAuMXE/UdC3O2lwQOaG1IKODdnZu7nD0k/prSWY55L
2xsyC60Bnogkz6VlVAeJEvADyjgT5XxpJUwwXxE2JG6G71lpXylG6+vR5QUrzAxX
JxCrVmwoZXQsj0GR0FYJZTn0WXhKsTkO6ODEsn2icCjyQteS3dgv5IyNiyE32cCd
A1gM6FazA/yrZOBiLZREmFxl8jOtA0UpJU3JFVTOL0m2HBN/Yqo0Ad6mNzNrZzK6
QCrC21L5PyA0/wmO1LBEd3SSKfBetPq5PPQzBXhtCUMukE+F5diD1140x0l6qBPT
y5JNxufn2jR/lWMGC5iyCkkgZulpBCqghbw3mQIsvgEKQBeS0Ul2NGp6mSnuSQEK
8IP7hJXAqpYff4G197GWG1gxVfUpEgQ3GEVqSWPYsfga4r2uSzwqyCtWURazxCLZ
FbGDeQ+rbjq4Web/b+Ow739EnbN848YvhwtXX+1m6X3N+qSPTZExFsJZ62Q5+D+o
hTU127OMlSXCxBKrvE35F5wyC18xIn46Y9cxREnd3+q8xU58+AhOp1iwbSSjjCCk
8EUUfdXkr2L+3SXeZh45/IZquz3zrgGODARyjupfG1H3YvfuKHFDdLZQb9OgUF6x
aGLMG7eFrqFyNHbxH569BtTmNNX7UKYim725v6XtnVrJpzcZbDdkdR7qHy9KTkX5
iwyH87RXpenJiUvPunu4LKYNuuyE24V8EtRhnZ4K/YdZpC9xccQP8pOxjwyCZ035
2xTuelo6M8pz6zjRTxdBHtAO+t56uVAlg1Iaqpzcr9K8PdCbCa07Lp/YvTgNztEX
R23m4xS/DnLLREzEJirYfzonDeQNucpEeHZzKldl2NDRi2PiKZmOlqhJWvydX7Yf
bElUcGwAx7jGHKheTc7IdWN1e4uXpiWIF5b2lYNRzl5nm73NfMngDvMVERZANaji
V01WlP53w0zj7Ze/XeFQtgGPSmdRzMg0A8j60bUa2v4TPQQeITgBXn7mCdqJ5UIw
VRWsoTVEGgJVJsTsudLpE/z7WejewzhYDBd/mToBs+d0JHF72ncrQezPcGAZDH3E
QQwf4yjFUiTkBrXvLGOf+76F9EIpQTvTe9UH35/Cvv18EkYJC+jeFxBSMAJVDXOD
z9pxbXytreEfqp744XIOM71j71YCoj62xNTgRKJ8wftxZC/EdNcAFzYGQJk1Lyg3
oJaunYvconwE4IC8rTVytjD8HCXMgGFAYdGVi+KzXCIbjBOfjPp9rJO4oXPD/mEb
OJbqNH3aAqEVV0Gr86i9drTUF3HlYAdUtBapfYuGXZ6X5FIgHr7MnZX7rsQKffRH
Odp6vdUijznznFi0XdbJi0JE/7JrvR/odMg2mAMGg9dKUwmm8bRHiM0PPWg6M5ff
9olbtLNiiHl996pMTo6N5enmNdJsxDY5+b4bIAaSwi4FR0GGnai7es0xxqEqajfP
YjGIyl6MdGieR84tuWPk5q4Nv4Je9Ch1cm6QnRvcFKhq7gJeVeAoz42wCRutF1rY
su4obbSjvJuez+VBDfJgoBmTEJNsp1OP2yNiD6XaN80HQEW0JTyT1Srx0BaWEvJN
oB4oox0YEu8uENlVDcVNv3H1vTHmi10DaIp2FlbUnzOx6Gl4IrdKRdJvjOSCXUNy
Bp1R++oPrGfn2jZEANUGXpFAK52IHu636+OyrR77fgo2carAS7bvQaamjoXXJdk5
VPMtqggJ5ByJPFSmugxpdXoPepvuob6UUZ0TJDvYuUz1X5OacrCM/FZggI40Xw3o
Y1lJJ9BrL/YyNNwsY+abV5kwoLC6CcmXf54QlfTCUFSCVlWNg6v8HY/7YXVKns3U
EilNP7M6F/nyL1l+zcr7MquBt0VTQ3AzVH6Oh+dTQFoqxTwqM0QnAJEEOoIWBz3c
Olgu/wOPMSBzucrFI9vc+9RjQ+gfOp54vq4zYKa+nRiixBaRWqYVXkQy9uCQPrk1
tS+phx5auB6nmPRh2zv6rxNgCJy8webJIgJGDR7G81U7cFNAjDoyP2wVcyGip2iF
GPT/D8w+F8VUKe1uWbspfqGSi1QvG1p3EEaXfWiUERPdZdUZ8VCrz+cvOdq5hZr6
fL19PXZC5YxDIyWSjsEK7yKaVIHvvrkJGHiMu7ZPqkEPgu4sGCMj+lydjGlp01Jb
h+u4EUftuljMLQRYG3ZUfrxfyq/GlA63i0lZVoyJII68MA6ncx//xTlYujBk5sQz
K5Oul7S854v7VzG3K4Dp0g1qJOTAiQL1YyKTXg75GIFLxCDp/ovQcjt2POI/T4Ex
NKzzpk3P1bJEuiTTaALqEQ==
`protect END_PROTECTED

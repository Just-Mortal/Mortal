`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rph2TUKhEdXCR81CtzqIUq6TzidcBr92/Z5Ne8NV0X5WW/IXVLVVsNr2dYDn41N4
89cLT+IwgP1LULJS/IqqH5POc3RRhAUeLCgaQFYMzhEr7sSxClLn2r4PDYtlkQmS
ZwAwJcElkgiqa2EfxP4EnFzNBfxKteW5lgyCbOUiRIuFG1ZchThXIs4zG4LPv6wA
QJr5lTq7Lh9dSiqTgu1G9XUIE/KY9eybzq3lcnlKmx+/u2fFE40jpZ2Bohf7ukoP
Bamif6SFHLOlc5OuYQF8xoIl32j+evF+W0JJkfcfRCg4sQ/nWia2+qdBBhoW79NU
80tq1vHFqoZg2wyUgSsSlbXl1m6Vh6807+RijtJBZVsT/M9+TfbvHio7I3MUwuDw
V9sCQCCz/lKc8xQCx0w3kptseTZsY7sqIbF3BgRxOKvMfMY8M75+vnDzofL1ZkxN
XSIv/0rvnYde3pqrHg7JKO+t3jSlVE025/3jJSLrM2fkHTIWbhnP90aElyHdmnfj
q82HaDL4q73ogN4Q9kuSEXFfXNboQeE25ApL8XyBnhnGy/Tdvgcxiz2q2qUFrlRq
dnNijmLD4UhHO8+eQ/wYirtL1hdN6aRetrmAch2+IscPv0XUMOKxk9VTtWIg25oP
wHiEfDJxC1OtDZK342dgTdiFVu0gr5/nuf3RA1vsjw4oYuTcpYLnmiMJzI7GL31E
Jia5z/QbzHUOP+Ylr6mRGQoJcVnTDtjQ9DCHUvp2DKHgD1RfdhQjz+2InGhBfGUq
qZfv7kGLrVDugIwhXFtM1v6xpKUx01fjWGS84hGjDRcHqn1vJBz3T7WUtNwksZLP
AMYuaNNhVpsNPGnbGe1uDLTZpJ5BL+izTioaqeb9GcbF5KAIoYSacF6TVxVm7jDo
hEzkRg9NAwinYAmdo3dQY6q7PaXvuep2LippERE8ecazdEVj3W8K/4G/sl2WNKnb
340Z65Cq9t0fdWNQPCo9tfjD5v4sCVt+3jiEcwbuhPGcW8PwrDLs3N4w2KjTnYrz
kraN40ii+5ne3vMx6nx7zxMfH5/N4St6yAAwmqKXqJd8qataPSukt2lhXbEAtbXG
ql1FUFNt2ueQ1li4bFNEHsvPth/NytY0LF9GcTQzrPCQc9tf5l4MhRXb0gKpGUeo
IZMTw2IhQnwUVQzk/ivq0wv8X44bTYRK15lPbpLgZSie4krTQ88Wjow2UYU9+uNy
k2u12cV56nI2W+644MlL1bXEM7ujyy6F2pPb+gsNPxzaTv244LPxOjmjGmgXgKbt
`protect END_PROTECTED

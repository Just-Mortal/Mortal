`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uhBCtgssAGv+tu5fiqJzpfRbzGdmjFxqpYd+zdHiBFim+4uP1jC0B9sRs/W4Ujmm
2h11manipr/Khyp5tCjMG86FIJ3OckYI8MD41uhVIedCBFUjBVzw9ataTFTWC4ud
CQdbPzVTsuq/MFezAkoEwD7NDgnndCKUFBot5Ypkg3cj4GziKtDq8wh4zi7i+LQp
MCAMpVWhfPZZJFNDXo/ZpW701jUPw0o58oe2AZ6yhpIsd7x6JpwPLMCy7gxiXL0g
AZ3CPtLYDV6ki/5gGJL/aVM9z7FLnJDTd9vkInCrwHOayrUH6b1ekfvQYuEZaBY3
nE5Ea2OGdnEBga5SQPGfAuUQWpq1xRAfryq0Ak35JY54ZHIIQenyRAymQaM7gU1V
74/6wIyKmj4Cdtzkx0Zm9uSsXkGdV81aM0GE2SMQO80/AqdFeU5T+v6hnxj9d7GG
YgeBzJiDPwY8a6M/CpWJD80qhy1URuL7OKcT3VjFO/ULxiE0EFEt9lMheaPMJgsB
Fn/4IsKdPQkuvfkNSJLa5AdXfbEQmuQy8Ef0qRH/J+LKUtXRJgoXPP2KzViEcpJl
OzFiAQIqjI8I4vd64L7hpyLyRp+MPZBpdyySrKvL4vM4aRiASOqFoTBR3/hMwEaX
cpr0/6AnXo6Dg0gb1YHh64M4dn6XwltVzHCIXekWbhHpxuoraTy2DVTD2GSpcWoO
VmlOJhjwjvTdYy9Pw5ZBQ2LMhRxRsoHCiyClLUC9h7L+1nTj0hqVMsmlR11TsROW
IAYS9pDMRSgDwSstECGY5d9F6EbC/Ltw2RD8RTy+tIPZ1x83Z8ww75W+gTpBaYN+
1BkqEihTSSrC0e2IxSUuDecAZ3rlzKa0GgP12Fnon9sgbmolVGzcFpbmMKZpYwID
1eHCbt+EdKthNqnEOeKu5auOg+Tx84fCZE0mLEyilV6U4xXseq+eLqGKAFfTGKtl
29sL2jTIUdA+jgu4uwE3Ug==
`protect END_PROTECTED

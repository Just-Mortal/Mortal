`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99sqewFaPzv51FX5guW1UXL3RPYLq2oPbs+Kj8z/aN+upNNsBU/enscttYfeitpL
HHl9ovbuAdExjKNZDi9NEw8uqN7KYYDDAgNwlL5upXyD+H3/AljbJevfzxNdr5wP
O8jVSOFUHmp3JWKPPdlxn7i64/h6t/7fAbgGx86PPsSDB7rp2a9bcDiRoQIUod5Z
7ojjtLAOSbNACG4N3HV+dOy2wpSF0yM8RYm4BSZJpuoZGRAo3sjoDY1JmB2G0g2d
sPA2obqUgl9K9PZWu9U5SZFj1QzQsDZxlG9hk+63VoRT5nDtajNxvKvumZSuRra8
8MSzwnQr5m1t3uRxvKKAe5Wl2zvKM2o+h+qDHBqY0pFfxrXuu2Wtc4uw9Q3k/MBc
eRJ7kFuMWNBE5cRlMnMxWVV40mlKqqWkBrcbZAHaEC0Ajd8FlcUqBUSU/htNTgfU
6kjkrleH9hySekggU5IpGdjgOgBYxjaMWezxrPYUwwL5l3pBDt5olcA73Wm1/RZ+
Moh+CdlBfH52pvOQ4OKo7FHzLs8GbWKUQ6+sV4esDkxcPO362dCXvFJ01RsZ1whR
MYajgW1lrDCqtEJAxuMwOHhy4VnNFKYPd8YqiWox55P+yeTecvVG+VAzcJhxRT3Y
vT1o6y1dTaV7xhZN/ZAf1UlJjxju5I0XCMywmSnTjnhwESfqwbhntLw2hXHqTMnf
NyH2kde2XMtPPXwPKxSxwxtrvbyMGMVJdc8SwDdldcGOIqE2L/3SqIinItTnNgdb
AUYwJpdQuS0iBVDkFabpi/U/ZAw6lNCfZgZ73i8JbuRdWWL2PbWE/rtBD1Rzv5RW
ji4KV8bB2XGwVM8MVmilp/22l7JQFuPGRk/KHDBqPdHKPXPgqddijrfQtXKXgyCW
wu6cBHoZrkwpTTVJPsGI0Qo9xm/p0DRyS/ExDqVgKn2woDmRFVqWwtKPNfVQeU9d
Ycac6V5XuSzuzjUkvM3qTzssvhWbUVIC/OUOEGR4ufjUBzNotV+eO5sXEF5Rgoi2
FogM6QrZk8Ij8KWkH9xrBTN6DiYvKWvHJAtxyVL5j/4o2M6BN4PiG7Fg/Si4ftoG
8vOnNjsX8iubptJRxhUfewBU9Z4mMmIRnXh2LvacERguchkioCpFu+Tc5a0ShCaL
DqvcGvmWa0wBiEsNAhwVlL2sOf8pOsa5Xn/jkpHTl+29wUhwnk2SBFNCqMMe5oIr
KF+d/OQmjfKmNAQQng3dTlJ/Bfxn0xu5MU86DhmHnC+ShKkRgGx3oraDGdNlOsyv
1oxcDik/G4aPxocDRkyjUcA8d4SS2M4Kd57Qw/ZQfPkDWSjxbKjhLSnDH77FAGjL
je704yD+YGngLlYzu5+0+sZr0mkPzxiMLbnB9tTkzF0WGW6GGAuoNvFfXzOCpyKn
LYF3S/v4V0D+qJFucpFyuqwsePoTM2m7wnQfnYVMYE2O9DkVQ+kLDzATgP3hmp5m
R3uvv27VOwvD8258zVZA+yjisdyfKY8EW9JFalbvRAEzM10lNlysMoIg4oJv2OFK
tLElNswEA8EvP+K037mu7j/CWSYA8wjyzVDtvKW0vgZNjPJi3obmN+ZWD9zFtr/w
Ru17fLUo9j3uSwwLHD0rkwHPeUSl/kKAvoTz5aFjO432BNTWP58xK6s69S3TwGXu
Uu03PMrk8q/QEP8Pc5PRdhFxT/Glm6mmPQOILXpeX9ibzpohhblXsO2xRxngScjp
PcTpySKbc3LRv9BGB1MePTEYT0jHeC8UrzrsuiK5CQTb/s1YJ34yBxrxh681Nuto
iUApI3HNmob9QnOHSue3ftgnfjTGXUm3mQIclDV8Sszzc+KoI1kx+RUnBO4YnDZM
OZOrVMQCiR3quYNZVlMrvwaggbvU0HghDW2ePtY3EB6B6N22mepZjw5k7wQo56m6
BECK6FvFerZBZw4P/KbXABsIISQm+WJldvz5cAAW3kIO9pXMKFgfk0BA/fRu3cKa
HQ9tCRGmCC2CmkcvNg4ZOWNJWpyMS0nLx9qnwynyC1OBxZJ5J9kE0SrhL5aUzYUS
6e5aGTED0jtr1vSbPuxvEs+N5iMdnZi4kW5TCROfBndiigwLMj2LLPEUTi6S1QSl
lyVj6iPNQsHpLtAsq8808O1WsDo5RJuna8mEEN9UfJCS9nfN9E8N3jsBNruFFbEB
3hk+psgPeKUQv4+1J4zdEF9l5Iy6j6UFg1cnWcvhL/pNO+70IcqPLDFQOHf8vF60
VtN23JzbPIOEiYB6yWPykOuo15p5noqgIs3YY6N7jG2dbo6Qf0t1oKlRSPiOCZHz
qtWWLzEab1tGe9v0yipW1rmLfqDRueIXtfC8OJ7IufN5V+x+BWYSGTYOI3lZJD3p
82n8w5rlML6MlHSfXWtqYk1YMZjHVRmj45cAMk5C6TEKb/bYjdy4drB3Cx/3AvYs
1nVjHHZSlzKpgeckXm/7xL08S+ErsFWlCo21OduvbFcaov/sdgcVbWXVYI3lo0Q8
xIiD6Awgcv8hh+Eh2w8Z3d4c3fQwU/EO6Qq2kxHhJYrNjD2KIpeuoAoakbc6GVz2
sRrrZ/woxWndGJg2rcD9gM9cZHwKyZHVMoH8NS8t0cb2n+/rG8VjTnZXsm0ij3g7
XM3O2CCdF1aiWC3unSjEwupdaYqTykTBlgfMsEmK/4OW48nrG36W5URp4ayTns48
SlxCym6OEB5DGbnPY5ekXflhm2yng/mkgIg5cVlnY1kFVvbPDSFtLvhc/LScaBBt
FiH/JW3ARdDG2UQI7t4O87DJxPclF4bLXtsS2Gqj7bfubstKuI4We1AaiR5cRIUz
O/n5u3yhXdNJNcEd/p+oDs3ykBxt4iYHwoLZKd5dyP0XJ64U+go4RKccoe1yDF6Z
sTNdAl7gtm8Tw42Mbr/r11k/PgfYAqWvCiEgKab64a0sNJwjj950mpSvilGOubHa
zRZnjYRoZJC4bkhwX9EqN+6+wzYz3Hug8b0l3McrDMlcsmsNIrfUiXsoArbP7C9x
KjJG0rA8v8rqgSoU7CfdOOR/osZzi7sORQosAGiLsi4Q4S6oApxkt88uEMGPS5L9
YdN+lCGmOxHqlX6Lx9ygMyj39vr2Tyo2/cTfzLQ4pDl8HqZQQ9h6AuL4Y/RylG61
wUlZJ5k9lBHmJcdnfyxDMnrCfzCGhXSZiahC0yV3/O37yoyFwMK/tbqipkguvdTY
SEWdJ2Eq43QpvYOLsO03WROIuZu34gc0FHNMDCBaOzb1sFfOakf1Qs+3s3Unom5A
XxPdXsB3xHgC7TiBho4hFOBwqUanXyjFr9XMTEILpXeiCZcE3J2bOCSnOjjoB8N9
2hriGu6NX88dpeqQ57AElfyCWeJmrkwRugG6y+O8Lp3qVHG311vi9rFioXz4ee3k
CiM86RP1L6mGGxDRdBaZxcZEUtxsSfUf6g23/lVYMA6xiqX1UAq80RSg2W+j5MUM
nuOKx0DRYb559RFPJBpPt/+VPm40M9C4kjs4TVH6SJd+igzS4xh6AZvcWnU9wc+o
MR+HbIGhWpxBN0z6I+jEZiMYqF8X79sp4IKOuNU1a7I1lDvVl9kLbMH1kR2ACWoN
w8tXLEHS42HZ5fkRfcCgR4fUQquUZJpslJ+ExvixGo4xIfEuOrdLrlwo0ItA9iI1
sLotgCC+1IajKRSz2jxs7rxs26GmcpnhrEvpHNHqF+tSyYQ8x/WkAiOgJETFPziN
Q68HFO7mH6MRk+Sjkg+nLeq2FAJWKTKYYgCE8yUc5xEaLmGzSy1LejyiVFS45YY/
AqPsrpVtg+kvJt9RlmfEsqS7oSyPRM4b8AblSBA6or71qnoz3TSKrsn1GGdEHL6E
cMKfzn49MvUsikZ1EyVaReJ9GXu67rt35g2ObKFcFVd3btX+kpOCJ33pRzcEVT93
IxcrknrslFhv0vD94m3cUEVnCzggdA6WCPcnYLSUlbHtYJu7Zu4uoqHa0tz4ByTv
7oIEqI1NFMOpnqmGK9lov/aJZzWOr/wp2BDwavZwL6FMchhXWEo9GI1D651se53p
WnfJzsQFG4k3k91/AbDHY+Xf9sO7bti+GLP/GDVicj0r80PubP8l8XJ5fdoVWFDA
LBFS+5En0pOGuUlJeBd6DyUd1Nxm7HTpKuIS2KnGQHcFhRdild/qbFS/UgqD3v9E
31sRoHox+i5/y2AliZWE3NqBFNpoiHC6LdTA3I0dessxky/HePsGFhrtBTSXN2b4
wOcVWUZyYjZoJ+pM/Z0PqmzSKk5iVn20XiYNoGdvV+o/kkqLhEfP6euiXBhlkisH
MNVQWU1hWP30L5ZJqzVs/QZ9Gc1LKuJIxMqIxdB3//mzARj35u0TG/4SsQ6kG20J
FpVv8y7ypjFdA55OO3nlTF/ZjPOsSQW7CzIMI5cLZFsiItQxVAFCmR1S8VnP1+N8
WL9W2K9i4kUPWaxoQ3SL8qvneo1Lhvy0Ga0Q7m56DK9vttIFXhfi81JsrUsfFKs4
SgeXfdP/y/8vTwY0UNG+zxPJsQb9I6o4jlxIwU3+27a2+rlHLgM+RmDS6KDi3XRO
zW7R9QVWOQvV39Mw4DKWvIS6jLL7N7Vi04hP1VkuIncgqZ02Bzb7S2blbo9jD624
wTP2nnNnMG4PUfmc15sCsZMxVpPldp/R0pEUjMncZ3MRuoQE63AxdVwWxRetK00a
6eDNGJ4IcFtcujMJScvoIJVSQ/3qTMqXJ8wm/w4JtL6PUfvoxxcNv7eJ318z4f3p
bguaJuYL+w2NrXknRlXSrAuSbHIArtrk+vwn9SfhOZnJ5DB2UnJIzMLUblhP/a0T
x7n7XT30zndsoY5aFaTMOWY9PCby27A2a1pHGmeJ4/Noq6l36BaXTrMInLWmfFGG
/gIa+jVuZsy7tOpZHtJI5RZ41W8zSY0PY50GrzUfJH+ExqJfvpxRR3C9xN9IJyIU
97pLCeWex045c79evJqXq6ZqYCgpAZFBr/XnjrzdGYrHWw8UOHJ6w4xfmkMRDQ5U
W6ZOUyF7kqVwYCME1JtdR/QOQuE79y0JKErQiIBCP+Mj+vVz8JXohKnLf+RHo0ON
L/DeIW+Sy27Z/keEkU/dUZl/BIKf3iEwY9uS6LRfqT6vDyjhbw4ZZ8H0huxyfe68
`protect END_PROTECTED

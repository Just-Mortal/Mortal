`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19dwlYGxDKJ57ymOcIqRI0X5zr3/pvnx7xaQLQJRlZ4GrGKd3NZpLjm3Yc2IH+V3
yAxpa6iusmkVlHVIoJIbRthtymgUFZeJqOofgHs7aX+xS9Lt0UI5o3M36KlPwdcg
VWWxKFL+dhOO48snET2lnIrLz3AN/uR0AV3oeqRJeW0vPunw91MH7TIk4fIXOHLT
la9scWEFng1YBR2Dr4wjukk20upj+s+LIv4wZkHB0W+dl9nnT23FfIylPio3UkBa
U+Wf7uQc7ozFqnivmO9zNsAmsJ2+tKYLXXefvB6uKapF+Rq0P/9MK7Tr1X0JsdhZ
zf8wgEF13lLtHxhgXfz2tN9t4zf+S7UppBdqZqgMgO3hFpOUn8qKr4Cq0Am5Qt+N
duk1+xL9hFw4iHQ/yaQYrMcf8PK5Cx5q0tzN9aPj/2jhAS03quYY2DvCQlQJEiBd
p/iDpuT5FXFB3vorx4n7Nqm4JLZwGEv6pPZai/x3140NAe2YqK1sDkwULNOfv5LO
IjGz9iQhb50xdlpJn2U/Xg==
`protect END_PROTECTED

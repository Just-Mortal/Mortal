`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCmOKp4wr+/JYtUGCMxUKYwDi8vS5jPSN3M2EAw/3r6dG+yrDLM8Q/bKtcbTUB2k
eEC4jhAYYgKYNoc10w4zuYEahCduDXH8eQtyhUevpeJbgKEYEcCCfrSXCUmBfAQq
RYDFnklSoI439BXB+yAtHGz01qQyKCp2ze7cZmkLmactsI+2ODskrMNDHMBhw8wC
Bpqe+ln3CAe06zslMe+S4EMhSmzrfez6n7pp9pmjOO4DlX81jFSQKK3G7fwJnLrb
p1VKjjYZcNlJIFrfdKV7N5jvlgV4SulT+41N18BSrhBxMtw+KwUsDeZAeahCjROk
UNfvBjtb1JnHumdbC+B+8zfWgZ0WE4pVFglpypEmkTlLa3Ot1sifAsibQFE9fNm7
N5ikUBLa73Ekhqw53O7eN1CcsgniIwY0Qwuj0/T//UvZkTTf5a0X6sbMeuxjArb3
63TFeZRV3mQFdAcSCIovJVVTWNt4vfKLF8rS2EZkgFCv5citkGR71n/6aM1JMTgx
ZWtkQPsaPeg5iwbLgDrJbZPqdmpL5cQNmx+sfP/YkFAVEYEfQYmDbVpTEidvGLbh
LThq0wo2HbvgTR6TBz6HJ2SisLasD2Mw0p4TIfJVjObUjQPelrN47q8sZDSmsFS1
zMVpPRf1nm4OKCEuKTF+722pUfjaImzOgLWDLqO9SEr2hUbUuIgbbXqj+Cj9ujMx
Anji5EqW4gqpRp4BkocR5nOnvpsbowDB2YEtyMMmsImsqTvBQammz7ARmtv7BxGK
d6HL7xxX6JgQJOVuXenhdBm0nqNbDh10Qx3nuWzSqq8zqtxGZ+YJ86xQ6nBcbVeN
4FIo7k3fqFNovBxzP22ubEkTGjPhMIq0oImoJirqFHYJgWTzmi0dhMuDYFG/Ic1/
JVSrbK7ehScO3SYOzV/xrM7XCpCP/ZUQJhwIcVJufi0AYqEMlFQhKfRTpoil8+uS
mv9ZtS2a+EHPjVfZhlNxnmU6nAX1d6fWEwn95Q4Ec6L8uS9M07lN+8ZA277EEtWF
25jJFGEUESO5Vb2QHMVTBFoBE6gVsYOmgCUDDLQoCreWq6RSrFwE76zrbQhPLCS/
CA8cpS99XEAJolKKRn3Ku7Qj3IteaP8FHqLe4p9w+hMb0ns60VjY22mjd9Xw+pS0
zVVOlbFmMfZ69IBtDYvtoIbHzvRq6cLIKPvLTxFqpXcgZOLnOXCUPNg3UJNDWGSy
1JXArxt+63TQPdsbSSH5zcwsdzkbULqYOljCpjgdqShYVdho/W2UnOR5azbmg1tg
bufCZa/7MbFU0qDeC+SEAkToXuR8ZPz7mQVzEyzlEf73d1xIbdaeqmgc8XzTqbaa
c8mSo77hjofZTTjqIGrIfoYpgGGPGGtxolcaAuiuVtiRllh0h0PX/JeDYWR5hqHe
0FFY0V6KaSfpyq91nvt/gImQn2hPWXdJTB1kohYRP+CD1BkCzW79K0RL1EUOWXWS
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aYy7admIU4W4kMdRJJWXCDSqpgkceia2vQ6i3g1+iTxz7S36faPf5qvAIgsZnj1z
cW7XyM37sAPgcffcZ8GNYDcY7gQbD2a+DPZsQ6F7BPPcczC482wV5zgJMQpPI+0e
pf+rBPln5DpurW/S18q4rGRgm1kFezbTnZg8H921v1zO+8l0dM0TSq4tewAWTCoG
sh9x3kLckfOmcsi/z7aKgaspcClS7AMhmYnFM2oNFuhhVLZWgYWA4Rp3ySHViijj
cBcEVPV3FAzX74lFwA+BOYwNuhzYVuZtTq1aropGdlasdz5HLgeJKOskxmG0AT2e
R7gJIGbMcKL4MK/xHSKiu7sPpDt8NCae9A1U0ORWu6DTM4LfZzZp0YShnIdkJBYL
6za6WK8G+dV/a/pThcSrkzPTsvNNaNg7GctaYk5faoR8C1TvSm6a6+G6P+SYhHUV
Dts0LSIKPHtbHTDeJMSdE8cu+litxXwMv/o+lEvNK0PqvAtXJrT2MA+wWetQkLqw
M0Cw4pWECaySOYbxmzPOvlC+sMftmbnTSvNj0u41O15QpW6apizyaOM3p07eRqhE
nIO7Ue0QID6aNYK9jgPwij0tXGOK2OVEheyr6qXoovt5L9lQMps9On9f0TjwfvP3
TaMMNwle3gPBL5uR3a2Vlac+6T8pGzprheQ6al2ZYAHuFif1ivkRRmNyz1v7oS1N
0hggisKCs6GraH3wgA86ys3vUr/jGR9Fbm8o22Ott++vTr5XJEzlnT5DEZpxjsYN
YlpjKOrgO41O7k4dq8W6GtaYyjvBNP2W8quocl9GmYOFJsElEg1mBEs3lwsV6cNg
7oKf4R+n46dFSKQLAzDsYTr1BE7AvINB628SxLn1475YEk9qFPJB0d5cj/+srpFP
1cTtUM+QuzHbGw4OaP5W9/PEd1IHqjrVfKeFiEoEWbXJnFowU4Dc+xLyMI1o1FRS
/En+EcEUGAKbzjpOlk3p8BDp8b4hD3Ey+KSqI4foh/06eTeTITuvcSde//JOTjUg
DLbKDH5kLLzjPM+gLEr72ohoNC63rlG5O8FlnPOXpLYeCsSIgHqR5+ZawEsPDg2c
CSOeCCeR5rxTL1/VNGVmy6rJbNkSW574EW+LFKR011h45Zg/VhnSRzaDslO0mTn/
AM5YbuGiJAVnCwacxgvW+y1v0fm+6MWUPaAbVxm/6/AYo9b3jwTRZ0U6xt0Bjx55
c4SS2gWGwJ/6DB3Dw0YEhnMcXWdtRC/nlO9ik4KdyQL+7V5uil4RJYsL7JDSiK5p
7RGilBUdJMtdx77nUbqsmWwAryMzp1ocSSo9/Nibtsmsp85dc6xSvZjetU1LCAcE
9NLwWmke0Mij0WFBUhsB8VolGtFijnJ/foJILml0/p4bu+zrdwMpwt1MP4mIahk7
LHlHGQcTMoJP+n7HpI2ktA0mo+hyzJT94E7lHCjZdVAKieGWjVxRtYGmqLYacTm5
bygWKtUvp922oJAKhrdF22faqGchBzzH+6OMJqQthiXHVI8PBpPaLTUi5HQSYOw4
dc364nhTrCHOCxClVZz+Cto7weL0rykt+oCdNJ12axFEA46jVE9ZMkphLFX8/mG4
3aS3flIE67fDvMIiIt+3QvneQJRkGEye99e1Dd0nCkF6ztMN+7r2SMmLEshkjIzu
BurH2u0hUVVCUqMGwvk/30On+FMA9MCBuNWf9eRapYeLGwQPMVOaPquk55NIH99O
MLcX54bGn9B64QrS79ZM1Q==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CAyHN2Y5kBBKFMIVEa8ZnZhQJc9mtC0shvKvp2VtejwfeiXUkl+M68+CzYqNcTE
U18WsQ6Xn6q49Sp1xv3LAkAkzzCqnVOo5VqagagOdULMkwG5m66uvC1LQ6kjwzhi
aM0WWttNqFRu1pCaUgAWyGZEwmpYLJxe9YfAa6iMA2zyXjd6KqBvUsHLUR3X9VA1
Drr5jrcFZF7MhpeXExZNXCmI9nomzk/GdHWGBB36f4/jQtKhuzTn7lxNQouYXi96
3fYvRXK77NNHZ/5Sp8VImpqcbiwcMUX+cDe6lhj6IN5KNAOiSLifh3+aBHtz2E4N
6smDr8hfaBIwv3IHqZQY34R18OXzmMGDq6Qp9Il/+urAThxzelZsblq2p/grb+UO
`protect END_PROTECTED

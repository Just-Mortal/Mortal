`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JpSGp7o/lKncg4jN12vPfjFheubLh7nRXg8MSKSc1SCRHQMdpHpA1MmTL/LHDizR
PfMpp2jdiaqENqFZeaMsLJJYkGB7v84X5gW58lLZVFJ8HEnPrOqIFC/UCXI9z80U
MmkkwYfDKAXhLVnkBbnN8cOZ+V/ZpSbmzVRjWaeKXGuRPCJB7Bj/LfYEqhkOkegq
E6qSflCIKVjpRi9eRCgUmhdDpF1kwf00D1ANbOOsgcpe48SmkBh8qoq8iFoxaKL3
NuxMCIorqjj9BYcMZRGUjsCi4EmrD0zeFegWyBEPQQfF5BM61MGXWSE6gaeynSVM
K7aw7wH/iaU0kOvP2eAYvmzyFM6bJRck81tmh/DQQDsw8d3uGR48BwXncvfCwKrW
RDOj/Wp8LLXeC1AJMs8XSmU3ETQ3ldfgBvo1Sb6nepxRZPe0k9FMBvo+GiaoTWvl
JAtnWsfJCOGsMuxdtQiOqzdvd7Y+8/U1dPBywc0J3ix6zyxHR4cWtBwWpM3Iqaa4
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vELXkaDzyuKi3EBO104Tjb0quEse8k0iWuj2+NshIXR6I2VuWO3cjahq7K4XiyRU
/Fg05Xcy1iuAHnqIb50TSFYgkUY70NDEBbAHr+ta93cvxUEyM2zP0wEDonphC+ul
kXARxo/YynvPadHI4PNw5dvJDqQ7qG2L0NiMHtgSG85yI98bzYRsIHfWCyHVG+iy
A5aVQFCn6opoliFxD8SDMruNZjIrBNDB+kcaQMBM1I0IW7nzNZXZWWv2e2MyDLRC
9Y9Vg9x0qH72aK7b1GZLAS+XYmSUSJ9/hVWtdaePJ6T05XkJt7dyLCFC0wS5KpgZ
ckbD9Mos5OTi6qmFZDoUtLwZE+L2Nw8yoPrtPa/5i9CkmTtH/gaZ4MK6wjHw0UjO
izYt2AmTEw5k1T30yh7tUPTOyuJhanqxDFdJ9sJ2QdD9UQWlAiqpG9U70ZGyHsao
gpGjgMg7ZtQ4i1Td52mE0Iv3zmLg9ctEVr6dJVCrcXGjlX0RU40T8kSPFTuGE4tE
xph2eACDdEeuGJxKBfV+PBR91bhdPpbHDp0NrkLyKbkyaN/DK8W/Z0g+SRPe0WjI
34DH0rYYyfsmGYh9vkEhk1K9hP97xIs2drUNq1JYgn63pdWn+1SSoNFMM6mcMY13
aDl4djq80loGO9H9FEOAhV1W8U5Q6/IS9c5EQxMHJg/DwwRGsUh3fIgXUwbwbZr5
MQ1BaP7TfMB93muhy4kzFAa0MqxIIkG5Ii4BaVDDe9smc7Kv4bPJTI17uK07fhq6
7AuWlujt2kW1ponXFBycXg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJrOV4o2NRFMEZysfg9yHYIMFI9h1bPABcWCxiyzLYWoGuncehffvkEqsVn5wUBw
f00szSranCqiS+wscQsENGT2J8RlCz6LJbNE4F+OrcWNdwqHMeeYzMBU8BJsC0yT
H9gy53ZcDaEJKqa9K9pxYnjEbOhUdfj2weLfX9ivzuvZfAj4vrruo5UufPIGwplz
40uyXa8taimDT1X8ADArPfeMHmez8X66HYJHs/Hy0lzD+R2n/4b9PZE2fPY9/fwr
m5+wyrnTG71tAsc1HknW9XrsHreVatpRGDZBMButvYBpc6GrobzeQp+8130Ubo6r
OGvO67xPhk0CWFkSqO+kD+ba641akphthzuH6A9u3hXZkFEAgZQKqJ9VdRtj2Qk8
haIs/2iiYrdqAihYPL+cAfN3WLHbuqPZfOr0zJMgPFQAsZUum7tRGC4nrBac7NVw
tZiszgDJ1sybMDiIwy6A3D33MHUag0RR0AiFXT/VafpCpP7hc9hco36zaK/WiIYz
HBa3R12lICaovBIGruq+jjUxVUKCyRsy/Yrk3hD8aaJWksp+W0aeUZT3xWbyhe5t
+BxN7raneE2AqDZGU7K1FdFWL1NtnJ6MiFrSzvVoYM1D4v9ZnYpeRqzbCS4LbesB
Fc9g20+7ihscejVJTLH9k3hMpZVvMR1oeRQzAyYIpO8dcXCd3N+o2/JKGPC4NpKB
m1nwBacDxoMx73w2esAxz+Z+GfkYpkDVMCw/7wWxbCPXI/SNybHf+8aUdrU7drKb
SN0GUD3oh2Bbnq/i7kjivsZvV6J7sUzT3AXxDL/+L40CDQbNDShIrXq7zTaXedP0
HdbS3c1kSvhwOK/Q5tY7vDhW2r0qnAEg2XBlw7y10AApycYj92pFlzFtHKF/c+He
DbVd/F9xAFXBV8pCV0N/IG2OFhS0si6YtGI/MXOvVbMrOyA+u+trkX2vbesPUGEz
IJZ5XmR4e8QF4XWhZ1vNfYsz7dNlRhOGviAjcVdYIGLkpLXpz4JezqpOP2EOKqFn
FIdR9GKycYoO3g0hrmYW3kTN9de7HQIAob6q+RVPEDiip1oZDC7w/FC7fo6vCLbs
3W4OMYL95j0BqGKolY9tjayJYeKjJRTsHqm5XRioYbd7ZMC8yB8bJoln7jrAEaJG
YZoBUdKOM5TPRQUUBY/HsBBm+qzAdaERHFwb36vC38mE4UIpiFX3iybh4+bV8IZ5
ynb0z9dRmZoaMJLclSvo0csZ6qRHjjWMwaYGky3aTKhPLT4srKN6UoW5QIGG2kXY
U6Ieb+MUuej5G2dWaPKdUTSkWxXmfqpL5NcgRR3Gu+K6JkD/UfjiKGYlEHPalkLD
DV5/QZu0u3vXxEZ2dR563rjdInVhEPn2fX+oYWJjdQRLZlD9YZObFMO5OAh0fVK0
c9pZcjcmS0/X4ShIiTi+C/vfrFNMhr8ZI86DfuTU56cSjIVy0geBLtqoLv6I+W0S
HRsvLIs7zRolNisz61fnVFMqpvVneY20yygahFp+/lQN1yPwG5V/te6dJCe9E3V9
XJW5cZn+TELqCRTZmc4I3w6kKTmymDKeVqxjaIR76cfUTMn7MuXH2Gvjxlbp9RaY
vt0ayDoC4tzD4WdLOBkstal59flHITh60+ny4j+dPMMx91dIo7p7UXWvr7ZEDkDm
UsIgRxaYsKYnhIAheWAnXjoZVHmukPDGUDKAZPeuEn+L2Dov4qGOtBa6W4I51zpl
4eVNCa5eeRCFCX+KYAkt/xdrhXo/2xNto3QPZElYay0SYwxn7phW6PEbSg9xVzaz
dYIW95eBhEiqPuj2NJo4mEFeRdeAgQGD11B/8inMpq3u50kDQ46qOXDO/ptJU4ap
C5Vx36//iwl3wXb5FdaDj2ZEtUv18UMVROsI+IC8kt8Dmew4pYa3c25LXZfp6DIk
rk6AXR2dKmAj7rcGcGghAKjhGlx1DLlx7W19l/EqacY/oT/y/xsL8X2IXQU0XDab
84W+Twjz7Q3RRaQeDlF1/bmcl/49rAdNcmQZa7PrzN8GGgMlQaOvl8+SSxSM067E
tbvJy9KiLles3rI+Klo6O+1WhrBFpGiSUI/1UVqJ6wmx8adu338yCt1J2c6SGwCd
0nLKa4ECD4gvSSI30AxxKSE9sS1lSaNJq5JkyA3dmZjjPPOUkSH0xPxtD4v/36DD
9kZ4QNj1uS31Nm3sbeLeA4GdzC/Z1MlC43DOXepwviDc4BbOEfM++mElHR3qayOZ
cRH1d7QaJ5Yhhfu+Jf6poBJeFz78aMJAvHXeyMONXn6vZ7USRJv6rNgqbAHoX+aU
l9g2lrmJThY7h7yA+kV1k9Drxr0MD4zqcUBEzK6CpggaRKrDgYI6DI/rYdHF0fSV
4wVoqM+D61FQ5q9StEshGYN5Azu56nKk2ceLi89TymLd8c62LOo4RWQvC/9GRsCF
UjsavJ72vP3WPN55R9rA9FlRwRcdU0fsEL8eCnX0746nWUtO04ZhHN0tDA/6Wnpp
ZddemcBVanhZAT0UGHzdDxYL54ZCt30P+iiMeXXXdW1fLOgEF1od/AH2TArLI3hA
50I+yRuIOkiEMGewIVU2Ut5rl96eo93Dz9LRMUQVqkO2H6s8/Sh3VywPeDG31eN3
oX5OrQlzKqhx7Ck3RIye5RvpJtrTv/PqlPq5anTKh6Ku2drV917mgmMaoPCJOTHF
KV88xdTtgcVSdNCCcUf3SXZ2xeb7MvtzRTFY+5EneVrLS0DAdcVzbVoYqEt8jScD
3GrxD30GtoSU009QGgFhPiLUgALcxZKmCKTqsoTspOHDF4RF6sKZxI6Ep/5Wdzc8
qX7RLELJMovKnW3FHDh/TW8T91SRavWWEM4KwansqmoyiXWrvCismLGB0cXjSLik
9NzfeD6NWY15FsmtIbT8U7a4MgJNcUauvpSJThYoNxANr8jQ4oHUYf2S+aZmWlsU
ykl9C+c4JqLBoHcbZglYyxIIP0x+mdfAzEIVDFMMzJSiMHRk67v4or4jYJZTtsSZ
8H5aaflSWdp7lOJTdmMO7ooUNzxgRJc9SLnQzaysGIO88+EBZrckT2z5wuwc7qRV
zLuzFR7wUw+RXvEXM1Z/yW6yFp/pbSY23DhJ8lWjS+JlJ7mVdloT80df86FtBCVL
ThhV3euacWoalXw1wl0z0J4BVsFPrNYkP0yNXTfEwvTeao9DGLwHv85g2X1EgL/P
pE8+5QJRoBp5THy8PDCL+gnEN+mXm9dn3G62EHT7W5XDWDuOp3Dw1Wxr3RbklhAr
2FQhaLqLEMqGiXiTrfLRyRwefpYHQOODg8ERvWJPNFj4Rx/goKLdxQPzxCy5NX40
iN2FuNl1f7/GAQirIz2gu5Bj8SX5IDItDu/uJq9Z1WgYYs+GEzFlbPtzPMc9+v4X
/U4SFQ6yJcte5S0oGZ7ue6p1JqgCBAOOLIXegsrXTVTY/kJimRZOFPrwyDXCMVJM
eCKIUF94asICKe9AXDAZHzISX1+3wJasnk3uu5qmMKyCRmBqS5zUNAP8ue8DKZC4
P3Wt6BYMwwXRg4qrEsWJLd8okS4HktFDGzxqaNKm9dqzkDKJxQXSCSB60W/demv+
A5IZs8Lq73uBsiZwRdknOvBcaC+WE7Cj3tQ61bWYeR4ByixvVAzqYgBirS4wV/Ae
am0L7FloVe5RpSwb0/mwO5N0B0KNY+Pefirlg9y3hcJ2pVTtmmlwwSRBgDVo1FzP
KtQINkCgSbiknfOv55I9+SOy7xoqh6aJswE1ZU+7btTapnzROGP3Tz8M6iZbVGo3
3thOG5+gdECIkta5D/ul0XmPrzOjNYg6SI3A+nAsBtgXebALBpg5CPv0OBNN06j1
wvlxsBEoubO018aacXMd8OAhwRpBa8bFSehBLz4XJRX0+BOXIRwg3qzdv6CxVMs2
GIPkFhPl+MssYbiai/W2iw6Kwns9CFpdR12gnZ5e+OdGkfqRuhRBuEZgpQ9wAgMV
7B2tBFEHMuontLuQHfuS6ERtsYqthXtaRe7JTntGMq1oj2umaVbzjpXRiML5x462
K3rLMOWfpom4ugK8d/aDSlyIMnANQz6Qr2BaP7NrcnO32ZUqFb0WdrO3T+I/Y7qS
J9MW/2MwNKPcx7IH5Xg+IsLonAm/Qwcm16AwotD4VHofNT8WoIIRhoW+ppMJdgIm
jkYOpryDIT8RA2v3ZtfV8v3jweEyqFwb+ui27HPPHzDo5AQrC/FaiawJq0K9aP5E
SC+FKUArzCXohVvSzrmAE9y77szhykq1iCj0kLuZ5qHHByiwy/mpMhNSxa8BgjaM
UNArRkb66mKBvciYbrleOHgbkAEiAxMFoCrcwopA91140mz3MLaGkd/GeTjL4Kdk
+sHTezZ1Y3QG4fky2ALRCE8Olu49temQlDQOnaN9YPtuLYi+9Pg+92MldwvwDzm5
of8E7UAuo8ySvMFCoDegQwMFDgzlMlvnT/xodnzr7mP7HIk1mJt6l6IAt2SKmaPu
4j1RSHaQCk660LCwI6CIl35b/x/pqv3fC03gVgDn8m70P/3u+zHmRemUPTMSXWcd
X6UG7MK+MbWsXfyCMIuRUN1pG2qY4xy8iy4rPrMaVLz9kHRxy3pJDX+rKttwIxN/
waJ123vrUhcqxVGt3N6Jv/63IP0/XdBDoFYu9W1Z1br6uHQm+zcVbaIQy6cuArfe
6UzLG6mfGTrbXyPbZkOmju5IzAYBYLL9x5bUvH/p3gm0FIgkfYNtIQfwEP8MeKxH
3pYMYjm/7+eMUz8QVy0hprbwVxEsY/twHQB+/ptuufvDwHLQ1Rw59G4UxkAJFlTk
I/cAZ4nYNqxbbv6kVzgXiktG3xUtdPfeQP83vYvuLJs9pvj++nTI22HAovM3Gr3B
8VzFmBvLP+mwgjRBEKbBrvzfiQ+6hlTF8PIqcQlRs+R5MT9qSP8gX6LP45j4twTl
`protect END_PROTECTED

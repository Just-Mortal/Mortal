`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e9gDooby3FRHilKaJ+avT23jQfBYWI5svqbWYXFMimP+hEm7s4H8reJvqC8llmZU
70K/Xb6VTOYz2rtUzJCMyN0pFmr3WRXFUs/JfQzBe5s0Niw0FTge3r7ehJ4wBtV5
CnFmaKZ1uL7WssiiDWWvCL3tVw8tc2ZGVDjQvQ2NyLHkXbKzMI1OdbgoMDnmasy9
vX6Iw1Ji75G/d/WSRgr5e5oqI/EynQH/GmsiSPiwKN1CQEzo69ibi6jTsrL9cu8B
moG1wnaZDXK9ENkXByk93kpNf+wxIbyOFuqXYZSecEHJkE8fNV8+GxeQlO6EILyc
6PVMA9hSjduUZ/i8CcfdX+yYfHTyKZcCh2NIS8p5DFRG1w1Yew/OZReaIjclakLB
LMiCdOA8P3YqZq6EvjnnTl/E/j6tS30TDI9BhpBdnJWZRJBjwNYGVoFzDCzqXUsW
rCeCGQxy+P4EwjCg1OqP2kELvCHE4Nd6CnQF9YpZY9CXXWxWjVUmkQhBti9fwG4j
`protect END_PROTECTED

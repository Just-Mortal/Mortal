`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5O7+YqPEbJylu6YLgmFA/C6rtggGLPKYTKthpJOZ8wCeumodwQB1qHtSuhh85y8l
gu+xq6VG+pyM5Qp42S5Ip7/D+tvee70cKNagAA5OOCdFgvpu30aCKoIYfAj8ck84
TkInnDnVRN6pEPFk2OIGJCeRETR8XprR2yZnwi1GxxtXG920OPR9mBMdQfl2HoXt
RoeKVBkc+G2kNQ8f3SPuav3a/yhu84qlLN8jzasqAAXVmySt/rLnQTIUwyG+eBQK
3ky6UR7xOOVzeLCA1agYeeSVPsPbmr4hA9qszZALEBGFdC+VGMhAHAIdMfNxBld8
TVvWcEOUOm8mrCKVK6vRF2uen5iVUEjM2xiFqiU/U9Y/cN5xYN1wxtc44ROGo+RD
AuSFDpgSvxsHHhpKQnggN6QnPWorg/FhL84Nzkqi81IICOvDf99nVVCjRjRXikAA
6mDhHbHLQ3qg50rpMcTvmzv/JfclkjaLhPk/WGd1kB2rZXLq8yP0mVz5DjY3LJKD
bIDhoFrvQ7x1Q6owByBKV7JPaHOstG3iPdpQg/7JT2DB3FTJir9AXa1x3UHIDPDh
PqKjFomN3Jm17/bdont9mlCPqxhytuTStBOGqqpVD0JA8YCtyFmtoce7xzuViKMg
d4cKSt73+5wI1FxOonIKtmayH6qx3ICGW7tZ97OE4mEQMjz25YsC0Yz9/p4HZahg
i158Z63xD8jwgqBfa6A4ocJGLXF9q+mkBgFYnesdcUYc+4oRGBUVGwg0e4fDCC4t
ZUhDdV7ktgUo08xeNcd0ZLgfjIpnDQbY9uZogg6M7sqClXcsvmwFW/dbi4C4CEF1
SIBFLWtMGPlbJSGnUI2ds6tvTZnQh9USwaSaBWndD4mb4qREBFUp5ELe6BoJJ4s0
ya/oERqvqj/8GHn7dCWeMngWLnlF9DgB/rFs4yZN4QgKcm6aeP6GozkJdmbkF1J8
/G+LR76k/Ruewoyca2jhrFw02h6sy+TN5RL/bXW6Tu27XyQ0iluolwThghKSvp0g
dIbMnwGOb2GW4vWke/09OmYjjiI7aQDyfcGs7/3zaFUtrtbZQASgMMsK2Pz3qt81
lSOpW7eRJVPvqyW628UB1nzs2XxSs0LeU3ovBwDRs7pAkO2m+Yy2Q9HBdhidNEnQ
5e1qel3UHKCuxCc/9FxD0G1EpVzqSUF8kd7fVXPd5M6Zr+K50CIDyLJkIaa4OuDQ
L+KsGX8wiOJ2dWminYxzlLtqdnFW9vV5gXwJIYHywiLHEJcIajhh2G6heKe4nhw4
NLZur9BChlVMC+s5FQrU3y0Xvp5/TFOcr/oyuo/Ma5N38cEQbIZ+XfGImDKYZY7L
iXW18tKsWsza7Hj4bhwbRQQI/a6GM2+lwGo5ucG5s+dEaTHEjrJJYAwLZhwoftDX
dgNX4FzQvld2lUC/pZUjv4aJDXNrdWoK/MReZiWop9cwCs/uv13WeTipdzt/4g2o
XISVB5W3qe1g5N8ogYpddiZSUlJXin6YCiwGvKv12uNgKQGXgHH4ngeSqTUCNi+c
TZS4jIlPXaOafI+Hz16Opj/KPczVhvugLTsHB4QhWLestANeSCGJ5vnElZqxC5c0
u1z72nzFw331yYHKM4NQFmqwYgmk3kCftQeyQO52twQBhSXc9Zta+zigPfFpS+k6
XFwL1McsYylLElppZ/QJxJvmbOgWXv9dxDntym5pcuRLmyEkfIbZ/xePsFkAwRHz
AUmgTWA0PoguNPbg7QZWGQtf5ZDXRRYEd4/vCCA+DqmnJfzPGWA5ed1I5qGitfpc
OSCEQt0VMkKxWc63Wn/3bgm1jxw1sTFE7OocvK1up7Km0FLdcXHHT3VqnUbIU0vM
iYytCQs/HC+A7eUz1yxYAkHUihd3Se/oPNjERGqn2M+bPmcN7TGFPfS5LnTYb/1V
1sHEUUyPSQwWJeiIDSYnuEZ2WoyBl+eLG5qqmqczWc8TaCXjn/j+qGwdify3/7um
M/wIi1I+nUqHtVuEAbAUYoQ4guZPLYXabZLkpgm874dygWtKd1VpHeogZ6cbH5Hi
MSr2zKJ4jvtLEXYRH9+/u851WJDhVz1K9slqcVDzW8S5VeCLccuZIXhPOYxmahxB
fBeuQqA+ZuVhU78BU3kPKBVewC7nJcWIcJqiSkG2GwQPTKkNVlsmci+piuvw6lMs
MUCD763M980LvbtTHi86go6RhNFg3ztCEKTv9hsQWFQIA5DG2VzDi8yOQLflavub
2pk8RV3jf1cwpv6ojHzHulOtfvkuovT4WiHCf8fW3CdpX1AqEe3AqTpoSnAuHJN3
ACfZhYit9A9z3zEZFGgUkUAGmsIN0vQxMLoiaQ/nbjz8ZcmIFw9/aM7N7RSCbAvS
HQFfSOxBfmt1at/seq2w7iJgXnvFetAapD1aNcXntlUn/V7uucJqGH0NHXU5oZEp
/WbkEhNiJx1cGxnZp0QwwCnNxXWEh1dZzTTuokhgR75JFJOAAaW6kufp7A/el7dK
dhWfLa4M3tAjVE1lOssS1koAonmhC4TvfGOdLGxOTycA6LqIgW0m5EGMAXTL/Fz8
t3rGG77/42y1tMiWq+3OC9QavZiCxer4w1naX6wqYtZnaXdYRB2uUXQw7tfOjiGo
lzwcJd5gbM3N+CwmYDovAPghsSym0kx+qvfNcENE7jLa8vQFBDKPcWMficDC3pbV
15lJ6azsNZthOK//aNaA+2gful7vR65ZbVAgDvRCvIblyGEXX8D2sQyiKUqUfP5c
v/Y+W88CgM2jxRIO7oPcVuJOev8nfxtIaZps/y2w+gp1mAgGXOX793AmeayuNUK2
MOTU3j23HErnfBGArDqvbBINmM0keN3ZZAzvxfyJb43RMreA0AifO6moj6H9VHOD
wBCXy3Ise2/cL1ez22D1ah3iUlrud/9Y63PxQcJZ3WI3lgZHs5bCiFwTFBl6tXZP
eW3Cdz+OKanemir7qKCLtOyRjRF0bd4LwINOrdOLbYzTcSTlI72s0E3QGMt2/bK+
6bfX18ZiWBaUWtMYNMx1ESysyCgzGXgqyUnC0S+otGHK3nh7LI/bnEhOKslYKllT
PqDP3cYSJcWdT+NX5anHCmJAz3lm5BCA52Cf7GiGyDBRRbnrWVoIC4X0jyx2/Kja
1h6a/3VF37sSns2ah/yH6NzquTiAV5YPzOUtXO8hDVI9n15MO+9j5zMyr2Z4Opdg
A3D9QA9OAsUKe21uA07zuDW7AQOpbCUoKR2zAs3gatqmqynndXXLcRRuWCIiWX3n
jPKCSfrP60Accq8MXGIuOoglmWTfIEZCq8XrUDRPUtQ4RJE/j8WlBlYpr7Sei2mR
2JgBuXUbI1bEddzqgMtltd/diu1A/N4cJs3pthLArrjqV5LZPpT4MTONBIQZ+qMl
SQJbnKXV8i5mfpHx9w0A3tVcU/XFiTHnty9l+IoYiSkvfFOyEaAm58G37KESu7+h
FKjneGKlvZ/rdfQopzvG8v1FaELinoat+RQllhcXLXCJ2EyPh66r1A25w66jvHK5
Y8OZq9QOEIzfz+YQjqCz5YFJ9LcgjDC99ajgcNrm2fm/+emHkISllWz2denhXtN8
Pu31JRxfPSLNV94w/3odl+MsZ+lbrBX+6DiRkjr4wo5rOnWHORTpQS7nBlWak4AT
/rKXrei8IYR0awfHrYZnlD0uDTNYgQEeSe2jQ6TpYWRgv9A01euotib36qJ0gJnm
QXYHUneZ3R+TKV9w5NBSMQwb67iGK5r3gO6o2fexA5uoYtpeqIZfkwtLOMYNATkU
y6fiHZwiKivhDweLDgnkv44nzM3YfVQZno6WCa80QxWp2QCt1JCg75mNmU+y8bK6
wKlEF0S3CCaxvfjvZ8cKGtyjDIkRnQ9+aWY/0dm5ji/jLzOXxCmadNzQiRICR5N3
5nn5di0XY+VjJNMwRO7JGnUJBYSCbJRqAWJEA7rECvJ+IpYFTJT8LUY2G4dL4gbk
UAHRldVwKwnSXyLJT3frWWzpu850pxpQxn56jXcUsEOCGAj9lfxh4aTDaNKIZQ7k
XoCHd1DXKvSQJOG1RxHe1ybYWjn2GwY3kzOX2jVI/qMzCW7tKGIROYPtC+nFCZHJ
bVBJIKbwadQDsd/eD4jIhMNx1fOkDhdry9PZwFFg/To9BHi/g6FEmFlCT3j4nh5i
n0LrDV6Os1/ff4q/r8dQoHqWtejpWMtYKl8/m1ydd/nA7oz/+GyFxMHTY3Hw+p54
/oTqWQKlIXCF0dWYXzKci+6dOVG/q5o8TtU4Rqs4663la2eioBWbzsj1YomGsjvf
qWk0qT8xdsAwZvBJ0BmTPrLtOeSENifbFC5QJ/vY8SvMxGU9IuLld9XxF/uWL074
XVQGzG0UFcY51YT/XRe7rlVc83v1eOL9Xcpfa/hyqkUgFmFBI9hkr9u4OrvaAQV9
cBUT93mbBu7FlJ9PhNDhOrmyA8pqU413TZmUrMIAr8a0+BsdjME7tVrt9uSbpBGw
fVAoQ9aSiHLdTJctFx9AyG+xj4Vr5oUWQ7fQMCnEwytik/9GWBJLUynuLa7+8lSn
DF6tycWEGcLlf9DhLEwXDSBJ57JzHdFlTLXTgUmoSwsNA3+3HVpNEa1gIaoQnzrv
Ok9n7xB2dsczw2OePh3+HiutmHB1zfIS1JpIpUOl3Oti/ucu985lmcf4epggI77n
lIaXwOGcUBK79/t4bR1yMJ/lvU9LQS4e9CbKvImn/MSz1MDW7iGaETZJT7ftzEjh
P7FWv1Ve++v67chyYQqgIpyTMtsn9Nif2sKLXHFcBp8mz9z/okSYNTdU1sE6NN+i
A92bYAUooO3AXFuqX3fKj4ZY4aWP2FU1kLu2YVEWLD6cszNqNIXJHMwQkpgQdlkB
itgbR/+CeJIFx0J/SrHcTC4DUf1VrZMq3ygTTR74ldKATIc661hdOJgWvjfmRCIB
zeynl5HI3toYOFFwx7qkabl8QmVMTqygORGGczzBI/JWcJls+KuhQcLed6FVFt67
z5iYrDpw8hQil9xcp9lSi19lj7XvNLVQSjY+b7Vkv2yC0HH4neAE5hXpUrRsLKN7
8/hA6/P3K3EvCHVkMQvesCWN4/g8AKYk7rjvgsUiAVDq2n+TIuMaF1+kuJ0LQWh0
+mDj4q92cOAAJLCzuCwxH9F+7SWAsxkIqMozwcPgGnsHMRNbOTIUmkMZTMah5GS9
jZ2ejZiFkyyiOhu1KKC/hlKJmNXJIUp6HquUo3GkeGw4RRmrM72G4oD2zrE3vsD2
5U/5OXCSD3XcMumc1vrz5Ebm5Kc3gnJ3AFoCDxKlNRWg1OprR7rWP/Kux3JbuPRp
qmYi4o3WfAuVsvZcCsPV17aNs0JsjYsW/j5fgP3aJPMJbll283ZRQHqWyKPOc5mV
u6C13jMZ5aSkJsivzKFuyNNM+AEuei2U2KOLoXSDWpupthWiBhkZSWZxx2JY4aw0
wHSt/mC+oiJv5fDjPuBSYNzLCMSxUg/aDDevTKty0aeKyTPxbYZ+WZbISUIW+Ul5
kdFCIyDzabWquW7F/YEkBbzbNnyoUdj+Kf82SOcTFFVBMcxfw3ELVruNvk15wKDS
H8P3EDC+7OCSMv2bHL7JeUr7bOfd97eBo1XZoE+/R0oKPJ+gbe7sECvjHFNA9mkl
FennMh9JJS/uV4gWT2ERQxrRuMy904OyNolP/XVeBCLvxUVdc7P1EsvInY2gzjd8
aQ2YkTbZybY8yYqD2hKlTPt5Zz9cmZel9WBefXYX3Z6AV5tp2TD8oYd7R7Zm/G33
/7awoZpv/TVMG2XFP0LAkgBkpRby8uwd3Vf82pO1gMjuRlj15TSZ2hXzyanqBki0
s/kxBZIeA43By3UX5QZwObc5vWsOF0KfflqYjhw/iYC9sEgWC+ODxr0Y+IcYDg0m
cmvPN1Nyz3+fNbp8SWSA/NQY5JN7bdNg6FWp4FJJ+Yrb9r2Rkzt+T9QfX/OmkqXu
SXOU2KgXV+bVB2mh5V/T7ygvB9MeOSF6R1WYN4/46hQZJpapo0ULUPhhqxBlyBxU
q6rI1eFHNK+RH7d11zkDZOMN9wG5Q5lc713fRZ0ccJrkDyooOw9HzCF4MsG3H+2K
487FPsTVeH8TFvYj1H7MsLrkqPdNoaaMJ5eqdsIAarWUSmCdvInLJdB3h6MAmdqB
Lj7bm6QQS7AZsV8WZLGIschYC4/FzuJDAmz/LtJndC0aaG0Y6wXg0H/EEqQvZ/il
h3llPn+8GnIACxYOvazogZ4AoHcL/LcmOgaaCkMCr1JkgdiC0LWzxQh7omc9DW1r
O/7OX5BIZ4cldBJifsO8Z3j7VIFmM1Iz29Mj81G4awXL9tvuR2C/fTJFsI/WELwj
35TfCGWFNKXU7tJWWJ7E5TYCiRLONl19kiN5f3IxsE2qkOxIR5VW83L2M3ACgGYY
UQbnxjIeyinjS04zbwWQlSefQI738F4Zm2QOQn7jjtN0I73PWTVFuEIUaWDrJg6M
u+6ioB/p3HS+xi7RlyiqhgLI0vtUovO9LYvhlAF9tYBKA+CaT724Ni1Bb67jtv0u
MFi55YX6TcUV1X74ry3k4S2LEWxkV8dF63DhIdNK1x7WVCeXSotIVvPB+flC3vt7
QnR32mkvOXBC/Ryoqto7TBBPPSwrzQO67juG877jE2V8EJO+7bEL9Va2ctVtplLK
k7Xhnh5tgQswY2T3Cw8hl1ThsS/ekMe59rJwd5bTDOyIlQ6G3qPKiZ8d0zq3WpsX
zPbAVu2SHqWVTL7D33T6FNORks16CYIYp1u7hxA2dk7jQ9+YGFHMzujM0qFsvR+4
n9jXkcL4GEQ4sSgpB+uep/jj0NKMCOXVJUXlhQddV0aVPmxr8vRYNPB/DQnSiFba
9mpkZWEda3ALMJqSHNPd/D+583Ko+gMjRSS3Rb/qPnODlq5FtV7cA9BZKQdUWKue
4Z8lycbhelqNJEOWez/WPcKiGgsXYwA3P5yXQl1RQ8AUSbnf3YZTNlXChLhm2QAR
rUAkD4iNkGqH3CZSBSnF5kIIHXp4HfU6Tg1O8r3DugxTHvnASGFyhcJCroNdVSAW
fHC4PXNNUVGM+E60FLllNM3yXK5XpCGAh3TOMRWvZ9hdJq7e3tzGUEwgaaOwEFak
HNMuith0gKicTUsL04bYV2QXheZcmwaoSljg6LY6+ByBSkS9fSqNcDhSU3jwguuW
EqB0o/SUjlRj6/d6BN7uvY6U1/kzfLbd4QU1Adplbl3/TTDCPIlykSXvbulDZ77d
6teEQ4MY7I0NlAD7MkeKNFESpg5MP8WMA/GE4V9ru8SyPmppFgpGyVmEt+IHOUX+
GWvxRJ6PHRRFwXWk/TZb1SsVYjYvkwoDgkSLuVUg0itrcpZ1wY/0NZR+EcTiF8xx
zNIhJ5+X6ilctV/LgQj36XtBWnSp/fQu4RqjgLdI5cgg291QRTirJP94mgDXnbCP
nLJukO5YJdIBQx3DCN6CrTRPrHoAsQaK/hfDYyoZ+AaNJJiforZL31i0AiRZsDV6
/JeCx/RNSfd9iVxtaxR0aDdTcGtHRCeV17dGBSdYfkcrqjBl8cFK7CNjgWi53TKq
8+CwTy6DadHB2TvXbndB8HEiV5lFHsem3FAp/6HpH5xqrWTmf4DKpbgar66UNWQD
PPfOdi0MBtQL7w1g40O6l/5F2NM+Ilf6UeL3/pCozhkA41GpW274gt1fdY9bNLud
4xyKIefPqNhMpq4nPRCRYA46TdHRXcauZnJIj3gSG0fIwIDQ+5SZBZd+Y0R6uVf7
w+A6GxG1sWtEBC7MSed9siXyXq7IE+Gvaj41iwOcy/fsDOG7s+JllhjmUjC2/Sgx
ZRijlJ+dnnyPV/3zx1MtH4FE+2TjpPa+G/5J99iq0jx8jh18ZPtFqhZodjy4Vv1L
imNmX0/GC7B3ODiEpfKxCnOL0D50xiLHOmPCkqVZsrMnnAEyqLgGJ9qk5e+RGq2V
osOsH/i1E76Mm36I/pQsezDvVvqpzX4mX09yJ1xhbVdwfKxTkzxECbNk5RRacLVk
Yeh/I7Bn76DMKJD9wNdzuHepIC89LDOg1xKEjhefaI5FsCzfP7SYNiOVxN+EL1RH
gJtqCUxByyy2mDsMxSNSRLe2ZYj9SNWUv+qtqbo0Oev/AyZ5O+aVLTaExptMmiJK
`protect END_PROTECTED

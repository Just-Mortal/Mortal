`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spu2Cx5HP7vlDe0Gd8mg3Unx5UNHfz5fLRvGMQKl2PQ9Qj3nJwqc0dtgLj4dISo8
Hq5a9WJa9crjIY0g6BNjfsJiXIGCoEf1RjWWfox8x0Huf/dAwPEnBn7RgXlT5FRy
ShpwVpV5G4pZYwbdAQUukKVIiBx1S0eNNztXlfDdH61NbT6kcYsLK7nmWMguyRu1
BKu6CZib4tBvf7lM02OPJso5NWgEaohvIDdj0YE9goeP1nGRMR71h6dyV1BZXkzf
qK6VG3YAUmzu2b7lD8ZdezpaECuDkMyJI2LwZ3eyqy8oaH1GEsd2SZn52W5ww/9+
rDbE0qA9yU2DUyAk49vfVroS+++Z531m0ejCSOPUeZbfiTtpe2q7+XMymBZM17es
yYgh3ftEsp5Y9J2Ut/8iux+hfjN7o4faSvRfrPzmAm5dVNsPXkMWfkRAFku4fpzW
V7yQm6RhY53vce+xLxNnaW+AlCMibnKiDIlmLyy0A6qn++5XMUv4Yugq5yM331+2
anVjFCauN2IBOJQMW7bDDcueTJjdGnBKp492L7ALtYnuMH2ps6O91IVarNmP+FVj
ab/gcM/VW6n+b6+bLf2wrtjdfnZCa7LAJCFEDqhI0m0eCqyyZj31GvyLo80tXeM8
ctvIjcgTPrlxZ9tXA6Dk8T2Kfj6F19dDJ/EPU/8kWuR/rNIgrnMVi29XeiSIhn7b
c7mSpgi5PZEUF0DvvGC4GZqPteR+JkCIqdPnhlksxLmwWDaBKriwIOP6UKZS0FIA
eS0+Zm2YHGg/fhvXqUg2EjajecwU3FRVvq535HOi0b5kGVKsdtH3MiIZrwQn5lHh
gTdc2r1F3nSzt1EdrE4pDr/HQp80h236hFhVptu0I8GeRYWwYi3Nrbyw46ZtpoIP
pz39UM2HGleirSEqh8WMH8Cfw6ZfX4OP3iquVYbgLRhJ3wfMdHPwcXxSjsBzmPy2
Sm2PSqrfgGzkavmZOKjSPQq61NG4/s83MMZcjGiOnAY=
`protect END_PROTECTED

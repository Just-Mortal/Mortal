`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iU+ST3RkwpHYrbUX1dhhE61Ci5OHPj6o2kYVqk0Vxbhdz/f3iXbJnG+V4llb7s4C
1sr+xOW5GdtDwv7eBo5dSIaLy4SIg5g5ZKMcyb27MT4dhnYDrdutQgSy01hUIuLu
4r8BrTaIZqiTj7PxRwxKu3P963GQTCC9ValbhT/QVfKpgrosU3ZNt9YLEPkLozLS
J1OQ1OOjxBN7aaApsd1N5y4XPz9jgE3xr3ujzV8679bqJWWs6GHEn2md/AqolPPI
/P02lLc6rkoaGnjct3/NoKje/6JmhnUV9CmkWvGjJBlOtfJ3bIqHaG8Y/O7rnbDZ
CdMjSsdc3kebeowrPRTQFoxpXo2NpjzAiol3gBy9S8BUxis7tjuIGspU2MhcRfZc
t38eYZyyDQohUpno0EVqjSHxsXBGoLV6qvv+IqzCTfdepy0Y/UHOoJZnhg2585vd
Ob9vxuSRC+qp/6g9tArrEHiXcnc0hoE4NjmvPu9PTe7QnUlfKiEF2SVwx6sNZ6d0
5BRxGKXr1PoXGu8SJ9W3IxyYBXTkxCkl2DdVUBBClXNLPqPPaUoy+Fj4Q9DNKNLB
AuSQsIzYj/FAZyEHol4SbyZlkElCH/6jvFEhblwIaOZ2/p5lN1c0RriN8tCJOl3C
lKvKrvdY61C+xIVOFhtxN0Ns2Fi+DG6agA9sDY366rFtd13kbX0Y7WgcUHFJGib2
pumXBdkiCD/hwIsvyiS8WIOjcvNYx9g9T/+rB7zkyl0IzIBHELDSo42kZCdQr2OK
zmBxqqs4HDjBvwfvGRB4CA==
`protect END_PROTECTED

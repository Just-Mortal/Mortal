library verilog;
use verilog.vl_types.all;
entity signal_generator_vlg_vec_tst is
end signal_generator_vlg_vec_tst;

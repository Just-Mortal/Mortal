`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cg6i4df7T9ID8DjME3CRvoFxsG2v5fzxUwmZr4va0M3Gd67PoNXZ3i6FIo9Lqet0
KtFAzX7xcBC8wcMkCpzw0RWazW5XLaidMEw0c1VgATelxAigq4PL3y5sjNUojVKp
zuTMrsdpAqN6L7xWrANMPMqKpECgL0JwqHX3qp0wwvdNgLeb8892ekcyCMT+/mhF
qIlp042p8u8XV7zFtoMkfioay/pf2VjSU7sfjrZwe1QswQGbGuivI0Unmx0yUTVQ
YfFsOjsllhjqNTgvsjqeMZKoQlyPQQdxbxIu7f/LjcyNaZCipSr9soDetjjft0cZ
Vs3h3wZ3s7a6QXYOx177OD5+ewwV0EmMSDHzu8iFKAXoxX8vCTugBVSgWeYfLp0e
g5nEQ1RLfPjmalZwf7m9g4HoKZbv9/ANnMigxrzKu7LjxZN/qOrpJjqhGDtkZBT+
/f3MIHgW3Vr5pOTdrPpOCutoo9FYiHRYfQdlxoKU8NXZT2UDsmTPZb0Brtf8BtQo
27yYk8Q6hp6fPaOhBHO+lnkZRQ4I/qlmmKMKD7ksYypU+YDXkMX7ogULO48gC0wi
KhzeQtG4ndffzcGHevS2IZgPZkZUmVbUpsP7HzGghrrUrsWsaMmPfimONIeQnlXD
NUPI4/8chBpKzvrO1ynneNjCete58MViUFKcfinM08o8FofPnBvz8W7B53lOCzNv
fWoq83syWqnFS9dWoHbl5WS+ZLnRqu80vxIwFwqjhCXxIhTzKEnZZDDv5NVZibxl
Tl2oupWXtmeE+QV3nS+eJw==
`protect END_PROTECTED

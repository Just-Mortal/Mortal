`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7W10gxhAyN9ehNwCmsB1MsSSytbLYgpI5xgGGVQvJhcvthbvNIdic5Wlz7qrEDS
xYSpSaW0J6DDo9Ho7KlNGIcFMYwAI04M0cPQAKay4JnnMmBsh8ur0/rwLJ/Ydz4n
PHKw6eCuELERbEkm7ZPu/fZbOaPURNuYltFOKHzNXce4ziCazWJgEiCUC4Ff5Bkf
oRxEwiD2ZGKNSzlJtIAyuJLE9UHTUByP8iDtKYNKoDlh67Tkdpy2DggNxZLcetGx
+MhtzDT6QwQvcb9qNnc/0LaWodJv7SPgbJcWBClCdRT/xEeo7Pso+7e+0ZNKmIt2
3VNJiu9CmjG5bsj47z85X30YnvnhQIq+RlyayhxqvH2hH2h3i50nRc7/Sv+gnmy6
ZlJw3ip9MelLSAIi1X3uf4G62hkr2TpD8BaRu3ldlnJwmeu6riER94r6UghLCiYP
wfrHRgqZn+hJQZfYulPQ/fXYrFx0k+rfvISoo8UdJCmi+usEuNmslM+O6ev6GtPO
F7HiKiN0wZFp+33pqi7/sVb13jjoprJnEKso15j+w4fP7d8v/kQQNguat9btd8Jx
YevtJts5NlumPnes4yeCX4rHD2ctvkyeU7hcvRmGxixbL8729r7SU6eLmEiuFSmR
IFhDAfF6mjkdcxeDSKPlpZ1ygHYH0hSW5BuC3a41yZGvXgk9RCEsJqfmx/utlG33
outiS9AlYW0BOOWl9AisFrFaTtVDXNThxj4k3AWmDHtawJ0DU75QaTchQNIX8MFt
YXv1am/ej5srmc2cogmbyMbQotfcULko6bmi4m23TSI=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/B9lk+fqvN5sebecsgEWA4IcoIFe6LKlpy575BOGLugsZzIQkRBOs2UuoyBlncz
YRyO3du7D7URYB2kBxslmhi/Ad11ibY3DWpbfPafCDj4OQn1Rk7xTzpeWMW4M52w
XZfbrInyA7jhTVLmGA8MObSw0+MgYAvmbZfF6bGtEvJLecYt/YYPhMCDgqLRlOZW
unLw+LYPG0ptWsfLHwstPjDvo4CgKJz9sLuT4XmunK9tVcnAO4d14YEiIyUB+VuO
qJzQtHHjvycH+yAX/TpNbo8BWS8DWQfMBwAzENpJDI+S+PE93Xe7QzgGYufn5hcU
K3kTTY0IeG9W8CmctouPrSQ4G43+oRkb6wnkZblqkcsElPGphbz+tBQSZpOonYMT
euzyXarVDtoZ2XDd/gAfwLvv1jPA8rE1kDu0U/jSCkclcjihf+LT4HznorFoerF6
z/n5nAQ47f/1Lk6XpKNo55i9IIbE+g9Q+6ipGjGK4qKsus/2uID+PeR5CaK7Wd9L
HGuDA3wtwI06irrXbAsuUFWIv0Ss2DsQCqR3Hv3syoru8D3uIgPv1ApU3FjMUb2o
eIO7je4s341osEEDSn9NUY6yV2hfyPTUCwptJ2qt6G+GbWqNUkX+rMUX0RrV7Aqp
iPODu3FyGt/I3wEQoN/5TZ8NNUiOyXls2747encsYYEr+kiNlkUxNqKC9NNN3oIF
l4OMiXMbCcBlgHbAgbsst68kk8BkYsXhy+2K58p7HqAEBVbybKEJLD8w3NNI/zUd
zNWo8qJV6lABDVZLxgx1xprZ0IoBxcoLCOmFKWZWQ5OHnlz7NQF1Y2aqZx91sX8H
ObesAf7XtAAuFci+Qikhfme/LyszesUxEnqSFmsYuG5ai5nECN+HoPzHRkxLN7oU
LmC6Ix6uyvSMRQikkIOQq0s3WtgM8rXSR/wMdbISHIZ6lSOXBRSxFpxbvEhxCTHy
S/RPBllSqdR5rdLgqyHWNqPF3Q5umocJOPcBrTfXHzSelfk0qaU1RQFTRxRG6gTi
izHap49URbPBVdAFmKTVP9AOjStFJMYKD9DYlMVBIczD1fOe6icLlw8gPMOg5wTX
W+pin4glWHgt6g6Ul5wmY8T3NDQPdWO5TZZ8NYy2RE/7ooaGAUhFfVwNWAp0dgjB
tz9tTjr1UBpw7/2XphoT+gEKLbs9qkupiJR660c04HrW3y5aww8ZWQmTW+1gHrTi
k9NBrR0mzOki7neEIhDV1YFmdiGnMH8JxqrNFtV+3EZvnNE3ov8zri/JqfxXhDgd
RZz36w560SWGN12b+BbqOyXqYI2CwsG4b+NmGJp+UrOnfiQOF8JhrNWr9yGDMgrF
QAO3s6qWAM4GtHAv2AvH5f2GdrSGsAdvKUNPt/oUcP4BBbM0awcchzo+8uY4eZU8
YWaC1vbCVfxkVTDPfs3z9tAUmieziG/N6bsAY9Gw7DmWD77Q86MpEl2pqS+owCBa
bBOFsHD7drPKI2EBTGRuQ+taqdTUGeRiO0XhoZlCODzocs+Od+eXzjkrQU46gqGX
y5phr5YRwP8su72/blo1tJzDqdnx8dq4xYImqnnSuDplB7qIpV/kvuFHX2Ql+vnQ
ZB5qOJIjl89mBovMbr6LXK2dh7euYoCLv1D6sC4vOK49Y2ai2N+bEpdCznDxo/oY
JBAMRYuiv0BEEVmo+mvTdQHyzocEgtFN8IY/4N1PJdNOS7DtlPmvpNpVPQAmymVz
nLCtNnW4Z5RjFPN8woB7qoH1AhqkG3ZRbmZuUPtrrs/yGOMiDr29UYnSOIz3aPxD
fTwVsAor9DqZjwrZmO0PaZmDejjG/K0nzBwTB5sZO78ilUhlUWzwRcxO64mp9SRW
dkmfm/pY05bNkEJdh4KbyuHcMbw96bh5Rh5IBRXkVUZq99xl5MQq2RZuHdIEXjc4
bg8lLPCa7ShrRyVhyazcsjV7L1i0phFX+MdPyJi4VFcL24CyQMYd0O7bFSG52u4x
i92I8ttgzD05KVx7Qrb1ntF/Cqt0N3Dmgc6eBWq05fXRxvW41rsr4ABwGjrdaEYz
rHBKdoOvd0yRh7PaOEEVt6+9JusCXYMlOJNLfoc5BfHb28hnMxhh0Xfo3i4H/Xxt
flgl36LUvrk7UHEbtiMTD5vcp50OrUCwmFo0A/8VkPD2CfrhH58WEuDh8JNncPjG
72nb0r5CwFVa0prpOAYaJeHBv7a5gWTzhwS8S7LwNLgNbKum/r+52023P6vEe+an
4PJO7ZbQTfjzDnqsodaDiNroCPA/M5KejpaTTBploQAchsEzdX9PRU8MiuK5QP7z
1AOzpHwGuboRZOEHsVKieP23VL1jcPgE0YPgqGowFFF6ZrjV7EKgCbVFYDJUL73y
DDr2v6gJXxK2HcW7I5L8XQ2Ps097JxrY0VrmmMewmQgVJOqQk7XYG4scYcyMdqWd
SzMZxzpHfSPVsk+dhD0fNh6TFq8DyiA4a+mF5HDoXUViYBGG3f2Hsil0II9bkmDY
e7R/rb3jRSW+kLauLhSR8hdn3H6dry2EZh3q2YPL62MJxdcUjfSDW/PL3/34zO9J
trOCS0qyuT1+QgZtXti0FSRPg0e6/XOnD7zbD23l/JSKA9ecHsGZIrTHKAEn0h+/
YcKW6N+Wf8sQx/F0uCPw0tWk3GUkqBqIjCpw1HUz+r2hDNi08RYGXuIQSOFanP8F
TYt6x/UGLgtBo/H5P43cwEY1nIePrds2zBjeH0VKCJ5QCcyhuFSx0jEw+5coXW4O
g3o6W2jdzXd0h5pQnCN492jNgtvWXjSrVi7K0pVHls8V59D0uKkihIh93MO86F9I
nnFzZ5Ig6PM7RQUqgbTjuqIq4ncex7YYixuw3qZRVOLvEd73mva3RZ9nCpe5FsYt
xqvxH777X/mLh4TQhU60ZCPehr1rMZL+jD8P9rEVFTdYUzCX8Td3yDx1bryDxEiW
wRdvNGATF2ORmpcjK6XXtCVmUbkZM/B6l97U1bm0ck2CyI4jUvRCNPXqKNshSbW9
YMsh9Fs8+HdUG4vQznOfiVVzLgfEF8SiKgYe1MdIxvzGorSksx94d7sNC7/MG6F5
+ZhT1bC07vMqb0gISh1we+rcbesv2/lXHQ2ra9uoKrKQcC/TtgK/MEP+kxdWDvV/
GnLRWYKvMTISCOFVdKmQCdMr3hjZMtEX6KoVwGXMdFEr6Chf/vWap++5qXeikLMZ
EIJQoB5IJOuzwAAlujiTgYmQgaGWi1q9XlS6rEEo8aS7C2Xi+JXiYpKoVH78lnHZ
njd+JCILfZwo7mePU4YM6+cGB2FPQAxoQBpXlXapfA5yoIlFkSTMmE/haI//bSi4
thpZCnyJstALHa4RROiAKvFmswYCauK8zneqzCKvzzj3pr5aPThO1WLuoPDRXKLP
eJBge3UpfMUATRy+DPWXDb+b35AbVoDi6BTEYxNaAfg2SLHmZldTV8j6FR/IG1l/
t9hjs2IMzIc2+1jd+u/nyzB49LUEWr63FgqSsqKjiIAX/m/+GQgvMGy7sUdrAMFF
XxzFRwZ9pv0lySf8OWi5huBP4hTo0vJKFshcKgzB39lR30IErz9daMsEgaqOSaKW
ZxkVcBZ42Ik6oRcKOAyMI24SlVvnUzoTHcItnMiBtfUjCYJ8b8ca2nOMRMbYHRPA
W87tnWX3oANag9Z/AKErtaHPylU0ItCPidfl7nY619KW/LaSubNfM6d11RXz7U+l
Xr1xQePgPPTCp2PwPx1BrkjzriAWE4a1zB+Fxdxz+m4JkxZa/y5J1GTFT39vs9jL
LrELIm9SpKfplBvs1JO6yKPocvvisbaUw7YMd1Bw/K0UjpwDXOWuscOatij9YaIv
gJwLRUXvpywADpmnI8xLankpLBGUwbub31JdjbsKVLdvCE2a3315wAH+XAaHgcIG
85jEy0Z9MlDpO7dCALAavOpMfYuafiwK9H+GiQLkCy/q096PJ7sxGEpGH6oX9B9Y
RxBy0iXAW80fnUT8q3c9yi59WsCFEcz2Kg48MK7B5o3Zb8hN5+F+hquniUTB9KvJ
PPATZzy323Ajv91bPFAzolanxw/KvEfqJ76RSvADTCXT+mwF1U2TpljbkliQ/6jg
N9lpQF5KgIe8WPyKQu4ZX9cRnNyrD0K52Uk8U6yj+D3rW/tdBgBOOm+3W2Dg7Vge
rZj5EqB40vz93MvDwPnOxnEWvs+Olb/8+EATRghyJc/a4luZK7q9bIYG/NPrack2
WgiYVCAD3fufQQKwNqMsDu8ofbJasjLtUVKgRi+MqiRJ8QPuFfsnfPQ/cHlCZ2lf
/zponDgIG1q0hewo9u0sG7sTagVnuWkuzfAEofso+GrSjFcfx2ssW077UDC0onNn
G9KKez3iDGypvCKhPFmq2g57tLPPfM+CYheyjfSmczyD7nt3uMsEH6Fy/iEWCMLI
osXp1wzXJl0ZKsYtgy5io6EaBeEStq6PKU3ZT9uiqxnyZiWeB4WZdCXsj+Lu41/t
HwPbvcHC8rV1evjwwIJEwyFv17uzlXVHKugU+8GyWbi2SswT9MxRFJKrn4JHBz/9
nGOPJXXnhLpC1qW5+oYYq+ETfHKjRiZv6SQ7N9gDdDAz76hXsi/Zsl+IH5khmDPF
`protect END_PROTECTED

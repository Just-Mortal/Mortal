`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyo/8kP3oVt4cztKiIBRSaGHtnKI3fkLolneTulxaubAR1BAtB234Epu+yr4fTm5
+ELrQej5tYfU2dwPiYGFXrEQz5lLt1FykRXpXsSIl944Gu5/Q1bRrsNyeKK4CY5y
COT/aOCy6XjB+kTAgEzXgrn23UEUuFQv9KYE2ALcZ3UYMS8sdzEk4ZAAu+3m3t6D
qVI2qtIh1pGGDai4QKVcH3v75iqtdPRbcY8ZT5r9JRftEL6n1Fi/6NQ9AVD5OBOR
zSx0aXRLVr0uklGUlhdeymog9+OUR1N9GUDPlUF9kqS2/ftd8ASA2b8T9WFBNE6K
eOvFoC0elOgTV+vzT8IMPgMI/yLSxFNr8sAA8K7FNiSgG8SzJeWWp53mGn2qdkgr
tAxO7DSkeujuMEW+NviOrzbDhaeVcJ/OL7LOsvc3XKPGhm+juJhmozVONUTJf+2z
7n3H6DFmXfDkIREVrMLaU6xKRmNC8oFD0fQjHu6FvRlitiRpONnaKlqRgkos2dyc
2MozNfqnDXqUoEoHN1hfQ1Lo0kq1lWVQ4rcFFZKFPjYzC7SX4ftsrJ67TKAujzWU
fCC1X8jCLcd3Wk5IShiR8cDPKk9DJKw+phoyWHgTcdzWTT3xym65dIDktUVp8m/z
P+dIg1SBO7bIvzoJJ2ysYQZcI+QWCG43g9S+J1ncdqwjx75dXFpQAux73uUorron
hIoTKVgVqXP12xyxDb9LiejdX37v8tjtAmWCNVnOBgZ+V1YUa9CNYOvzxB92aPE+
iMB1/vifMckFw4mBu+E2aKbh1AMuPqi6fUJ/+8VwFxJYcuccCXWbC3pF2+XvSBo9
t5Pk8dhT5jeWooVxCVgKUn7IhvjxBz78PjpaRkdBEuCkKfSnBKNmvC4rp3+Td5cw
qDNpJBtsymGkbo4Pjf/n3rp/5sxIei2d21mhbsEB0cE85lEkexUp1Ey3ugfHCkB4
neZ+PF0TcNkTez0ki300Xwy2O8Hz9DtHQd/o8rBvHI0=
`protect END_PROTECTED

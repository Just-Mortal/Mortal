`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5t2q4PvhWUp9ri8uZX26tVfG3X+kgE97RMzoEg9NbhgW+6XlGGanb8y1F4fZ9p9
KrNMMgL9S2MWVN0Zppd//XT5jN3yCgW2XpY+PR98+05qw2I+ID/+RuSSc81cbYdP
f3ln6RE7arOilHkcIqQnPmrNc1pfVF38DxiyGPxPNNJ8eLCxcLWawdJyjCEN10Cv
crLWY8HrAwBrVYNLwjlhLdJz3fFt+/of4pltVj46Cldpl70LnzEXj0nTMEbgQRpO
VW4ICvxI6S8aeILDhtwIqUpo8PeH6dduVffAL5DzbBvt+1kG3rZDnxnXe5Htfg4q
WbgffpnVzAj8uZtky66hqRQPxxVlOjcdRwmk3qZdWnJy4EpHvNpOz0lpvdGnWfWg
U7X+pTUn94FW2/9Mq2Y3gwSKsd6pRcj+S4meWrlQoLgsx6SZBQrJbGIabzWZCaxG
wSGBN+4p4A+hnEENcPZtMAUySt7npXuSE31KFBTTpRS/xs1MdnNoASRsBrGOAM8+
AJNUSv+QaZkwzC30SIogap0Z6M06n1ZSn3XFRUGc+2eswmGXcciMMVbcGEZz9xQU
KXrwsjigx1ctUP13dl8YL4ANU33QB7AUpxjqGUgYtgzCtlNqajDmaAS1Kljmet61
oyimw2qiyG1p0iGlm/4Kq+3ml0y7ldSMyp+87OTkbWwEVYnfZkdez8LEWt9KSXxS
uWNVtl3o4Kcbj1tLk2kvfshDObUAqequOz8Vvc2A63vse8oQ/HCq0mg2Fw3Ino+Q
BK/9aEU+dCcECyELcxSIUi5VEwZG27jXM2Mnc8YGXaHABeCMIU/ozsYB4Du/Vu9v
6fnGAlLG2oZkqT58azzIQ8nXdJ3V+iGATrVaO/56ArmIYAtWSCYoLHUnWbkCDsSJ
LmtnAVJnOcovzqSd5C4ggjXBmVn/R975BJT5rB0Cy+movklgt0E6jgpeBzDNW6QJ
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFn1u9Vd6Dl0DQXlvb/cIuYI77Rp64Pwg/zEHwmH3R0BYz5GQ+eV5iJjbcgK5un3
MHJ1aKg/a2kd1kk93o7LngnJWVtTsCXS38yFcpwR25YnLvZuQ7Nn+X3qe4lwsn7S
dq3I3VVmtRChEN/RcllOlvK/Id83EJtBvungtZtOM0TN7cSY/zZkNcDYTzDncIWb
PtzewGJs5aEWn/QSWB385mD3I+Q0XjUYKQPt2/2X5Hm1PGXkxQ/5Es71oKA/8LGb
qZpvgnAsV/BUg0Q+dGAb3FFCNHp/pW4WqJYL6dafZXcbzaQPJYN1UbdQUXG50jEP
PMgVytgWMmMm5t0egVKrdRB6PDhak/WritGNWgaUxyaWMwIN1gMzF1YEByDfvbnE
HPTwIzJYa+/p5UgtRjuVoulcBkHqkmEblW0ZQdFWvW1/MzeSVjnEvOFLQH+zY9lq
6Nah16bhqrrbC0RMGSz3qMSva+nfyDOiqaqyyp5MuL2l/Xoz38DnQ63e/+whnnZV
M/AbU5QjK9NsvkXGehZxQFKFWeHbSozyvBhWYyCahdDak38X1EaNWgiE7mv5ciSB
/ZicAtsoyfEmohLfLvEWWIWobfgn51HKJBbUM1iqD6EUA5B6pytfq/npYJ202/jF
4YoZDH/yQaZxcvOyuu9q69WFfv3Z06Sp8V0QGRMKF7LDouJEzEylgfz2Tf5W4ZsX
CZDVtp5oWKQSIcJIAuXzno/8mjpOOUcsAlyF2QNuZopkBrjvReFrYNwaaALgZn/E
9QoIuFFdzHJ00C+n6zeUHSVXJzxlGlvAi6zCh+MLl9pPRyQ71zsSE9/medTcNWva
GLqqOL4FU2aWiTl+6ADyi6yJ/Hz379qqYGv2v+UKXMe96nyeAOhoQMj1uqamxam2
1Fj5zXSuTcsNlcjKIlSNyrCGkIWmDNbeb1b+svWvT9xElrNVArQs/uURIV1mKh+8
rYagGzNX0t/aG52AWVuGO1C+9b3Yq6Tro/IcmuwnqhOyMF2yvYwodoDhHTHCXIPX
GmCCaACUDspwsybZOuNWuu2yB3t+eqODVW/htwIQ5aCnmtNQonjdRo6OaDOIJGRq
IznFfNcrtmfJcqykTgJvZs4EjL0nmPaIwgUVExf+S5myahBLpmPJQkOAqYzx34Qx
A5wQ4UuIvaqAlzTsEQ8WjKk8dbydyIt8UfrTfpt+ikZGCo3//DFeVOO4jqJ+RmSF
iPnQsv9eSp2Om0ZEr78x9wL6V6b3dT9L3UJJJgKDBUjBlH4vyWDqBB51MFwSgrkm
oKfMcfh6n9xkbVYt+IDExArNb4Eqb05jVTQZhEvgQ1xJK9k9YTAoCteFvXf9R1h2
l7NplFx3DfF3YAEpbpKRB3keE07Y8Wr2azb/woBMwK+0MtNl4pR55lwSXhS/ElVo
uzTo5jNy8ErfbqV0QgSPTMOXhcvfyDPwZuz9H6r1xlksTEilEFSkB9gPni4rVkCT
MeMpvGp/M/p7BbZHkZTWxWeBEuV5K+lbMNrCd0XpsQBLNss8T/a1J5ywsDsmDAGK
OrI/bmKjKqp1HJXwInylny1nzKHCuE/zUQYTO7rf0DbiJgP4BjNUVIEFOo5/RfLD
SYLa9PF7JuPcQJAZ1goTS8zIsWOLBuYjv7pCs4Wa72nB28zUa4cvPvKIWR2l4L/t
LVxU/FA5m5P4902sD2YSIuCDJgmCTdMBfyLv/iDO3GwA2iBR4dFcAc/lrzE03aBa
obK0Vn/jK5rKHPuQlUHY8bxA0ZyPRFDYEp0dvnPSkibArwoq9lVl6vxFOM0Vv531
qnFti2IIAqMOjiTZBIedqHzo4eku1FKg8UW/6/3ZZC2GvO2ciEFHw3+nGbn2kGyk
gcwkJ7UZ7/+NVlU9pX+PJ58dl2EFTTaFIPd8j/NRWnmwuaUSOteRCtb/7iac+SQ7
Zxpf51ffCdJWFZmlUmopTFnXYOtVvKaY/FjdHIi8OUHHo3jXVXVKkgIhpnvWNOmA
ORtnnTDXfSeovZ4fOgqNAbYvkP8QVgsiZhSAyESa/2YsvtTj7Hi90wQavp+w7bmu
x0NbpmeoX6dwMS+/pNEjGANrMyocg0PMK9GIjApSDDfXHTRmESHs6zF5COBd8TU8
UCfBCbe1mERRQbFM/PjcQgxsqKJqvar1UDxfVZsluNhjKILgfnaw6DsL3uqBfkpl
+ZMWy7k+m7iCbQt8w3inYC8eozNwaKqa5qoZj2l1cpZasfwtP6CscayxaykBEBk3
FFJ1a0LwOHzEof8B4JY/iGkUnOs/ByPC3cdgks1qr0y0GNQDujFzN9e9FcQPNiQr
Pqmg616C3t9i0juVo5IvNNm4bc8c3aUpBeTbVgDKSUG8TN3aul1F+BrOsWO2AciP
RzzXS3or4xE9Ks7YcarX6AS7ySMfEYtxcAnO/daln6mx1Gop2FxErKb/FO2XV0xJ
0OuLubX22D7MZX+7JtA0ZLaeynDs5ZCDUZdsX2SI1rzHLtjJMIkckNjmhpoV0VPM
CR1VyNRIouCZYfhLC+YnXJGKqEfu+RlI3q3aDDxAR3e5IGzJLqfkYleybBWS3oTz
FFMOtz7/zxfbm6Io1kGrGkIctA/OOywGFfaX8u1pkhX4gwra8kWwxeSZ1pDF88cA
xdOH/n7DAWKeqGT7CYAlrWF8a7MUBhC0AKKCiGPOB81SqDD2JG4OK0n6Zsr1R5Iu
crmuv01oJFbIDjjVtY7jCFwJy0lRCk6V+55tVcf1zkcOE2/ZcVdcWY23XS7QVgJY
UIrV7iDlZbXMaZ8rYX0/y38iXpzWxUwFHl6RNZECxmlHSZ8VdENRiSu/gdq1Mcfs
3ueik5nSGtcKoKy+KF6U7xqanwbE9EIv4DcH/bXHFGOYfdHzLvEqJyaWXQlZL9Qr
AkBrj0fDiiwvrpTfPjKvAtov09Yqa8+qk5l7d8pBo16rB1fW2zpVymmEITAJxIqZ
GykmvUZ56vzz8BSL7j63v5tkmLVsS9PPnONvtj7QrcTakiOaq6zt5A5pCUOm1UML
YjMdzlsuHWgn1walsQoGT/E3b1ox2OCU1r79rZbIKVAIC0EqSmm/SZHXyg7EyJT8
79YMgjihG5HL4IHrOdlyV3EJhQ6l+saWnfxY+mBSTgbpHWeX4HfFEiwHD164+WQk
4S11LM3Dms0R5qFnL9HJWdW3E828pxnZRRTUCjb19rmsyEmWAgTk6KKz0FIaxaUf
/jtUm4LbLa7oX1Nw9flBjEIRfkQ2jkd++bmu4DKjWGHS147H4WcY/BIUSSxDyljH
amGOp1idAKX5C5saO9ySPQpauEcFFHVUy7HYS5lKbifcROI5Pw2yCPAIHLgExmqr
B8nwTn7KIHGf1rF2/2N/0sdvkESfTWqtdU2MfmsHNMObcOJ3LKDsvblDlFk4bH3y
xBFvDOFkBvS4+mOvWaG9RAStf14zUGQ22lCE1OhYeNhTrW0CoVMCXfwpYYU3i0Uy
i5awJHvarw9A1986f2RN8ZAtRp7lWNl5VTFTCZdLTZj/S5F92ewKSBoeitXdQqnG
5zorq30/p2pkdj6yu6tA47XZ/HO4FEDLZU6wLeL6RSEQX6qLB+/TZE6tnKAwGWQ0
YOQAxTSsfndTpLPVjIM/95QI0Mlo98CLj4MFGMJbNchwthNubo6ljSGiCZcPQWHP
s2psD6mnErvXUq05cfiAw3o6DbckILBUpPUfIbGj4hsEgojWqCa5JUdbq3q4gIaA
VCHh+IKYGobjlK9P59UxVlEBxxVElyzjg7BK8tKEMu/ZHRrqGQ7inKwQrby1zsKZ
GGXaKhG2vW+tjRIoRQNSbJzjAQ/LueBorCd5yPNuaI50mX3NH6vsTqJiDJbLwqoI
HwAvdDbToPpMJM53CrwjQK8w6gl0bbaUJWSbOtynqw74pVQnAJw/SrLSIg9ANXtO
5Migy/946Msstne73RUGWOUmYUyJ6wszZ7sq+INfYlqwna7XvirlA1qXJPPLy8gp
V/j/mv2dCREMInV1eD14YO7mI9Rp/haUbZUKaWruEL8rtgiMD09qi6amHzOWJ1fB
hVMK2bPKZSiMcrVGiIjuoLifP7HkuN+c7a/cTmE0QVV3tcMJ+rzMD560vzSUKxee
fhQjAelMreMnExBHzbraN1vdcNx9neXOWGVbcAajYdDHRz3b3+sw0tuGXjP+afJA
aeGLL7W6TFd9qXXgxsY/fko+Q0dg5YbnPPKlj9GHkq018TzZtddBIcBlpVFvmoYg
+40ZTKoXkYzD4KbT35DpEBxpiGX7MNeOxJB6LBo6HEiAOIR9XXIm8ujJJ95iEgu5
8d1EZKElYE9BsjoTGRmScas40q8nOPXoi9mkhHBACSxktimFrMre/v1Sc2zx+lyr
GydeCRuFbNzPfnSgvbmtd11A4W67rTqiBeDtpMVT3Zb4r9i+4mRj9HJxMMKG9iDm
J37xzq3PuO0OgHotiUPal8u4U+wa6PCoJM20QjtPdqiAMN0/XpyqHKzc+R32FPq1
FRM3goDHnBNSB/4KFOfRBRPZdVIA7QO3/SG2Me6sSFEgxONMrMaRW4NwVPscrnlB
uQ0shSAZFudSHhZIr+BpZGThmDq0D8dmos2BUlEAFdxVG/Wb5jn3cwZp2PAb9lEb
yZaUd7MTuaWHSTwsNzIqUFjjKXnH8Y3LzAxNObCs1zjSgoq+RNQ/a6UDNDAFJ4el
N4SvmH2E3INV5yFcBCJSe8t/HtPnnAq8wWWqe3gIazWaj2Yt5MRCC04aJLjt1/ev
CFrXToIjj3ZW+uueNIvVXHRQfw+NFw97HBwWbR3VJG+/+gHFqJzZfy/BNVWCVUq2
EQGWqhAeWC99z9Aoa3EAktdAYe0jENgJksUkwjCZ/hyk4UL8AubOQ5YQK2X7exrc
HW6tVNYVotuCzGpE8RAUFB4rES3kWsqVjZA++uIcLby6NsdBUbN/oxpON6lV2V6Y
/Nr9F1NPupKs9PdTOOMeseW3tazN4xSF5c5sfAnaklpUKm91Sv2wN7o9tnc2tdzu
kK4pC9i1JYe7ItaDvMR4WiUhDhc4sUSCXpvOCRGvfsDFh7nYl+7dlXjXJ7Fsv/d8
tLTGC9k43jIIKN5Haqw+W0RpzjSftGPB5L+fPF01GreqsBT0sjPy7iYcwNF0tpwQ
S29YatIJ6aVlpeHbcKj/ndXUMf8sY4e87SANV4jM7YlWC3YEt9wkHSIUxLJbj89B
UtcL42KzmVNZvJnYDtLhxjuw2bvH89DBJxQDD6rxkWPe7Es73ejbHgIEqJbLe4/p
J4WOMkqw7sH+LkH0tR8rn53ftFh9q+PC6+RF1gg4KrVoQ/9rzVChy8K9Ox+dcMUg
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJDAvf5Z0yI3JdC6yOtEmXGb903ge664KbgG0MdlfRp95o6cWHeJVv5hZa8kzenn
FAhbakJ5OyuNGvEZnIU/Xqua6ImWJ9NbdJaGp1zwseS4X1gwagEdWW5VSDa9wu0K
lAgiYZQghtr7GSZKd2q7fCilQw7+tOY9mPrASP/bi7ewcXThHnOhqhfkyL2BsRVu
GTI3q5RqETj2i72ld/x6zUIxqCc39DsbENlbiev6RZ55BnVQsSLQUKiFHpnGvBWj
M1tAeuovfz2/pwVOaa+jOFWB14LTPK4jMwvWN7pWUua2tSYwD55G7XRYrifwkEBr
qiJOhs8rn4HXjuRdi76Sk22gMnSJMC/KQQtVqviZlsmP5jIYm85n/kocnctT8J8q
PCoNYdxwjEFqbmgVBUua4Ny2uIcKCNNDt7MU2IAtxh5CuLiLU5li1qM9rgKeL+dY
pzcA7aw4Ea9CwbdSHCCStHr5Hs39khWhOhaaEWGNtuOk7hPwVYlgIWMsc7UCo6iw
l0fuwx46FBm2m8vJa7viK8XtpwUfPGMAKgXO1mnZ+lT06HaM+RotcOzSo3obqDuS
+Fv9EJ9v2BEaT2Aj1gIoHF9/qtxjCpHSepR1tjuJZAZHUODo/M9t8mtPR5DEldmY
twjv4CCRN7xmgO2meUe7rWUjmsLWffP7tpUmsMAvpCKmINZtqDXMVNhQFjRduQBG
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wTObFH3Je+9I+pzOFpfe3f4sx9kqrY8V1Jdzs3CIf5Q+B7XSmCBnfX6BBT+HBHxp
/rBLuU2VpvSgqxJHuAPAbt7cmE2pYbJi1qkUzfZ785dh9EXxnodZOb5KkGf1iuJO
/DHune/XhLfpjoXn6tEzva5JPo1KrrvOn33rh6byABwVQB1opWv0rqC/tE74RJFP
hAvJf6C+JkxZ7e740yueU++LgR6rN0eb9dYBNDJrB4nrkmYBFFTnPMxeNfTPp752
UoM+lqhvYlDuerOtIpRzNhssNS9+JDweA5K5gpc4BqUrPI9IPmVr29EuC1rztEP7
H6LldvY67fclja8ibuHK3Ps2g2C2jzwHP6mBazllLYDl81VHPVHFFKSt0SXm0wVI
5I9L1HHITnEtRL3x0MqBrxRwv4IooAz3rhhS32fU8TDgzusTpNmebleCAx+GEzmj
4abshlfMwaViGx18KYIsnV1ZhvMgofKWKKusKMCNs0u85kts2D4qinnYf5IrcEZx
ZBiNM5Njtx5gXHW/52hc/fd0xE/hSyE+MhCx1oUjQYcvUPVmQjjHcFh0rhJEvAmR
ArH/rnuccyU2gJ9SvgG3WFtRXu6T0lxvpUjglbynyOObm3pjwH2LJQ1px3++n0r8
MJInMnouzfz7kWVIR33/n+Ar1D+7Ykbv7+zTyvdUvhCSHZ3mlas4OLrTd9EUCLLh
7WgY8c/I4FGzCo8158r1c9P4BUBbR/kfboI57JIq9ie4nHiBKTCsvfrt4S2KItWl
gsfI5Emk0Cd397c9qjM2zme1DKix/k30wOy26OSYGf4405/7F7ACP8EpIRDjwVsc
rgPyudq0XFf6M7xJqzn33g/vzNmVgcA9+wvj4untt5h/yVzi7MNbgTT2bZ51AvL2
wqz+/pXGQDk8tS1qLns1ad/eleuDdifZa4gjkS2MqISWTg5ipRjog+HafSWkB2we
TMPHaX89PhbiwNSRpb17IiRVmybn7v8qLsxGm3Zb4IqPF1ggUSfZV6KLjraVxHAR
ALMfN9UaeYgvEzwRus4Vigr3nhUDZUXnJAuBdOjkSnS0hkUF9CuZrCDzrfU+Pe63
uK2+n0AWLaXXRkty7Cyz8C//VVOTpE5jvyo5+373OIdoQvH6p6phcwmuTjJwIEvn
ktfm/B5gPW8J1iNwnTNIkZrC9TfKBOnhAkZFpKyO6wAXOOLGtnc4QZiRgacqsgfS
Pe+/4eO9m+2+IeLUQYVssSWbNALCuoTdRg+g+9TzKBwz5fixVLOTpPvyrlDTO/M+
zOsGaDvSSzKapAL+TJUMbbYT0im+sY5kymMaIqe2/R7dNJv+zSU1oFYkjiuwf1nA
B8EzDC9ByFIiki6qIhoKUmigVlEFla+Efd52H7Ym7lxDJwu7jjcBWnHKohAxqS2A
y56gTotXIQorXCGWkhWgyeIMINzDw1FspZsf2jqmFnb+VBFFH9+YQvUJmbp+4x/Q
HrZJaAuCl9/n9DwTpAm9z6Ah1UKK6sKhtOBxQJK1gAnhJn81VcfWIF1OUa5kKYEr
8/HPJ8wZiEp8BS2zS0ibo1aCMNS9aaHhZ1E4jYrkVpGuSfkEc9K8Dk9V7HqYAhep
bk2bfQLb6szKQehRUaIjhLsyKRCVPzojUKO3PpF0QgV+7SubYfcYQg/jxMERMQaP
VWwIY0bNM/gYdYVCZe6UJWEmu8rnizBUscR+kcgoNkQvsnaiLy4zFF5EINUIIzoy
PlqRepU/l6oJkGVhf6Ah0dLI5gMWfoJ8ZI0lnKnWhoj8ivXzQRLW5cvxR+x8617O
X3EFl4h8sYigMAUOYmmwqY+FzJYHvBbeurtRU11dGdzi4FJ8zOj+BZRAZApeXnJR
FJs+tYQAJq6Ehm72efRNegRNH70HuhI8piF67Hoo4Mm9/nAhbZjio/Z/dofDgdrg
Q/ZK4e7E16RZlk3iFBR6pY5tf5ixk9UlQQg0y/oYZQ9KKO1JCJEFyDcLMACHlY3o
zsspN6NyL/9mx8Vz61qWfAD3LI1X2A8kghc+3hYku/TBblo5AcOzy/0YzzQWnGrJ
58JxdC+PRBHc5z9ZE2zd17JxSV4vSrzauByL0LhzKPgw4n8Bf97iCDi69WYV0quS
WlvR/xsH6KtJzq/41ABoZzlUtzFX/NDZbFL9yBcnnSYNNR5am3cvc3MxylLmcyI9
KpwBT0mSRXPXOCWfb8oxASNNpwfaWaXeJDSGopF164EwxjHzoKUauwffiyNhNiwA
jyyRra57lm7tw/JLDNuBpUpi2wMGumJPw0uh/1PvOUHfGSHDZTLAJ10abwkHbdtF
WtZECVWnMHJvsqGp1tPE+2SSgkGBcfVun+rEPXc8vp7kqk7KMFFCUMwrDCc3UTtD
3PBSAFC/M/fBdo90t6y5vrTArvK43Md8EudZ79AN6ESxvv5YW82KgTTMQnCTZvfV
vCWBj30s4uzWWK3oDSk54gGkwQ64uyRdzGm+/tfV0I1T2pyU3MhEVHjU8CSBlpHn
iQwmhu9wFWrFUon2Ghb6VNDBpRsTdFJSOgGpOU0H8a86ogccvFiAT5SF5vLzq3MU
oiTXT7UcLZ60yUdzKekchcnJ7sdnzTFdbP4fAyInsK23I7qvgWH40sm+OgBEuIMG
/QmzRb1YWd90YdLE/JtMHfogxgrPKWNfiVeweLGYiM5DSzKXAor6FgGWhjVqQY5+
OFbE9wH5cvQNF1uul50w1zaFulbHkIjksLIXSf+L7uAP/kGwsJpw84rRqQkSDxLX
NGk5KT3zYb/800nkgXxezFWatEMzwnVKfrdCrt4Mv2dNga0EKLDFrFnoXuJu6K6b
cLfd2k06l+rUI0eQxfQa4yvWOJNkdRj5dxFtzGL/4KQRe6ai3+wRajIVdpv2I4oj
uaQmB9d5DOKFHhErxWnOO171ElWe57guf6nVJX2phZ+ztJbKropzSZlrxSzIk4q9
7yTmsZtRtuEorUkhX0D+M5ngOOfNhaFc2yy/WKHcGJKuwD7rw2xfHuEaFKP7Jw0g
PQTGhslmBnC4Lwpme9WfSA6rAYMSvJFtwl2Kr6TynBW8z6tiJRkz/X5lsT7lXzuK
EMFx57PG+NYmy18eozVSS0MVGIejKgX7xU9snPGtBm5qB5T4NQrlgMVVw3G9W1BW
fxLmX6H+J5Ay6+aeQ6G9UKHEMibVkxghxDmOb1wrbqc+r9PuKn9TgG3HRayx6N3i
bbYeJ6U6nJd0UV/FgvPr+H6UbXAfDLjCLuTU/6j44AYPvX+KMsf98cxMgIIOKVRT
G8ONoyAoQTue6CRXt6TNwFSTcpECF0Lyk+uT5AzbfwYo6LWuNWWODpK9DF0n9ApW
5mfZisFzkQ9NPJpXQxselLXoXM8Oi1MdRk1q6Z5jWNAIW6Z1PjtfpkFk8wIhdScm
33NXzZ4Pp5kQIWrVH698CR9XPE2R5HqrIOezN2uqBwLCLNbB+nm67knBWfSh5J5x
DnJa8dRtgWqFGYOk4H6zJy8h4jCKodyPluo4A82yuZPLsoNe+xxaEEWDQsP2dum4
ZhNl6N+M5i9Cd75w3VyC6CJTJdXeHzZaid3LMjsiHN8ktCsX+03cj0njHRy6x03e
4gaKT2bdCqW4DgHarv0CojXAAjVDSbW7ruf9keHq4KKwRqAegponDg3v/j0pJAuG
ReC4TP2RO0VmFDinKx7146jHddALMeHyLWxqT5kRR9c=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xe0zsaegXAQJ1ZeacLMJddL4h9kigGeJVMpF2DF9IIiae7R2uesk1uD8Y8igH/Gr
3b+10uNspjAeLCoVh7uim8ByH/ckISEmOfKbE9OOYhe4sXJDxO5K+EyMDm8eUMOI
0FO9MFLfj3gxYfHeWLrAGHcxZTTLj5zzDS/5oiLSzI5k4TlHQzvqR0MLmN8+3Ng2
limTCk0LWFGdxacDuwUzb509OGx7079mskZywWkXz2vwfSIvjAhqE4cWiOW4Vtsx
y0By8N2JbRbMVilzKJnjt+haEX4g4q+5FVnqCrzMEN3+B2A+Rbi6wIqvIRv3lyiy
tapMwbLlU3VXK+2bbyOhilWP14UE+XQ4chcBidAYtc9J6d5bu3OWlknwUsyaNgVe
i8rT2Mp8xwF9CDSC5vur2uk+19z4yVxNkf3XKF23kGkJWj9JfPxY9AByuHzS5IYl
dLt2y/LFDrMYD81lldbIisUSZIxjLxoGsIGSxr6Ge2GPpRTSzIo+7ADx/g+XMjq4
4vHsJ5kLR7LMg3wVX6E/XEtqzNS1Jx2PB1aXWmw5DD5auWoHdVJ7MxcsqbSXQimG
B06Kmf33NvB0S+/tE04eOfmcqkiNC6xcwR8RwMoe5uwAUI54wpZ8vmcFmkSjdl6t
qquCZGXm4ehXAs6WLBzJGXvuXP7a0W1dZ5Cdd0oTpEXTIMpVEWFl29gOVXET2Fq+
jSvWipjeOeME6wrfQoodNvfuHdYfQ6luPiE5DwVyyABaxZEHA3YhHzGgmZL+3smy
DSQ51//41VoRE5p6wGOVng==
`protect END_PROTECTED

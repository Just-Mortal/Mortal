`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZdgX66i4F+p3RQA+jkDat2s5PpqMTLZ2HS4gMWFyUM3eYpujRlpzjxFVdY9U+kV2
kS8QKHil11lNDd7fS2QL+JeFiuMbludQW6r2Lau7miZVcGjBXN4NOowRvmLr+k93
3L2LDVsfvtbeAiyrZgyzPhPsD1XFS/7zZ3M7MRw+wmYU/YVCqfWW7IFDvzBJSH3s
3l0SKbaY/B184n/r1rO4aayvYKsRkEBdw55rD1kwVc6JZqN+bQkLk0HnK2ksK1Dm
Pnf7JPBP8daQhKLjLb1s1lfEUjzYOLG5SdLGYYDWm7cLel1169VG+8hLPeRn3WB/
d/Tk5yrx8VA5A+h3Sd7SzE6hc9zFkMi3BlFv6GQZRcxnZM1aTkLuQGa0Yu2RgeL8
JUbwJ3/UzJHkn5XeblkOzmzKe3hLne11p0Xt23a1MBKmMj0TZuBJ/pCU3a8AAuxd
/urMRY/eyfTISBi0fewTLDDAhV+/mOizWGKKQ4DLpEjbiU7/M3uNKCoGLluilyXn
MCdMm1EcgQYpPMroZ5EYjS7ySbPmE/qosor9dnJaJWturLe2BWxkEuAJp+y7foQF
uoHdosLSA99dKSzTXVKzFD2ifBsEm+ZcJEg6yP6p9dVjC7E6t3JPhqQv7wm3ZgUm
ERBg0Fop5vbWBK+UloOlX+7V5XHTihMTXufASSMP4myuam/sksrBcAFtlHIxkdE2
DzkkkEV+jRGfMiEt+yEWDlqgxeC9A69g3fGqpXQO8fi6v8l7OBc7T9/1DwvfJ+R4
nEHJFPoJ6czuQEMQi64aod/Qhoj0UlVp54W+arMtN91ct2s899xzw2YoEGqPnyws
bPJaMczFA4ZShB/lsSF09UKfjGbTDoOBxb678o3Dn1us84ZfXU3lABJxqJWScNNZ
uBCeWPKE0PHiiYBmUTO0TM2djshgeteWdtMu3q0xgD/RkxwqxDa9t6HCbPUUv/6m
2L9Hl2/BkIXnbgM4sohyjjKE10d+EIMrabXEl3r8J8jEKZ73WI5Sw6CMCNEre+Fs
4nIkdpYDA5Ix6aR+pv4EgTmgc7sC98QfIZ2X5UgQTSkmDfTz1BzXq5SV5+tgP5Mk
roD6sK2YD8PhT2I/XVyddRwMErZjSuC4wSXsigmN7cxIE2B5jpIrz0rpUe38hAb8
u1SwfZBu+ZE+SsUI0PynskP36ATKIFgrLhTlKDWc5kbTZNEM/g01vUAfrtKrEF7t
xv1V9DTGaznsgHO7deeP6QW8/7wKMPnNl2Ta3r/DxnpUqFZiTX9FxZRXsYtqZG2H
Q6Y7U+dhl7AqXNn76N0hTnzlR4CgNXFxaISUpYVFum7TNkUcav/ODq/fX8pPRdtA
SqePPdVciavY5wYXmJ41c1oO68efSCzou1gXLvRrE1iDNGZKD2fEteN3QQRihPAk
MJWpz281NiizEfi8Wg2nbrnBfr1Zs+IPBZmDz2lB3ZebD7wGiWkjYJBnNpSq11rP
zVeXRL2vrZL/FZw/Y6ehaCR05usm0/hZ8a8xfbt2ZINOJ8hGoIWsUHBTKTPJajVB
zQV7TpfX7eKKuPkNzi2mOFcVxkHIUrC9r8sph/6RSOk/uwIKttvi9rnZBZAuLii3
alHQKMbIIKdG316q9aOKnO2OZcZN0WOwsubN5sSvT5hbpjIGkZN9Hm/GtWRqL6e/
rW0MJYK++EjyjrNS8VvZMsh77c7Y6tdqExUUWD+fq8tNHczWhmLSbhDRTqXZA/1S
l3WOz3rxOU2pC5pA9opvdVcbLT1J8PsRm0wbdtixM0vX7TKOiqgQYM0iZF9I527r
5n8kSYMOsgYZvjY583/LpFh+TYrSw9webPYkA4GO/1lpWeNMZsrIBdIkiEF+BF7S
dYsbz+dOJ/yWJfwtUQhycT9rBQQ38oXAZVFUtlSdwnVGxhoUY1oiKVUwg37AVHUg
2aY5WSo7fFrzQdPaxoTVeJNZNiU+NMR2b+f/9ojuCW3Iohz3tiLB3xF27lPrh1sX
eifGSHJbgyhYGNVn/p7oU73tM9GVJTpfUbY7pcC3WHpNIp2178aBQeCpOvja6a6E
PixOZwUxju1LI4LfgsByAHgH0xUQMgN60nGWUfddmWlqUrcOq7Aa/Ofx847QGl6b
4q/Ms7zgljZDrAb9K4lKl7j/HbPUMwWBpJFny5fT0zxaMX8NYsV3ni2FmOlMVFAr
uacItzk6NGnidwEOgB/u4CF7taBGo78Fhkg+rNI8HxL3pNquJLQ/QHaxLqsq7xM2
ZVTM9cuSLL9ZrkDdln/6/m5ewjg7HwMnuEdWnzN94O32MgqNhVfA6uUybqB7cQwo
TTwwVkC+lS1eWmgaRxpkx8nCxBJ0Y53Kfgic34DlhEefvxWepLjCltBPAsTy+IQu
HNg0Zj9j/+nZIRytsery6gpcMSdkv64Yog4iYWdggIgK4WRa8+gDNu4WWDLY1nyz
8jFm8WUVr9P8jI40nXts0ZVdjPKbbFc5qHn0///Cr4bJB8bKdG9EshgylkvU6mRP
1ajk7MrAu4Af7Dc5ZviGjvtoiseXJQjeMLzrDmBY1zjjxL8REQFrVJTjRyGFndx4
F4YHoCqoO9/eM1zK7dHVm7ov4TBhtpytTgjQCk62OLbNQ7tr1sYgsCE38Xq5oFV+
F43DXH5EvKZtoE7Kaui+Jd4cfl1t03g/GhlxllkoJZG3ekPTJZvZeELYX/SQumJE
9u6sPcpgQwvsQw1yQbSR5B6EQAerO+EFTHHCHEuzYqyIkc8GlsKfLzfPX2E9624m
DVt68Ix65vfyKdYGKj5P+1XnBU4P1ki3GpV3YjpiX4mff9AKHeHz6Ys4lHiIFYuR
9V9xjHoVjxgT1oR6OxeV3bR9wmuLcnsq8D0VoZvHtv8Sj2EFUVzMqq/ftGv/mITC
HpLzpKeLfN5ffDj5VJP9jBLBMOVZwjxgcYPyBWpeGL/QOsqfNua5lSMgv8RwKKAI
23x4epqCcW4Yjrk5Uc+n/oQ/M0Ekoko8kxEcqohZn7tzqeGAkiC93Ne6HFY0PFO4
Ky5IDr27thxtB4PEX7n4jC+Mz5ojd8rGHpQdIKdSz7tJAdwsNAtASWlfO0sDC0MQ
vatB1OQzHoL6FYnZcYEIx5eqUi9pMtM6/Amvo+Ncg5p9EBzKZ/PmJIvcoi4tdNam
nETzV/EODpHbEha/8SGHJUvLq+OIGUL/EA3UmtZXnCIkuJds5kcs8L789/zYVWw6
IUK9p8UXJ52olRezITPM3G3PgHN67Afg0BFzgS/bMHYwyLt4n3Iw1RTmaYDCFhM2
o3XqC+4zoJNIgTtqrHpRY7aV5MvFkVqxO+xf/tKluMjeX0SSebdG2mALJqTibY+9
qXR9luL6fJZD2IBu5GIbNfvaIgOPh84gZ5az1QJE2iuEZmf137uCReNZFHG3d978
k7kG2ibvJ+A7m2Y7WXt8+nSSGe159Vp3hW42JWoY0xAkDkmDBwmxt3yDvJj8Qyqt
k4P+DIX+u+UT+D2iS97J0zC1/vqBh3MhrUHxXKcdqRjZCzw4ER7cRVVHW1Tc/TvP
yPVvUf+21ImthLFzW0soq7O//m9Ucykukt0tu7ii8m9V/mSwnrqv8aXnKfnQLdXy
lQ/Ipx7YxZwlM4bQADJNeIiY/TNDEeM658IkpUMQOCWoCd9H1YCNzPBH2N/xEi0x
z+GcHg5LEan6a8o1lCNcg2n+a1Kfwc3j1IWYxiY3tdMqzf+82zJcCm4K8BwsBTkW
Ktxf4V1LA4FhPxgQeRXrwBooKrg9KQ7tNr0ooJ2UrzHjzQls8iKKciGZe5wUL0CX
4eFtnOFr/YN4mRtOlu2qieZTIzKjwqJ/accq02MOyd4CKzt9U/UyTMnsi0m8au11
9UdmLNoCVRB74vrJBy8CppsSwzNVWT71m6DGkvf1sfyqwghPsCQQxSLl5lzBECV2
XBri4XM47KV0OKr08+Wb7c/+KurYOIL3H/mnt8ZR7IB5pMPzJD1nIODC2+br0RCX
oZGbm8+xZBiBT2Q/CnGAk5TWzX3cwVOq4ohGzzj2h82bu/h+mTgY6zUHHsHWrgdF
WIomDum/+4FT6Ggqvj9ll+dbxYpdxSZmGNpFSTDg5CvxVjNL6gsacWH+LAH1VPDi
39eVdlyp2SkA2P18M8NRpkRJAoN0Hzk4wOuk2S67YtH1DZVNEsGiX1lUyYOyeW8T
WoVkBt0EBukOZt9vfsZQSWDYzp6k4dnrGZYpZ9VdUzvgEDKCZ7kwGQHTWNjanW0f
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hMmONAi2vcOmh6p8+m7G1E4cQTH/aCQdvoNpzBOXExHa9juspd0ILjXS1zVclIKL
m/04IkQ9qA+pdqL8uIELmfJ9IcSR5Uc5kh04gF1qlM7vvGSIpxTXPxh2hChWNhpz
TNkdTjUPDnE9cwGHr23z95DMFucBcfs2BLleGFU9EsRsn4ZNUaZF+ZkR6X4W+wEW
cFWHaXPUm08bcCu4GZbgEQtjExYcm6OsjlQch4mT2pfTcTBeqED4b92pG+Rw4sRw
bT7p9xUQKsM4e0YLdbRn8cL9ZLm6srF/V2LFwt2+yDeB0+Lx7mZ5V0CBt4RLJClF
3EMIMjmMrmTCv783LVGAhowsoxO+6HTSsomQn5v4Z82jVhlj1cnDo8VjrV6PPk2k
y40rQWs8AHdHY95KpQOYM6m7g6U/qvB9XNtK3qDOlvXRApd5kMk0r7Zvk9r8Og3j
tEK+Rv29g3ooyv1G7ncCCGNEDIUmuAfkxsmmVI8PyUnBZ3t6zvj16//yx5ZorbGL
cx5JqbJiLE5Pyx1phT3cSZHktwfoordBfIUJ6hU1rKrTGClJh1ol3hRIZ/9nhEyv
s4CaUS8+TQop+qDJBPpRc2G5wbV99aXq2emjfKeeJBruia3eS11F65s0sLLx9QIy
7rvRRyuNysP3qZV/Mn2J+uVFDa5fF7XSK74kHzynCNwx812ohva4vfFg9t85087Q
cI0kL3PklxoB3Pq6HDaLpaPkMpz16YC0nGcdFjcZWJM+t6eM/aJYFbfMQmRTbnI6
tGYxxtmX5mBPERSvclmvmAo6NWD6GobxNxL8p2SyqI74RG6WMlq6hc36YtuIuAtg
qITFbzxLIembe9r2Vrxzs+K/g7or0LfCi/EDwoFGQnMhuZ6umCEMhuwParKq+KAt
lNogF7TKPOSegaSmFH8CeQhzSCmrYr4vv81Q51BrXSOl/A63K0z2ouxaDAeqQNHA
2fGDIf5zudA2O8WdM4jcs8AAzdYF6UxAQgO/P8ZE1FCAnRfMFhF7aw4/Oqihh0dV
hUFa1YICVzFIr8TlLj0uSmWxDb2M62UAIwWL0XLYz1QaaEJOU3/F3B5uRYcHV8vF
pqrylPwlyyT8Sm3FDbASkbDcbIk/WG8xx9F1ko8Vz6vsej0xUj5vvuyXzw9FQGsE
iuykvcZKhwHjYZg/xiuH1/pmGWgPfjtRqmskRP4Q5ATOU1csZS/Qjs4cNoZRoOVa
4p30/8QPk68ZT62uY1mW7VZuTGGbXKT7t81a8RbrUY7YjEAAj2Tz+7L6gjNQg7ec
/+fN4RfLIF3FAk2n6JK+y8x6lfO5kgDE9U1EAEauZ1Ad6bSDPA4yHclVNPSIoeMW
Ol/IrA44jfgDQ9LzGoci16ZpknKEQ4PLtt+FlO4wCEHhovhv52O1Ozst+5rQxCn2
cVKydADF36lV2a0knqz6UwFSR9ybbTU4obrQVhkewvXJwDXu8ndssvsi9FlQvie3
7kdik83MiW5f9N5/v9nmHY3drmCt4JR3WFweixeN9ERzfaf0l9wEA/oeQRgEvwS6
xadk4dUYGLCI410km9mpzMgbm/4n2qPh0e+SbU2VB6juChkrksDxTOJ4NDmyxxkp
JTgOjp8ImO5gPyJkpAW0Rc1Q7pBpJ6fKnVeOlhmCjp2JOUDJ7zVNEHYkGJYDL0Dn
kMHa1d8AzSmwVkHeSrTXm0xj9VcKm11XZYTNq7o2FikCsttTbSAkbm/0QVNBgPiH
QYnR9rjmTmnU13p7zO7I3OK9II2FhFP6NRUjHT/upWCkGomQXk9o0khiJWLYV8p6
ZJMdR6SbSXz9LijBpKYuyOVBZzcT50/KLAY19qbWjXmZZTOHCNMsAVoYkxHDR1sr
j84ucQe60ISBKN/LvznAjiVMOsg94GKkvPk5qgOVZibmRvZ7J0RrYo5LI2X7ZsTS
wZIC49j8xXbEDP0aP5H3nCX+huCOck/rHTHKoBHUZjtV1kt/Ob4wawbcE31rnx1u
ymkzBVq4/3dJ1u7ClSXV9AlO1LCOb7mYpfuC3exSo+SGTzRscbvmyiTgID409/bR
ROjEUhjl6Bll6de3CTfc2WCv2lFKFOQ7mbMs5tbEbtR1YBhgzNoaEeyUth5fKvhk
k9/g9we5to0LiOpOsYj5gaN1/FrZT+6nZRzRhdY0z69mYFQu9s3j3E9OnyEpwG+B
obQfgbpF6V6h2m00VQ85lZ3w53eF+aEefdyjDBNeYO/PvDqfRA9Uwr3eISquyayx
UreuUDzzo6jto/XH0ID5V7PhlZLjB3o/PW+mmdIlH72GY/uy5s1SEdZylUWHp1+O
qtmrsk9yhrzO7TecOrr0BayUcq6zicMif+v0kADj15KBX1Zwlz/ap2PvIdutmHxs
szRI5wxGJjXwv4EbLj8WC3syxF9ZKtT/5uAuJDbLAlGjGa/FJ3srLgcRoljRsOQA
BZUA2v34f8JHbKcY04rl2w3N7ERdyy5F7c03iI6XZlq0B84Z0g6Vh2hRLT6M5BEC
vr0SNq1/Fk68+GJAmiivEUyWrHbHHaSFa7O7jciS4lfqdNv0pUaXIOB/IXREyOLy
B3D6MiVqpmIELYvrBOr5nkugD3bNvMLR1F14jy9Uc03/pqAdMxqNgTNLUNZS0N0Q
fadyr2fQ+5qYqalYg80VvQMoK2Wvb4KRTY5ZqilNO503wS7A7uYNKR8R4yWQHqfc
d+fqOQlHEj6qrLmDjnONR2+u8WoXaigWpgiNQmvqWlA3d9Rre29A9BXGaAbuS9MN
125/QHyaL6lZwqERN/yFA1QST+JiKaJ2CHKiN3J3wpfGlZgpTYo5/8zHI/mrUkiY
Kshl3Yx+azPLd0skbADidtoEgKNPDk61z8MBWh0rmWcBood6THmWdSyz1XcA2PwF
GVOepN9a7HvaA+a8m+e4QU0jxq/HCukNrDW4ZCBVx2aDOLfOl6kWsrKk5XXvJD+p
h5q4fktVVmk3sIDEiuM0pFgkymfP6NxB6CEdY51/Wa7AEkuX6vLH5C5MkO0qJCy6
zqp8ePxNn82sKguUgmeyT6NsEaQAx3/hELvFWIvAJMZrWPptt+gEE8iwxwlxQ32t
DZpMZciuFX7E9SZMkDSAcfc05iGn3Zh6qbx+OO+JlmdIX42WslKQj+POumox2mOM
D0gMk2Zex3iDFpdZ+ooLR4nR+yWEXnyhDrB+h6pdfSA0vUPcPQCKn5fY7yGQ88kl
wilg/VpxAKAAv97g2kpdCWN2kBl0V9RbmEEuVghOkIdJyTc6NZvJDj7zOZYuGrXC
1AmDHtulyfC9E0a6NIxP03DxZpMKWrJS0j+szZF044EYpGCsokfoWnV51RX2cNZh
dsvCDRb6hLEaLK+fa4zhHiGkttA/KMbCFCu+YNOfsm4fsqdnaSIA/m+iAXTiaXmT
ZFZCLjrlEq2J/ZFpHLgXOHf0syBrZHRhi/QRFgLkzOPcClmvIuNVaJ5YACxCG86d
SJVJDq19wRPCVHQpxn9123jp69cNwRT5Fy7jWhvcJlI57fhMVjkztL1Nva9ZyK1V
STyNzq0P4TkwSFWBKCvA62jdJS7xRRrG193Aay4CMUzu35ogBs6I4TZ5kLCACesP
IZ3FowamMf5+VtoHQ7J0No/p1ftLsUS7t+5FTZ6PWwiCstyA89zTPXsZCcJ8OWif
2c5hnE7Kx7p5fXLKH5+wU9q2hQI2IXnqp47Av0JpI0S+RuLKLRWZPQk18wOgnC5H
w4abPQkoMDE/v0nG7V4FEELoAlyUJszvXJBipWrNEdHHZ+OFdpvUmQfe9THf2kKY
Scq/cj3WRr7W20ekMmalSHc8/U6Hoy8s3TBZk6X96UBw4ZF/qeCksmTt9cwjpBrX
y24vNSFbNlCusOA/kfaLtwMF8S3zAPjyByjUqUcZ8tlmFES9Pfunyodpee0CTiaj
WEfc09hVqKGIllM9fho/mbojwJjJQUh8eAob3wzFY5/ujHY/PUd9psIvbRARMk0H
c/n9MOzSM5c8+pDiRwpsqLmP92dvjLjnIR8POCgjNY2EQ1r28N9lUobLkx/6Kvtz
EUx7VixRlSQfQvZTIxpAVJDDOQfnUb5A8nPry+CA5Bo/eCNJiXoGtewThuj0eN30
BPoDKvidxXWfpXSxmAZBkZ2yHAY15Xkq5HrjHEozI5z4Ty2hu4fK1W/PzF781qvF
O5O/URDDC2eUcilGcinRZ6SqP+GNsR0/OqYXeu1eBuFxBSliqpRt30Jw9TMRNczR
Fsh9rl2VoIz5FjtIzagoZo6ELJv2swJ+KeF8zMEt5VmqvxW99b+uBzp1ZwR7hhYo
SW/VfnkfeQIgoLyvHk8H1jURkDDGscTV6jUatqKho3tKFGgUow0pJ4XN+ce/JgBV
FKwUUiwKqR/yng3RhCH0IYAc/AY/P+fvqSxxRJCZm5P8OYTJIJbgNs2rJsPBwlKb
i8p+QMcGA3lCfcgDjUzLZ6X/4VNA9oIiCngqy+Mn9kBlkEOmpid7n4XFn/ajsryB
V0Ig7bcgk+61LhvMYokWB+lY+xJGiqRc4ewdd/csTYE0VIiUDe2XBIihvsLV7Pkm
5duWw7q7/1jYVrLi8o6IYBb+m3I0VJrD7RaNP/nshCj2A7EmdXTYQmRZ4kBdUFny
lxU5HPpxp3tRv4W42dUqha9cwoT6eC01MWju9KhQ8pOhhZ+qrWX/gROFQ6Pn7s0i
G+6zUomUunlFWjXM7UwEZgetSrtNqEJKZ2KPFztoB1yt3gRtEu/iTgvk3jBCakMi
FmQKvEPy2rwoZ82xNQZOeoVgu9gVDkQBkwGqHdWuPdYwQpF9gzqek/J47shqVR52
IBlkVC4W1d8Cl8v6Bb3FyjJs2OW2+0JzwZBYhOa1GuBVhPJF5BkxB8PsxbhG/Xz5
9WQgAVyvLUtPn2UdLPgD33v8Aw4/vLCsh/f9oN+5CYbVxTJPDURYMgYOVwjAxAPy
ArmV2a1mJTGtiWHoIeoa3hylv3oAub72DsKkRzO/VUjcvEZQQV+0uFOdHTxCghxC
7c+xhi7Ik6Xi5US1ylx01W7jFf1iPPvxbwc0A1ll9vNtjDeqdoiprDL2HotNW+Jk
z7w4LrQvrpp2U8dTSv5ruBvHk411p8mtfOvnO/XCNrOxQQIkaFxdpZg2cSiQ6bRE
bQPNP/3QoXxGzGelVBH8txdHWJ/ozyRjJ2/2smrPKHz6wMjBpAB2kFqMGJcAlAx+
BzjJN+iSSjl5ZyBV/wwxD8mI+tL3YUwPR/n88P3ddc9NVeKc5yW+oiLlYLak8vi4
MErm/U6MWAvL0xbOIEjM276q0/TRN4Aj2mWj4PVfuq5LXjyt3g7pwWyGdxhgkvSG
OXm/gRDrDerNtzwnB5ognQHf0oSX9aMpP7GrLQjdAVc7cLiWbCBx6eqGGZm1+RHq
zDmGgeElF9B4KjDPZww5sHd5pvSkbnO1m1lH2o+EFn4U/dd9d1snoYg9chaasWTi
ltc5gL75RLn8XLBsavytDOoAfUtdzdxaiZNePdY7q+Mwd+rMyK9RWdjOjEjQEZN8
5O0e1FIEFUWvBWOlyJVlVFY+vZTyrGpoviXehyORTSy7iV/XgQN0k7rWCoKcsYSM
yhT35zHsVBni3zzBp70SW+cKFCipF7zGjxIkfX3VJYphCPORIo4lBUSxv3qXYmHP
hr89qsp98f0kKpuYK9icSXeDqEiulItvRJUZAF0HvnYqpLX108lhyK05D6qdFrg0
rmqzoqaJpipgzpi7E80SctcuuzkuIVGaifcAqm8prSEMC+pxdmkG/tadyyXMNC2A
dhYzHoS2ozn5QDsA9WpuIDNk8EuASjHNG+EtYgM33gmbMie2CtnFbpATTHS4eXCp
fNIaBuZ4IozeXbPRFC9au7JotHXpbgSTGk+raIVqQuEX3y4Un1/zdRJtA+bSOvuW
9pMZvvphrXgbuOodQcqptTdZYWg+7vMTjwCb5prH90azZmUoeZ4XuvlFOMZ2TODR
ZeOBNCbdoW0T7nIQTVFGIQm3M7mPTSIQWKisoVDngs61m2E/zKiCrJ324syxgSs7
2+NE1RmHOr5KHmOnK5TV9EGiq+ft6g7oP/CKPVmSU82VumpJDbpAzW9GpK56g+a+
jMXPSK1c1bPrBoGTLdZUYZbODuww6n1WsQLul3Azh8yqPVL4Ym4bphUGe4p/qLld
4nz94XjFzq5na7C/kAhQpBZGQJyxqkyM8U3tY0mWzBT/FOVcmQ8Qzm4t2jmxPHtw
GFuM0IR9RVjm/9Df/TdeRDg2sL1rwvV6842wVe4+KF7fZDZ1jsUGyHWlMu/50OmR
R1zA7E8s4iUGnsmeexsfFJg/m7XkiQ1KiI3IeoylCYocwAzHiEjH8aIXV2qIT/tQ
OaX8SbIo6TQXA9KHD+N3C1K2W3awpEPGngwPpWfnLlsjoY7R/9Yds8gqpuCEP1f3
51FasS5kLU3uZwASp1YjOs2zJXXuqAu5uf7mX3RC4lesmW14wDEcvxQn7Rk32wa5
gP6oncbpsRBgaA4YoAWfo67WIRXIDjXISdD8R7g+VpPZzIIRvsiJL737trsEu1h+
Vuzl6ar4LgfCQpsEb59k53RpAnWzI/S3R2Tnmaw9r9A2dp4rl1n2fOeOToSAGmD+
EDPdbmxtOAYWY+e4MQ2erKsWR/aeOYYQ+akNE2evJHBPm7jBv17jqka190pbLavt
K+XQ6fk/kgZuaxyztEpXDgVRoaRGocNGTHXdXbjRutEiMa+6HTihpLIiyXo1tdVm
dXo6HehoktmXERVFz4BqjY/elm/lzApuoVY15v3+uRWVU0vU02zL5+f66sipoUsQ
jfcW7D5MMzWgsXzEj8I31+gntbWti6zmlQ+0wyrFhri4PpF/UPN6EU3r+koeIjSU
IpuodRhviU5FD4Hv0nBmfxXuopSrF/USqLuCPhMBfKXRaNpE1buyWRHBJLMTe6LY
vwu6sfv3X3yAVysTDaEbmrOxNkLg0VExi3JPHbqQA27ljc6Ek51XokBuA+F+RJZ6
ae/5L5/1PEnFjFlzfbyBTyJkFP9Oudv802aQd3y8yY9PdYtbJ4sqdR9ElXk9mGEs
aKwIyF7UoDBWfPF8zyngjE+qwk6UwDA+DtvxR4cBUQBN4JpcIuInMnWEjR3Gaf0E
IE2+la9l0oD+axUhD2z+VBc1cWISOidIskwj1fa/zwO23lY3YGTdUZAhNDHKEUaL
esorJghm0/pEvWogXq2aN1xmx1B84Qo5rtMvqaStzmQbKFpmhiqXP3QfxVIkl8iH
7bdr6cBeFaJmSYaYrh7aXQPZj0thMGK+FecQfakDkuaG4fmN/8TwGUC7YqHT4xXf
ylfLtzYWNjsMFERnHIP87Nm9mkUSsgFSmIDbnfR3/RXXZ1MsBYotpxT1KL5hx6Yv
Yr7sbvcTHAigbtx9N+DtKPj1M555nELeN2wnvtvENOOshDY1D9kmBcGxGcm68oFW
tWe8q0bLcSCpE68EEzP2oXAFenFPQ6k7PQeF4NpQj8L3pYKcudTjGm4+hWrOMiLs
BDNPfl8i1IKsDIQ+KLVU/+Z5xlOZs5gHS4wFP6MP6Fc6mzwyFYjpLpH5VXUI9KvG
AW3HMkkjv6qvU18DYX/yd71eNBWKd+Cwu46Gr+u5hUJyLklb3YgATdwC9X2yyBO5
Jpx1VUTQQxxFVLoFLr6wYq6LS5/3LRLIaGKtLoOy62q973dXUFwuWrdpjZ2k8srZ
DuLOiQlD/OxOzXx2naDpCf3Z0i9gJjyTKcjxw0yyU48yCDAReMCcvNwFDo7N1K09
wq2gIc+eVlyvMYueGK3u+OqANWQm7EVnrXbNDhSjtfF8clK95K5W1PdmAbsUQ210
Fr/rgytEybKvxsC6fTagMFOQi1s/jCySnLcgp9hiCzydKw2CBc+WiYQA/WAx4cob
nW7wuAQ69QvobkaELhTB/0jPAqdWceCxDE4LWPnJA1coeDLDz9NpcswxWEHon/PZ
riIt2CPJ0iKXAKgITGxJ4BgLJ8IQstbJNIH0ulR04xObaAjpvOQiPoHoPaSWFuYM
Wmx1ltDDTEw0wp1XOh81Ksz7r4pQICYnQiXz/siemp/oF3yjLzcMaHXSZdcPQkOx
y5ocOVu1tr7EbGUF9zmqW4AZQY+G80VktD9y2/eARgJXMVBElYckIXXLaEi4zFsv
v4XOfdy2byj1z2BW84rFvO5OZLveNumEVUdRqt+baNb0bL8vuOKa/lxsFqe5Q4FL
ZSj2zbZCt7E4KR603FEEiooWtPpekCF6jn6b3nQL0CBI1ISlD4zFCk9yr/9vg9/A
QPTJmi3YricU7ZFlRIT25evgCsUD58uodmalwmvJcaPrPI8NxLfsj1RKWLaUGGQV
PUsnllBEJCMGQ8Vluq8ER/upOVg8YGTKbFX/mBt/8z8SxTzMf/1igpfrdvl3VXRx
GCYnp3SCUSQwvW1zydUGXqKPUJsuZvgWrgOTVS8NoPvL4hPAguYinOPfwaXTJmnF
GDhh7UpQMXyVTpnlISZuO46A6mVPT9md0+FgWTycz9GFAw8cNO1FTd+0rPR4kjVp
W4h2ErubbzltREzGCb0yfZ1Ff0HFSU0Inn4htlTvuOk=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xq5Thp7q1DjWCLTTmnrsa/jJE2jRnkx4/Vl6mbGW4/9ueZdYP8u3NRuxH7ZqyXRe
lc/LYENfY6IMZUTwrQDP7qQbJB2QKo4hujLIXeV19Q08rVsW87R1l4tD8L0K6Xhb
nDNrVZDPQOTSp+YISXSVc2rFkXrc1lYVAiRP89sY/YqxpExqLjFdxFPkY52SsO+/
xUdNla7wKOspaYF8QWgjTjjGowHQDFoMgVeoKJdkiwWJng7aE+bI2CFCdFPDBD8w
imogV/s1I7UG1de+Mhd94WHPH94IvYYFfXqATTRFq61mF4SWQZr9jp0Nilnv1IPB
KdLNIfm/z1YhEXn4pMCdi52L617CXJouJfSux7K4RKxyqPo8/EGUOl9zzL8yAt85
70xj4hfzD5PzzKkW7K1D9jQd4kWvNQmCF9pJJk+UHs51jjq9dHTxec7xey7W9sjn
G4fi69wGdDT3L8cF92g7NLDnOashb3V970Ppqu8CW6oOnBwKtUSHfL5Rfnr7uh0T
0BdI5MFA9myvLlASoxPqbUkXsKWA48M3Y5J3Ex7kpt4XVkZoDzERdToiN8fPm316
vQguLRjoBYQEMd3Jb3CxC0dl53hKBjIiqV9EAV3pKU4BKhEQjBxCnuufwIkKROFt
tf+8/PQ/vb/cGsaSQc1Ey+zkH2qK5ESK4kt69MPFT9rgK2RTF1j30mWnfCB5c2CF
UsrK/Z3TunGvgaDilIA4Bxaiood2zpHcandLEcIko0lz6yhqtqkVGBB6F11FiwOH
XtuhWiYERq7qMLW6L7GIqlM1XGIjOsor6uu6Qz3+eOFNqOARzAylOpxgKLaBSubq
VIVqqpVaLeZsRJ2AdzqrUQWLEMhr5RhUr0aSu5QxWyKLkZgWdJ36WlFtH/saYkqe
zpiBJ/KHHjR60qk5tJvRd6XMINpDgqI1wEauzBjX1mDHLS3cFs4MiLblwhaLepei
t0nC98cl68Bl4/80pypXAmQlP1x3RR5jXaZd1qnkXRTHiXSgB0R0Us/Cnz4IQF47
JmjG8siaveflmDTJzD0B7VRoBP6BQ6qR0V82xWWMscuXvLgsuXqo3+wswMItBt53
fn5B9Q8HOuN8ggOIDk/Ah4cTBbNQEGMMabxzzWg7s8rtNbC6lRhzkxTVwIMqQSDL
N6OPGW+lR7JIrb9v5oRwSokOhCCN7e1Id67Uvd34m8BVuADoLfmUvxLAMNwh3d6B
TptPqktYd+3TNpXIZ0+P0oH4px5oN0whjtOwD11LQxh6AGafdE+W599Mibm9NQA9
PWRrVMYB/jbpN8rS2XoixCXUSy0G09NoKlyey0nPWFCcRhsLiYQxFsitHbJ1swNH
Rs1O2fOqSjActGe3JDkBwLeTxSM+vdxzsE+T0szmvC5j4OdKIww/9BrAwEIn5gLl
p2dtEE0DX7bTWwfybaBaO/Ig90O8z9dxP8Q82vzM3bDozvmEGjXCHxKcsZH36ob5
dnYV5SLSCcSmnp4pwU+MoqYXc3OxLkmRJ5RNXf3cR6w4VbJ2KPbnmEEv8Q710ddd
JiUwI39/KS+RzFpJbN3CLC2oobrox0MeCI7uaMh9UYKbWbQWNJvZ7wlB5mvjw+5O
t5ECb0ve0uUYGL70ke6shyZx9HahGwozqp4B00IvpQRtrcKxE/sxlOucJRwtphBD
0mSRaSM30yoYtkxWCQoTf/do5MztatS8VbeEDl3rBXQWjK7WjM2l6xc32k7Fxmhd
+C1VkV8mFuXmOa0cIxkykZBBJXB601sqS1sQH6pHMwpHGe3fVDmITE1fbms2zY9R
vPJWWGLYDdW7emfM3E5eYKK/Ew0qfBlT5uCvOdUNuq2Yhv2ZnX22DE8RSkWeukDz
T8nAeNWFa0OS8YLDjQAbCVN9GX1BRtB1MO+D6h6eoMFLG48z2CxneCDUaUfeDxSh
unPqwR/Ls0XNSz6X5IVQkLhuSKMYDIfEGyj8OI3Su+HtHwdpaqwaYTTC2X+1auql
d6ltR5rmBXTkmpac/JxC6yznysvJ4Ex0v05PBs2JgED4Ra+sa0Hcr/D28FKg9UAN
TzsJJbdpfIHXy2MbTsn7mjKStjL2lwR4m1B9HUEHh+nvDh3qsdEVLKlDKTBPwcms
g9ooxW6NSOTOnxe7AEjrB/undszMVXbsuI2UV4qDlOzkU0Dvt7UG5jDUZfJBMFK5
D7K7WYrPO0OIKseD0TuqHhGEIoa0wEnT6YqNx0PA5VV4KliYVAORJ7KBy5fXPRuM
eImJUnKFsSppC3Ge/MlPJgwCdfKW1KpKKxjXkAIG3qMEF4ZTAuM4D2Z7DWeKrbhb
wxmPoBCThj+Onn4QQkYC3JUKjRZQ+dOGdFycrmlwv2j0yotUIgiFh7n1x0B5GI/h
TXPlG+FpzN2250+3FD9BfWCM8TQ7fuUXGadKfHt2bBJ+62bJsQWbwD92Urx/b+Ma
yknz60kmuwib868dQNzzrBI5GhUF/3oChyYI6qfwO0OXyNaP0STL3X1VgHiZMg94
BwLLxJ4A6JoqBEb6xjOrfWl7CoAZSNf1tJmA0uw8kcszlcqDuwAIJ0P6bxXhfugY
tKoQyNkmNxKh3Uahv3D60/f5irVp5/JiXia3vEO9LfJKRAxuxrmSqYQ+0majTOnS
tsNErGtTjNSussh1YE2sVAy2AMaXQuJo5xEF5f5fHoG7StyyGym7s5qm8IvnEaDa
FpRT5womrFG8PWzHFaeYQkzHa8GslTKEFDOIAQt7uMt6UpEuqB4jVnflavJA4NII
1PT4379S8F9RvLBQItXXKpUerWewbddgv+FeBFPw0CE/mXhPc+qOzyHsqPQkcTuP
pihfcaGx2YIMJsfLagQFbOPzt0p3XSTTYDXgJC5NzWR4asn5mS8SwfV0lwFavnlG
dSoGcXgZXSd29yu3BvPeD0p7XE0xq4s6puKLpECspZPV9WfdGraQo1KB+HS+qmkO
xnvr3mHneoTsKgH+4z8Y289AoNMvvaUs2f9dkltDB64ZAVAuMfJ6d3sdiRbd3H0V
1+qcgUySV/g5QsQ6PeRB2ehyTl9LivJxJEJAAwAXX1FFWpVJUyydw7lmYo3JaGfC
2fZhuvn1t6d5pecqB2X4X7sDqF3YMECXtPmzKkNE630jzGdpdxxVWtXVGeUEPPVj
Ywu2PzWbuk7p5/zfdZ+1ZqwzporoIkaEVyp8ThbGPQRj9VSZ6Q4uQNMpJyjW5n6r
/v1jrdUlR00QgcHGKde7OeJeYEJtD+QWp+jvENP+RNiL+sUi7SLWFJTq9xuKPP6k
loBYiZn02uAYSLvK6blUQmsSu7KxnmNLGVdbJQjBPrXzz7Sony+kgjdoHmSqQ6So
AV7oXg/heTafgpyLBP5a8kr5gHDD436zkfa9WL1+1co=
`protect END_PROTECTED

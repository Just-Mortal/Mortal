`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGbzwrY9vvHL87Bpdrpe/EaErjSzqiSSFQayqVtwzEyH/4bZ7ovBsnxVyUrjcRZX
O+nqdceM3VDN50CA5K3zgesvGnjX269uhynHfxp3eh5t/yu2fU0miUAPYy5szyax
4S+KMSX1qcaAC+28hVyApAct8xSiomiJ+5rw1XWEcRZyCtqB9vCAAXEIG2WIfvLP
UaI0x+m5U7Gzi017bAQ97GIS8J0pDbmH0lVHEuc10jJy3Qb57IFqqhZRZ+3WFJFC
sxvhBZzEc1BOmvnzxc4Aj2Q4dBckeJN0znZqB3WkFHS5zKv233PJvLVHIDyq1sks
KkicA3CPezqH+n5eYL4NJ9MVGciBC6ncU9mEriIDKM7TMHqr0eIMEj52vJjxvYLF
BXblb3iZhp5d5cdV/zMHeJhlfaQ/GetkETBXWQBMZphp+e9gew+GUnNLjMRCn33m
SdHTh0HD62vMg5VyyV8gOhuFuvg0toGCyEgBNOb2bwulufsCzkxNTpCvegN9H2Hh
ejnaqlbJvosx0n7o0V7JxQDq9KYpbDBtmPTEfLyeVR6CnTzLqR5ZIfkdUBBXTpfo
iw+pLfOefQCOxjWWbbFmwB+NIwv1FiFnvbgFLbQCTPN9YM3y6XQ47vjeqj864nHj
H0yiLdr9gBahdFVVQ/u5FiWiaTizxMzpx9NKvwVFWKLJwMZ8u7tBwkLeOXwGP9IC
vO8Cns02MstHrl6WE6bmY1weZmKAsZoRiPnLoDHeyUsP8silnEf/UNIVwhmIzHIY
nanOKm5Fkcsc/J3NMrmy7nyAGbdtGXh2EWety8Hg46N2dsjCX05jUVo/5TDEkgMg
HPhtzy2vlfQj1z6dA2KESykZQustQL70dKyxOSEi+G4MjDdfvHzEHuQUz3H4Sc4F
EpQ6ZEWL5i6XucB0Vu0mC9lPevxPcSjkgv5bI1MM66eNItOLWwLeEHm/988kgCDW
hl1+9VLo1Gdshu8+7TOcHLZwNTmfxHV+tC5emK6u/8s0pG6rESr3qXENdcaRulUB
dy4hhue5t7KUVCjk6qrD/+b6n+khAYgDcOlHJJrQ8AumcvRhAI1B4CMc3KiiYWEU
rU4M1sUPXeCZngJM1+gWcOBV1ysXeEfGZxJxW1jeLKIz/pn1xLGeHr1zCez/4BLz
V1Hbe//YbOqEB1Lw205bxCPla4D2ML/CZ7RikIICn3I8/4affIrZJ3jiHregBRnu
wzUb+1eo6Nei3Bsp35HCC9bKgS4cjzMng3VMMdaJfyPoElNZ0dKtrrClXLJkBjVK
otfdVRb4YgYEU5A1UwXyUkTBk4lU/4189igILB+bxRG1GioVyNa7ZrVuwIp5p3Zv
YACClQzWJhNAMll/NVLQH/IKnc1KMvnHxxW57aX3deZw1+dhNPMiI/d+YPs+Ej+u
peIMkKivcSw+DcVzpCQwjdqdml/UJv4Egoq1iwH/sSpD9S0aJ2q+AMAvOaVC2aI9
2i/I9TIo8WmUUsQc0UhuwP9FzLZIU5B0Di4ypQRTwMXMV8pPGtIbMxhtjgXdMJhH
75UlCi8qG16aONANE2oeYSKcyZIV83IQprt09gXEl3BlWsKx2tEtHMJToDA8cCbF
Y6S7ZAb2VRcJxvFbfdxIzivRiCIsRcYMQ6sJuX/qq/Jq+4RXLAcaoQyRvOQ24wED
rgULPC0oGcgA9ncW6hef4pC6xBMRi9hs9l+Nlia73+45t8dK94ALVmo5QGWIiYWN
3bjqkc3A4Z+8V9ML5PbWcK1ejg3XMsqNljmjzYUUP75dEB8x6krNMcKFtUr9Ot63
JqKapAM2H89dnUfEqh8GenQG4iZVaacQrQ+bzdFHv/nT6zzRGcCyZe7qjYza1Rzi
8U2hm6JQK56dDEhdtLeA7ANJovZ4Z1rNiOqn8A9fWOb0RZD52cJjqQkIqCTl4ZHS
m6Ry3D5UCDjNxBW/wkwcM7hiEFmSgJjYeQDLnHhROpvD7UG+8yGCqMpvBuP0wTl+
5Yq0WbO9N3aEniR19e8afYA91OCV7EvkDKISuW08JkCNIWNo4nsUgr5c6hz7tJn5
jEpKi6KKVr8zSJG7B/c4sWuW0lFDU2cZfadQ3RHQvAbpTsMdOLv/tQInRhhcD5gq
h06CflTBhUXbDfp2q5PDffr6cGN8LhnJxEx6tcYEd+AqQ/y2Co1ItpqptgcW49Iu
jkv97bXflNkmoDtoPOOxKr7PM+nTf0vWkbNxnHCsTtUXoJY4ENgPhIrA3VgKxpJN
K34qAB6sR3x/XJHNIACChiDO864KBiGXjK2wWaue/5PVgpcM2Bo8LOGeLENZi1vv
opu/jn4gSRwJgTnP65He3ZQv/5dcgcj48fh0XyWsYb0AnIcy+IU0olxm1Cfvc1Zh
FXdoqtHvo57dH4WXR/jiIAoxnLjBoleYYQQGwWBbFg6Pj/MyiUr7fdm13l3zXrSn
w/d1NB2N1lJGhLN261OCt2C0nE6dChpBqRjDoE3RF9IprnK8sP2jm6vs8mx06mu/
qzGUq2lo5RDVRQRmEmu3BBybbBZY+Sa9VgmK+s61i9rX6MG+TwUyzvqLbtB9Karf
Et6y16KrZCFf+eTF8xMo1LGpG/heexSM3saVHary5NFP1WcY9X4vOOtM1QCaAwoO
YVQ0t7AYe0Rd1vMfLSbFdaqgZ4HfHWrUPYmrtiJPVJsKVetgHev4Wixqs+xe8MMv
l3Qwx5/+roPOxl7KqIK3sA4/0LSeTQF8bQltKYQ7M98tluZs/xqQxRgpRqcrThtm
JVNcOTyyKGpOZTgQj+0Oc5QOFOTJv+RY1EKlQgXp969EBTDGzwoICyi1uIMDw61P
99eYJh1tS1p0dT+M131tSNu8KkIoPAZJOlraV9AckD2w25PUp9L8XCnSAwLVqvyl
kbvv3RtSpiNp/8Uu4LnThbLFTpJmmuE61lO3Ai3j4TPW8IsbWNdM1i3HcXiyFHm3
8whjcfEL4whsOFy6G37lFf50p1zVafiJ1Dy76QEs2/WE1MB3y6H9D2OqeagsXId8
urK13C+1KaJLrTiGvFJLIVUK36tP59EaPjzV2IzvCeTnHNwD3Xg9VK+nZ8xQMB+E
sO8uL9wZ2a6cNEV/vwNLCQnQVVMs4b5URk4qrvWoeteYS/fQbrUd3mB7Kby6w5sx
5aro9NKrXZWGdjJhu+WT5LFhZL7S9tFmgiwTXv8GZytAFqPIXXPz7qqIeQ9EqYME
n0oYtaqSxQfl+mY9cA+bTcfQilC4BweaX0L16abAMVnj4pffHGbbkmMo2iHFyKf4
DtMftD615n2hNivzdQ112EPJD4Gl8KsfLBuhzkr4ynJCoGphM9ZUjnazcoYcJACg
hmKI+LG6/DJ4iht0O1ab5dyQEa7xzk19TCpRH4T+UDkPkJPmgJfvaW9PXCyQZAM5
dnHhc2T1IPkDILhx7p9yJbiCk2bjSOBlIRVg7gLtLCP96PhXICXStISyduP0Xwd0
k99efFdEF51AIlqD6uy6W5+bbEhQYyRJV79yP1bM6rNSEbtq8neX6NH7ohLFsc4D
nxRu0gOfpy8VbQJmgwol4zTJyBb6yDXaAZgdNJ/93Rkd0EP8NssMCnsBSuv0kDKU
VCIrhbuFgltya62hA6dUtw9QSFN9XTieVm/0JDLnA7BubCZTJYvjsdXuaMUi26Gs
OOQSJOR0gTMNTDcjM1zbdLcSVMXJfZYAgV0aF9przOwxAqJtMlP9JClXG8Lv8PrP
xH7kvnnPwmL6PGb1k+PF8j6HyK//Fi+KK4uiQ3fZh2JIZAK72v9ttJl57sz3yhnM
iL58GSfIKdPmk/XwOYxBz3FUronxdyYnz2rER3nOL+MoCHmqoZ2smoGn3AKzdU+1
CkhdDASVWhNnjcu1lzpL+R42ER+cWxJxcuP7ifwY+6hhbxxOpwmq7T5LHOIXI+Q9
ZcAL865rD0JnbnOhRPgriCj+br7pBj/Jvbgwf6DEHnDw9tpdumzB0jHkEEekSs1c
ZegTips408yZS8InhxCBeobrt1CZPf7T2P+jPOX7MMBlaS9RzK4IewHtycx+K/7s
YPRgpItz8AP0yxUED1xgCw==
`protect END_PROTECTED

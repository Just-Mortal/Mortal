`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scoYDTkW9wfgvJOQstIcjwD3DY/E6fs2MkroUd+6iThSdgbCBVUPWslDqmHHjRZY
oSMvBnmMHbvxjQpQOLvFMkMlQuA3n67cRBm6rg97nvqOb6yghFuI62rGV2NFwOIr
8L+cjvgHjZvjlLSq/eHBSPZK9P36QpGGIxj2XUJGoOsv1BP7J8UTjC03w0+zLukR
DuPMfx4pbDWi27cgqLoa3q67sqg7iVb8GyEaS3nm+Tbcz5BfEstyL47jV50NG1c+
wzscviQo7z8S+suQgxzeyE0wM6TVA0jML8qCO7Ak+cAEK2DcmWH2RsJ3gyeYRh5u
mKSgrBP4sc5jgL5dwtWeNYYFpuAMIhszBA1Nf+58K5USFyY1yny0KzI4GhbVvP5U
KQp0749ktnTyPncxCvbNBTxs4xeVvHf91dhHvf1IxSsSSLzEqJHAfa71/F3oIzKP
OJWj49q+lii3Z/TGamCsV5eACYDHSA9jSYtfYJflG5ZjcsQKK1NzBpbyv07bhALn
9n1jMZRZTAb9ck2zjgH/kCVnwxrvBVACYzsEPT/evSiBE6VIqxLFmDF9IiPfec+/
b7eTapr+LB8SOJP71COre5eaYD/OvPM6t29Ew6RrwGyFUR0MEKhdmYqvXuHuSNTr
OdRdT/2Zw/hJrV7dvFHGYtuxzOtB1G7ZfeD8/LREUJGsrY6GOMm6ZPEqpYCbA+tA
ho+r83gjqurP06vR7UHnnVscsl3puCK858lla9uAP6TxG0g83nozV3hVvgwl3r/q
0dc/3iCkZ1J7413bBEoZTDn5pMHJH+GFuevk/ZqqFycGbYG3Y/gu193vWPsgeQRJ
iq8Nq3wQYUKoGAN/keJkMbMfNYrEceNZYbfis1HDChftKhw12JXl705dDbxvO+77
VaH4XPhiG41gclCl9a6xV+kuIfGOgmRbhqzMqe+lEM0JgOh4txAFW0S95ZEwXjOU
n/MAVuOthrbqJ612XTRzFoUW8632VN7cSoOgFP69peODkMCXNICSB1mcexxiu5Gs
ZekNRHu2xpHntS8IIctkC1VF/rq9HaQCEye3SaPyG5YJjPQ/NyBtQJRIv01tbTKs
/9JfGioM7ojmPO31YscX+2+KcfzLFvFzs+HYIzgDzUhI48VvDnsDVYmQeRaC3vfz
/u1VwEe3mays6iGoV7StAsp37rbi70kWxdV5JGP25MCcmIwNu/tFTJzcONHd3zhI
uQAcBltAZpt5nH+DtkSKgoa2ui47cQ3IRp5i0xJ2R/c=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8aGJoKGFC3UmgnmaQMTP1B0mtXjd0P+bxETWTunrNloTFgQ/3G5Mkc8aJp42nJg
4tnWBOXBkrJBD1tKRvawt+SuOQgsNSjtPE6fYTy16TxEQgDGCzIwthkdczTFMQdr
3F6RY1pFLnFa55nn6c73lPj8e3N0/O8F7SdBmiqDj9dv0zDFFs2POsTg94+/UZod
VZAiybWa/Tv1GgTahBcBp06PPGSY7I7o6QZjHiAmAlguefswaMPaEIPla0yV8Yt9
ItMcuimU+3CIl+WG/L6NEkPteUWYmNLLu1ILFYzi7EXG2bGSXgL010PZwAc8U7n2
tDOM3RbdQs7NQTundM7+e2ZzGVDZEk7KACj4GQ9CiE3HuDBol8l4JWxgt1dwgw0k
YouBci5n+mAWoIwmLiBYdoxndeWXKvgTX4AfhYqtgk9IUktFvOjwvjEIduHjeFHu
byg7s7BTVNA7jSIiArrIrbK0fUmWYMRBX1O7Gc8p4aVH31u6p1DYtPmyMEdwbrpI
PzRWHPq9uSfwS3rOQF3uGiblupG9bst73vMK3OGmg0S68oAcwZoBWHUq/ZvzGjxI
gZd1aTSIWdupQKgXmsa5+n47u9OIL7KkUFsGRh83Q06PViuXnCGJyrgIGerNSKbg
9f0cQzML/172AaSsGKij8rZgMteydMTCAb+GHJIgZ65AThRTxFwvQ9fpjKqWNoZf
Wvb+dGBfvH/Nl+lLoI5qtOfeeJxvJed6i22GjkJ3bI7wGU8VYltwSjzlkYJks1dW
iT9ZE2VDi7cXZmjRPx97dOvRJYU2CMdJ/EN7V+P5bW96Q7DCTSQgSB7185x5I8Gh
DktfSvl7MrZXYCij/iItT5QwYacwveFfx27OZ/JdaZv/15hJ/4A2dcu6PQlxlAGq
0RYKdLqW+ZI8cZvP1nUqfenznwMdsAQ/8oCizaK2JATGccaAhRSSZIFE7la8UB4H
8kODEchEDglFKOvDgJI1vuaLk56DLjPyPgCzHCBqpgzpIIC3sgkPlMq3v0GvWMh2
xFii+8WgyKrcqw9zlozvzX/+CqWWXA+ovqp+xnCBLGZ3CN+tvwmQ60c4S11Y1esq
rntxyaExV4oJLQijmcBR5vV0FuodA9F4bLq0369EK7gCaA9HlEK7d+wHc26akRa0
QyOhWJQOo/Hvh2wH9u06DESjZcQ6pf7RsV7uhAIv14Bds4EoKFn+VT1wtm/uSbUT
Ab8oEFHqT2JmYONDleNtR7ufxGVCEn4/5euwq6k1LTH+xvxn/H9QCGId7ytQ9q+Q
XTxWrXnNhLXHDkFY9sxMJAGFNeZciHA0lTjB1dX21fbrzRZOjPEFxEMvLhA88bvr
6XUKISrU0eRu0/vEG6kBem7rVCM6gXZFX0hjtkV770zGlkzRsXf8gDrPDuJjlH37
+skpj0t+aNAZ3ZYXXxaOQsitmxFu58VZf/Dus1PUheDbQbKKZjxsUe84Kv9R8tSQ
s1dNzQVwfT7cZjj2rGe3Yg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wjG8HP0Heoa1OgTn5C+haUnVyGmOtj6Czm5j5WsLYA38PTDD0PzCEfT/XXx6jlb
f/haeYWJEDMc1uUBWQ/9x5TND/Hj8L4ryI+EdASVm42k6VPiPOSopXQi3M4vs6ea
mYclOcax2iNzw+kkqKaEtGuG6UjWIAyjAjZLN0neV9giapw4O7uR0MFVw4o4/mLM
GSyU1epUUmUP0Hf7jZ9V+ulJcAu8+lYvmVw3+EXQrYlMM/Fwb2DNHREscstNr3rX
8t7VLYaPBxMYibUavqYh3pD36m3xw6kHKK7PtcVS29D2L93rWGkv1OtvahPh+GoF
5XLAI5PbkG3PA+rCOQGGoA4HbvPzKg1eX7SejmlybaEP+3mYIkw+TnJrWYd2m5rQ
/VC+7GecfG/z02wT/uZGIKPQ9GcJZRbbyNXWWrJh8E5dQwS2AVJebyqYB2VUksYf
S28NfbHINi40TCMlLE2k74wRqWdDq2/9wjFO+5pfuLWBs4wO8q5mCneqF39InrnD
sn7qMKPm7rGvbkVZ1THtnnG1UkVP4MuPKRKIISdP0RsQmXtejIEm1RTad6oj1huh
8Os6nmCZgEJZbRJCgE4zeVKcwF17a3WJZrcGyQRvpfZ6AEYB4egDF5e7/Z8+Ca0U
eYavFGHwNaUUITQQ0HzL6r8mYCDv0oL+wSN/9yn10cDbGk1SaonjEMTinuzXC9Eh
Jn0PKAIAN968jR4eq0tSUb96IqZTUXV3sVpk704oMkHqngKMCvCFICQblaJItxtZ
uRjMKGiF1rL3+w839u5qfJL2Jmbe80tlF+P/1iD0ET0LSY5x47JSpWaVHP6S/aUy
n9vGEYy2hss6U7MHTtLrBxIFzb/0D/xkG6OWiwEPb5jacBg4feSGZBH1Un6RHDLY
SbydlXveQK632N9fG9WsWm/OymdTKc5m0THUTEdJsIm0RNwzzt6nEh1vdyXfdEOV
Vy4Y6iuY61k5R14RqC1iQMzKBAlT6USWv5uHLdHWGxP96ABv25C6L7CLhLInd6Td
QY2/+kP25IZs9McAijr0256oNsZwief2qLsKG2+Wpi2QYIRSXuTwbrns91LK2kvl
dc15bWFTfMSnGbcyHgvtCO1J6x7bEUCntxUaQQXWPP2pG4akJnCf46dcC4hk/iCS
Zj/xIOPCzUdWgbmL/nM0TA6onjSsWKqM+io5UArlhnCEkODk8HxyYXar3n5kSO8h
QyoCuFdhGtty6+qc++x8jEr2U1yX3Gcyva63cJ3mvCquZxttcUWDy4623wA1bgUG
4Wib4L4lxVmnyuIznHj0ubrPUrIIAyxAaGEmJ3fgIoLFwaU3wwqVZQDH2nX8gDFu
37QPP2BANcWLfFSqcAi4msDr1ndNfUzQoN4hqariUUjhrK6lrL7jNtpCx8jF+1B1
Yli8mIi6e44hIzbbq51AbDbF6zsuKCx2miVXstbfSFMMPVzXkG7rXi3sZAmAamE/
Fw/v8DfDxhbjxeIUstowzosppLtHXdmZ8vWkZCCvHslW/p2F3/MPPxNUmzu4vgTG
PF6bOJENXOO8vUNzQexqYyOLYWrP9pbBye28WYpInZ94jl8t0KNLvzS67mVU7t+w
NhH+/2xPCk1Q/GPbqc/CYzdvsYRnQx/3CyzOU6xyA90lZKuR/yqD+qwfxZ8576xz
mEH97TfOzcJO4t5nN0+I/IrdQBiGzal0BszDWA+mJwknOiT7s6DpdYpHU0J/ylDo
5M0TihNkMSLNp1wQain3pUwdivKNlYQu/HKh1uQ58xF4YJeQk1yaT5RdFWwAFPB1
hq9JeI3ncXWUkPONz14du4GyWtJbFBFIqsNfERtnHpBYRvh+wQBZQtuqXokU8sX8
OODnlOdaouu5zJqTZ455UeXKLL0TwSXRkTmTsDua9MbSQspySXsv1IJcX45c2B69
n8snQvGIYmFaO2vHl759SjoeriT6C6C65QXWXfeu/vwZLXTsBIxqFkmGFDhXkLyp
4RaKq73ezYrAVrb5zM0q4PdOoIk98jKXK55twMkXqz0kiHEqtS13b3JyJaE6Q9fP
mSMyAPBS+9/+CJWkgphuTCf4ajAn4DzMEGUJ2PJeuC+NOK1+Os6Z437m3mwgTmMY
w+dKI36t+Jv3I8Njt6Y5jHLzIY54RInVDa+M8RuJ3GO61NQngxoObc53XQUvNLgS
bc5NsiTBjy8nqXHLb3wUnxDisL+7OefOQi7J4jpM3S7uDx2ZY7aNuCrbGXaCOFDT
U8rRdDUpsfYAb4eR8w58xgum6ZzoqW9Tge9/38KHt/srF7SAM3Btu/llub7f/u9c
AcsAED4mLCOzDSuVYSkZfQqakiQBe1ggpWQJoQL8HnJJ6ksU7X4o3lNlijWtOXXy
lhtCDumiFseUWSPQLOLNFSEkgzm8UoddQXHchJbu+XsXyXbJxXkiHYroEZ93bJj0
DWOHmHpiQoZDwm63bTTCFxRKF4PaXXIgHlBOcXGgK8s=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1sx/FlJuAWvsKxJjM/kFKpc13mbQDR8NcalbHSBwSmMdKShXPItOu3ytgCWtFRs
ZkDb6UKpdEP0vH3XoIeEpVyI73inh+8UI/QKjif5Px6uETRde4x+DC6T/x0YPxpz
/slwl28sPND3/NUgnmbQZdFOUnmtV0q9v9sNq9ji92++bB9e0uNlR42Aw80sXOue
AyJcJLgFO0hMF0Vmi/fNP4MhQlXH9xgMPk2tcrea/4aPKb+S2+/F5cUg+XO0dv2j
CGBLHWEjSE2zUQPjYur00r/2ux8B9JP5TSA4O1tCXY3VPQS1T+Ge560cMNkg2vcr
YMJ4GzXE8lkZU5obIZ0SuR+mSS5/COq35f7iNCpBsWP1DJCmSp+S6v1+lDkOKz2V
HkJ1Uz1NI/VBieLA+wvss4d7o1knvVmmcY/lsy8gtM5tISOUNVaVJrL48ONQi1gG
/N88znPeFQwhKgrmlZ+E412fKwGcJBQvrQeEeQmGHznV1NoqMzJupPTc2+vys4Lt
Pqv0t6X6AhNAgl/FfZ27wmv4OvDX76n28e8ZXNuG5ggl9BrbJ4DDLYJKblEid5xa
iwsHg68kES5Qd6UfztzxPDgo8RH9MhcQiIBdZ/zXIOYToq+V1jTtdYDqkm15DTK3
G/5RUgtgH2F1Q2oyZphJ4tjvfT/OO5Fd2dsMjd+7kR2aoGPbFgmFLviU63v4cZFa
uFeit7H9AYH4MksBZWrZPBfne32oiGVCoHG+l5prMfKaIbYimR10Sn5gJPFEI2E4
NiTyTVK4PNfFU1tkA4ETAr6zuVSxl9E9gNb1oWdsadYAgqZKR7Gr1OAtb8Dm7ya/
8hLpQn/CKJNCCgJvlJiXU6AaMLvD/9/Ub6UwufpTj9YLkAQ6/TWhmZXtixBenOOb
r04TrXkJr9j22nMaNsXbQqPE3BB8ZFlJD0HrKDmS2jk8YSBmeRGEU3162bhAGXMV
9zSk4bNps/zn9XJIapnqI2zHqRcaqlSDK2avOGQx2ZWZpnd/JwvlWc+oUBk/45PW
ej6u1EJyx+eOZPdRAJmfWn1vsbWdsH7T5TsZY5Jd/xgVOTWAcLJpLLFI2YrFgrci
GwdJs6zJ2YYYszDPbvdkVSvmo7Nbsny6uM/D5117agPYIReh3wqvJJ2AvhmOlY49
GMA1biH40v6L9OlWacK94aWrQFxRB4S9x2ks8lyrwFzDpkyFFe/Br3WX38FyKLdD
jCObBcwyl1MdRMElRxoJs3WeKPEmpUcBsMJw4LHKEjPYsjb8+kVwazssRaMtL1fm
RR9mNCq9i9PVWiAldXPtcSSUJ4ns0F2e1AXjMPeozmyHSAxXcQHsHGu+KfQB4I4S
24z2hxVYg7SIA3Bo8RdG9k8wSeSVSeCZvRHCHId5uAAYqDPH8xvtL6JE4LoqDOwN
uEId/oOnb9JrQS+O8IswKEuMSbfCmtj4gw8AyKpiqItZQK4HqMjFZLtAnsS/0aLZ
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SWCob1i+CzbG+zR3fbFos2zTlbcJuJKLbsgX6QSKZH4xliHGP/tmeTlc/5eWSE9M
lQNRX5gY9W0KjkqAIblmOhybo2Nx1dRGXKh6ZCS2fqzvJ+mx8OWgtXZuuv/BuKXB
XpJ30s5V/Q1LaYOTuTRctPYPmEm6NgwQ5XBeVpIIXl6RSrqpEL2J7jNe4Rexm3iC
XBQSKTywC2iCjFDN/lKhudFt1Sqf9rHMP2CwORRW74xzLDjJJ3OZ46F2by/cGWxs
H9lA1WLBeh0WXzVKRWyx36lf6JwDoquxBkvjzYkbkHAK6E4eaqHVd0nPChzgjcP/
pD9mptWJojAxVAuchGGYc5N+5zeT9+MJ/yool6TvUpD1AsaICkYwyAkf48JQuQlD
3nLRtWz6CRrESuSLqydnxgu/95XYzOc8Fr0h/iYOU4ulkGffG12NgtNdMTZ8l1u3
YvKCmv90yoVy/OKK1YquL4VRu3AqnZijzUu/VoOjZthv0Sbpg6byKc//iL3ziQOs
1nf89Apj2/cSh3AoRlGpdhTeFVKfviOEVae4zRwZsDuk6qT1FNJmX2VgdM9rsI+E
mcSR3IOISFeAEAkprNuMpYByrWPLN3a8+Vvers4nYhB6mnDZ2u0N4Oi/HJndJT4Y
1sFaeiQQtvguaa17C27m6YVSpcaHFzYc898VmslfiWnsDWGVUH0geSEYuNEBL/5b
35KnxUZrev2OMaLUIw3L9oC01WAkbsr2iqwvLsXrUh8XUeR/MfM6gZxk5/NtE7ub
BYqmCT6Dt1vpev/P+AhMAHC7a7gqUGryWPUmi4XeZtXeDmHxrDD37gqo9xcdUb49
QmGDdj2fl5EVJtoO8EZZGDARmv4H6ajbboKuNPM1D9eeV6haq7jNU+I5BxJ4X/bY
Pgx+65rMXjiLhbMVEc5Y1AWmEQOLXv3J0aBHtMdukGNxr6AWMHPSWUi32QDcmzy9
wOP5o4I6XM7Ly1yClbplvfDpcIMRRvZ9FHQOrJ5dL39DJqH//9fNp7Y7Tx8Uq6O+
cn2V1km2M9pUT9q5bn89ABGqQ8VTf2b7Z3Dfx6yJ53a40yBk2GmlDl00ZcF7dx8W
5DXTvKSdAgmM1tW7kDObv/czFxfwF1YZeOrImLEkQUsiA23F0ISlhQ0qlI3Vi/kr
VrZmCzfJwj+Amnvg1R4mj6ecTUk9DEBQ3fX9jVA/6Zwu7fi1OYmNnh66fzpCNBZT
J5+7DtAOe7oz3A7YjgmikWU8JPVW5l7Es0PeIPRh+gdvZwMIdvstbgXIWA23jnab
p/FV7/WUeeSPFkPK/4Rbz9GU4kFX4ICGrYeeECc1N26vU480x7SGAKDA3s+dtaAz
9Hqh6EHNq8T1rpppAHeugZNmQgwGLvqHb62N91i78WrEkdCgwvzKrIz0dbZq7/UD
ySrffmCYbZFcIWQsm/V7/OTK1T3YzAzsVXMvTqzLjpAlHEqLZfMBAdaJd8aO7viV
1aXBcPkONJq441wbXDPA3FACuJLyyG/p2/siioCxpx0GxV1LpXdQnb1m0K4tEkBG
aU64H8WtsJxC67ZIwG4rDiXtqNompwj2fA2WqY9x4X3YXJ4ErScCfsSwKibJkc8i
8mLa5L45i+Inz/Ii81QwliFOCP1Z4DiyfkXzEvYDRyXW0EFaJlwJPaegbiFjfB0j
nKYQ0JXnQcHf/dptkhKKn+6hwgANkScpST4lf8LzQ70+77d7A0b7gMOKpS4AZrgY
9uedg8Ea3/Ztzl4p0t5POpPpIftgcqZDr2RdSxfRvjc=
`protect END_PROTECTED

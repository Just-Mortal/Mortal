`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQ4lOQ1WZKzN5w+S2/91Vqj+yRuBroFmUh+UYweAubcDLEvchyPUKrpvif71wxjr
oIkKedJ+gPHIKy6wPh2RvD9xnJsrcdAjmKcmNfIcHQf8Z6XKlFLJLcIoUxXP/ZGb
U4C1ljXzaehtgbD22/9K9vnfhijG1LBlhRgZwg7wVgdoypGgPTwoijojHc7wCb89
oRx7Jp0z4CYjwUE/FhY7rUcEGSnRjjwcR2qr1+2rPswADa9DPP6wksfZkwoS7bw4
QG9RgXoxLNVM1KpumZhmT4oSSQLVolTE8PDXR6Qu3+7fH/hlHpCGMuiNB2AVgHOx
jfYl+Bl0WOA1Scun7gHlbjB+WkdFJpTG7CPVOfKoYMlMEhfNy9GcWUtqXj1RTk7/
3Q1TqebzPqTaA0Y903UzZ2Cal2ql2trLKp7yA69hCi97v8OYVeNyzy5WJcY39mFN
MQLp3CoyTi49bpXYfVGPoiNojUupsxcyDsYjhgSJ0qpR9foupd0J9gPi9CqWlGRu
ZGJyEysGtqkLpsiNTM823Jb0L58y9r87h7eLZXPt0PmlrtF5ZX/xTc9ROP52DV4B
kWpNGu12marJyowSe3oJTxmAEWfU+iD4QEBBCRj6OiTZOr8x8l8+rhVDhf9SpoxR
EFNeEp0juS0+HNi9z3aFRP7XgfmaAkit1P9wxJmue9WAgIzWbmMI2VtzqVaxG4Xo
ikomE/Dm5LnC3VXBUWLgXEpgIWAtaYhdmtexmD+K6shnRV0bVETD2S9ua+GWzOV2
HSwVr/C8QNmFoUmL5GhXp3yqIsDXqKB6+bNVE9ZRlDWRxyIdNVe5vLgG7SUcNGl2
cqbyudeGgCrCP2ZwMQN0exrAFiiM1iWzIriY2O/YNjOYySiSH+zSf1BRw5pdf1ey
FUHrR2FQQFiNgPR/wbUMx5kqhb3RBsHCHpIeHqAbkI3uzd0Otii4p0B4G/3C1MIe
`protect END_PROTECTED

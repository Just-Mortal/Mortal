`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vXCRJ8/igRbPX5G5G31RvYkgdpk9E3B6d6SMH6U+T8noJNbVcWRpWC3r/wIZSm3z
5kaHARi+0zIInEhtbMfIKmHK/SSzGMsYblDdCoQ3ilvxB3A+lzgg+1RgZ30CfU4R
Exr9pdUWCYNhf1FUAOosBK2d5wCjc8ikwGW2ae8xtK0Mr8qXNgdvxD3wRdtKfUcQ
YOytWP1jDlv/mXx8SEIGuJjzIJoYXE0+smvd0ZGG1RshmCjEqU6qFp3gX9DzWWYh
h2v12EhL4SNU+edqrTMNlHLuw9dXwba1Xk2j9uL3fBPzWpod34aylet3MzeOL1G/
+1ITnGJD1TdBWW3v5QeaTAXiYDt2U3QFfuNb1zTMXxzB9+QGMR8jDVbUcTshFFOm
HreN8mbKOlV2NzFii3r2RWeVC7S5GMPqIdsPY4hhBnfERLruE6VvNSG09p+k/BHd
fZEW60Ab9JT/so2/I3vX2MU3oyeoAlOuELKejIexpfgvimd8lfIDpuwR5N/Niysj
YfoDIxLE+55snf2vDhUp5vxDLkFpc/G2Z3ZCo6gxbKRrC1ORJ0wwDlNaYHD58K+X
7raH04XZ1KhD7NcoWZ+Dfsw0CFRoPXz/JYyCxpYho6OEvs3Ac2TEwgt/e2LFx3h0
53Q0U1inqdtDg6tAO6ZjKdU57AAnuLjOtbrD6tPEZAsLODoNBc0LR2swUdoRx8vE
6pEYyuEm74RKu5dhUOhDp4Zw1HWQB5p6stXnwSe60NjkDgZMv3Tyk3GNGxVAMrY6
wydTyvmAF+96jeRrQVd+iPuU3sn3WsHYA1g4+7ksdd1jCyh/+QUOHNz0vMOUJHCS
5yNpM5knam80LCJPZLK3j8b/xz4jpUInD0ahm0KdsCwl6HBV3jbW5md1S/T4n/Is
kJgomLWvDG5jcgqKO87f1mhxWJXZ67S/M5ZgBjLmDeyurMSjx84diqcpeVwBIOd3
2PV8/BrWrnzveaMiP6srbRHOB6hGuRi6MxM4clDKxxANzvhLEaAbUtwRglL4MsxD
Xf/EXBUgyuOZhJhgKe0g71HJ21kkvyhThdHKuSYPSrUZF1ssSwQNnFCPX8LK5He5
ZhrKUD8scQTD94lFYrfHorpe6INS83pFbjz4+lCyHWCv7aAveOK9Uuw4+2Iz1aOz
XlyDvPZ/7L2kUPOZOACtzdQbvpFA5OtyXzsHXLRO7OVoTzikj7fNX4v8dP8hs2xu
MeD7eNbp65fMWDJKjZ1lwPuQT2eLR+GiHo6u3CerCBOkZ0fWcklGKIEuyORvYdQd
ZXe91GAvL7wmvMTIcDWkr01zjcc9/P8j6ZCqvcvRe61QLbJHOKt5rBp/jsDFZPL7
PAmumkjJvXl6uNR9An7I3as1/nn2L8rEN+kwFDpYDcd3bM8je/OCgBIzE87e5EWl
NWw8j0CaDTbWoRHw/AtMwJCOWRtto/6LxVcYHjWGUr7vAQkCPbe+t0iTkAPfXaEM
v5J5dAISABLCCgH19QZLA2DqC9Svetjn5wM7QQ+jDNbGoRkvzac4cQnDwxH9+gWi
rvALPZ/bNDmK8Bd5L3LmA1Pmj6Zhywn33+wCLJAJPs+zQ72HbuDSTLvbUbVzelFs
kvIt1dDvcJ/bpQZ3VNRYm+dNEWq3oYChhgxQqd4TWzicyqnUs3RDJ5fMci9/xfjM
LaU4dpK+/NNPyl9mZKu247mip8mMMrdkDmOlwg9bMREvNzTWaI+0g2TDXF77z8zy
U/7QELoHatRyMDzBhEz3YKThAllgyNZeBkvaeEbAi1BKa5afHbC3JhGASjnI7yS4
WBGnkPy/mS+JpLSpUObrKg4XPCW3Wta8WFS67AbTCif9SrzmfxQKJ4fzyvmUfugv
L8WQCaINkN4WeKnH8NWTDIZOfRM9svtihytlRI3hwOTMFEY6Kpsd/dUEB6AgeWGX
glSh4oDXr8aqlZ0KHGmsj6XsH4QGfaaxTK0FWlEkbeIArs6JJXbEI8uCT1TmAyDM
GIuQ0bJROXQZyrSx8+MQdDx2Nr40qhno0CIwvqFTSG41YNZtB4RTtFlqDaVp9bka
2Z2Q/MRXwvejlDwJhS035kyYUXk3oOEIOhzxYQp/7+No72FpIy7HgDsrPeHqX+AQ
MCSUOH5Nf9Yf1OcCzheG0hxWDtxCYI9IqkFP+ag/5bPU5M0kD0wVXQxXJKmgAzeX
13HTyO1JvKlXt8eX6LiBy7zze+ZwyCiZfZBy6QxyAipJCux7h/IDXP7hOoCtUn0u
TIEIOaDWNVM5ybR+cAFDxN7zj5bJt4tZU9tcb8ocwd2cymY1j/qJ0WQiRHN5T4Mw
N6TxgkA2Lmk4xZteSuglBkR72PJGSJbPUu/iI5K+SIUTkbiNoCcRsOLoR9fpPls3
zYYidLU1lVmaIxw4/BfQTr1YYLU451s1Zg19fZ7it/d9T09hrlvxvfAzybb3jHta
sl/0RmcroxMJ+BwN/gnUKSxkbzUz3bQ7AVDvCSE/L854NKFjkdZjQm56qgKiyOXN
HXAy+EE3ult4fPpby7HcoQyDLjN7lXa7vPFhngobkK0iT/a3HnzcwXTvXVVdbX9O
kF02ObysDZbq1+zJXH10+q0ntNC0d9ZzmA9QT/r69vsNVZWarC98oVZ209Czc4nZ
uymsEuIa07UNrbT2fIcEytsEm6tXVQDBr5uN15AalXbD/+crN8IFX28hB4MU73tR
r1v6mlFUmQLHtliDLw0rolf3Q0MZQINkPxPP+H79gNmeu6/KJFLh5+h9Hw8xmkft
oaHBZj0BFEJiioxKe8NC0BlEbHhQ5BjjEt9hzR0yO2DwAWJ1WQc3N04QzhhsD76B
+PRaYRpYdBxPLE2Y/QAFjkpDt0tld6pAWNQNXkESrbFAgfSi60OaLqVM2fHDAlec
ukzQEngEEqIa/5w3mqxQTzX3jChaCAyExaERN2tPIDxD10CYyuFYqBRvc1ergcI5
n53u2g8mJ6Y13WnV3OGmDoenXe7BeKLYovQ0iD4A7ow9sytew73KQabb/PZVazlI
SbRXUtRsVzZ7YFLKtjRdjYtore+RYTHL6WTmvzkpe5c48aZr0KyAuL6etndBlCVL
D5mPvCSHARGXTnCaUW5/7fX5JPtN2FhBIq4oQfKoaAwI5WrBzCYmzlEddt+IPQr5
Mhmte0o5GLj0pJZxkyNw0LDJlK3rRgenmmeh+lHdZcB/1J7yhdC0QzMY7D8RetuP
9hCAHaIgQuWq9cPPjc5rDXlySOEWCcvTTh6YWHeubabIO7CQoz6hM+7SyC9cnUIo
VK4e54hIK3w8YwQqi5WWehQW+ccxrHbZYXSwkLsJb+eY1D+KNv6QCFRVIyxKQZAE
RsknsXaumioPXvOT/LPHIwgwTAB6pXZy3GoFeLQMbNszuUoeDQV56Di8XAQvbNiV
PUdrZfPM1toKv362wdyydJWvsfjjLj8NHehhUib6sLL0W4PhRkJAt6Zi11n585RJ
HZjzx8nxYwP9B482DR2RLNdqhhlbTjQ11/SkH4OLcMtNfOeCPO1dqxrjU3ffLOMJ
u24KKl1+IlpSLZUx6ByTmwnNwLL3aaFh2toE1fPRWV4LV1xeo+3kXlw7N2SsRCMn
jSQyIuDDdwyWvaThNHWZjHdVj9sFIT06osif+KLt3FufxYqbRP2C8IYxvlX1NcSF
RtoU3qOLgTGEfszhYiJtrCYbnrPdPMfqW0mbgek9wgNFbVKfuoYBdA3NVaHJISwq
NTkY/BEEfpXusdoABc/2+mKN27ed2Wh4oQHU62HU+wAeihMO6MkuTE33Cl0A8yem
gC/rocMfpfcUxoGpJK9ub4TTR4XL3npLg5YbIfwHEDe+LcieG3Y+8IHEVWnITO9/
8bpCM18l5zhVzVHoI5HAd7PmHwGbOiLnbRBx53e5zA9xxAQ5DsEDvBn2/68yRJVP
vnMgkJHqlaZTOQlDNJ++YwxqyvZDb9lCohXU6NrL1tsufa2DLwOpiiqVxjkzHvJr
06sxHUxOLmpaOfF3/qfrSHRXwK+fMrJRePgsF6x7Iq0VFXqfqocKHgwmj/w8P4j4
05ydymzS8TgefXuymhWAsnztUlPQiwbvNq7Mqst8XL8/6vk9K1mShh9ubFpWmW2m
C853HUepCJdq9UitPHi3Mazh+wLNTBsxj3VZoACZaCZ0BRlKxahdOIq3yEnEuD2d
HWmHiMJzx2XAipbN6qoawyWOzNi9thDWzlFqwl/1VmLYIuspRmnZqmxrRXBQRbFg
tMbOlaJZ9LeSWMKXSnJrM2plR/0XewuAPpFdT7viltShd/IME9Hue5LuZA5o62RD
iwjiu5i2fyZ9w3u6srOFSfO+Cx1YfRXksXnc7GqDbtDzJKngZl9R5XNGFQ/3mOnL
VEyVeVEEPzQmBFKlp0OuL29UWkcfHjq+HQvWce3zDcFykNxKGaxKZN4aVvFUC3XD
exI9MRAv+jL79b3zao/6FE7FuIjTf+Dkpo5bjHDh7sousnfDjrYO55ebm3CK9UNO
BKsWo0XYpfUqo8NJgnkYhQEL3kMUdVPF3Jh2V89mhkwvOOwqtKmMqeWhkHCUNT6e
wiS4Rz/n5sUTtMp+FHErcU1WE9Bu03btCErDwynFtIETCoybOsjMl4nuufIek4/4
kHJTXEtb+iSspHHNZk/PJGRVaZdgbVPr6CpifCwJ54cysOmKrI4w8Ut6LD7Fqjl6
L6GoKnNP4VShIeuXuzDQGpWFg3Bk+3ASdgysbcnFsuXg66G7ilb/47gsqT5Y/NtF
3gabLxNK5iRK4Glta0wFbcoNZyGnwQUhgW5AW7mpCLZ/dNfLn15qBoK68kprGvc8
shaglmVZNtMyPMBOnh1W02R2Ly5CdhTk0qhtKo6oXU7q/GSVM3qWHUNX8YfIMzLv
PBBtRc7BE1/0Anfcji9LMlp1zqf28ZUzDReGsvb26Ejk+GykPoxXxxu0T9B380q6
MMDKYeu3zV+vfOfxvRX13bm2bzJn7BhsZI6QmTi3H2tP+yekbZsnaWJAdUvuRjXs
d3f8Rgwz1Wpx6lQcjhCvr2N82BriAHnuPfSJYEx2LazuSqBI6oFg/NSTRP9Kp7j5
RMrIdIIOl2EXvorhdfpFkbN0W7DMklRgI13t/3xLcDwKKjOOpW7k9ji+EO1vpAlj
+zkpoTt6/mZaPniqNYzIf8Bab6RTrpzffVALG9iYSHYIUfeiCbcnaMeCCi5iPLAn
7cNRUvpmeYxipiOKHD9QMD8J9NvR+u7lo5NcBErU0xg8GrUfAxqR5RcvrJXHZwhq
/R5j8fe6/K7Y9xL6e7L7U77yWVBboaP6uDWx1m4SckxEMXKl7vG0ABE2n+oKdInH
jVmcZ7ErP7FEcTujJTfqFTQswvwPl1tsmAz7Nf9TzN5EgVM9pUIEJEHHvV3DIfB9
jGHc+MGPsrdu6UE53upE3DonPeIvj295eKCsGTNGQLDgF1i/8Y1H67CHAOWXYgWw
UXA7B9WyV5VlaR2c2n1ge6PFmUgLkqFhLpe4pPjDvSHeH2G/gNOgQVPbJMcJ7onX
dbzMlGEsOlWNqx0NsKGG0gLk1At5a3XiG9KOIRul13/aoHx3OacAAUp8cCu/ODl+
AGH4bwJoQQw7uSwJcaM0tOOMZ7qs9DIQkGLeH2ydAGDxI8W3FwbgWgbi2mmkRJqF
eiC/cN9r6fc0S0u5KCdqeWUTUwFuFdLjXqoEZB9G0B17XpVC5IMIzrMk7Nfq5VTY
X+rA1xETKLgOuKxAx6Ej+c+67JxvZG+QlFDu3i+BS91Fsqzs5iDtHPXGS1PZAECB
JcWH+DWLXlLMbpm4UXLkoWXpW4PmCGcJodoXzOXWPt1NUA8vKeT4TCV2IlK7QqP+
IH19pIjYYaplSdIRZN2jrjmmvI7Sa7zC47xoP/fjCUmMWhNVAl6b+YYGgMZBXQvt
z9SjcMC5sHXAURX2KD0xrHotaX9yrW1ix2nHGbe7XQJcVc3rZYTSfp2pA0SKpp1K
fer9GmPtn1RRRLYqFEVVPW5t99uStWFcxhULSBy3o9mlskFr61ylxECopQe4RIl5
mTvyrI8bWaF2VLVqBzeFkGlGxdfU3nzICOTXlSLSLj6jridT6XeXpWKEKn8a1zzd
4FxhdprmrXAvB1oSbqy/CZjQN+HBT0UsN5vPsvUkL6Rh0je2dpIP1DKnkXS2XLFZ
XiU0vhsFVKt9vmUKILUzVC+2PDokv5BdzmlkdhIVSbQVj3sXekr3l+BaD4B+p2BY
0UikKZyUx+zXXV9wHbBM9MyA2bQ757VHCIsUCYwBQIZvujjaYpt3TtbTD4YomfGh
9qs05aeq/txjmssjPdibWq/9Lt/s+4fviF8Ixi/JjrXfQjEWNNB1dFPYmTI4UOzE
PFj1YMhoqVvSj+QZqZp72mnkH0A8PB9Y6A/LjmEzSLN2fsY0ukDC1jZUct7wy1Ym
vh0mwB/sy6a29qeksN/iJSI42PX18kvS0wUEWXpVO1PMthDqvS5eZUguaL2hojaq
C/cXrYfIZfI+mOFakiJiQR+JkCaPPOyVvrxzFI93/T1gBbguEDFWS36dKKFTH1Ph
0X6Kw83bqoXgo8zjorG0X5tNQrDfanhgg+pL6Wp9up6D7FujwqmzcKjDWD/BKdCt
CT034IaGL+2raQh9o/DB8UqQWA/+nlgHzpbe2ojEpHGispjm0VtdUF6xnLjV23xp
ZaDDNRX9CkdVxjlciGcMzLI8JW5R+PKiqYqHp2KhE+swXJuySIqRKKGgHWbme0Am
6rDiwri4WV/Xb+CtTZKVqr8BigMnBycJwwimjDdP8H08WNjK7JJXDmav8pnFZ7dY
vuYbz323cSH5T9xMDijGFVLuMux8Y93NtZyMSbCRYp8Ke6p7CwJd0CNfHFBZMqjC
xvgEXpxx1fVHEDEpzg47uuxSe9cu4ZbU9ux0R6eAQfG5A48lbfMztOydsf5wLcr0
J8ueQemI2AWN7eJPGT3spob9uZMyHmJSAbODEHcdVvAeh+j8uLe6dOya+fmTaauM
09JP3kaXMR+74f9i520Gk32Wt4Dez4J3+PlvxB+sQPIDt6WbBqIp4YLXdDN9AOlY
R9p8skP/b/C9zrXUW2QAGPAPE4iChmWTgUZ6kIzot3w3758ySGanIy1YOak/CaTf
c5hrR8AaOEmVA5V2W9N82lMh1bzH2s1ddetjpjhvyYVm2HFtfHN80t2qQtDPJpqh
K3fkZsQHbYCp+lYJfvfn8lrgzrviCMyPeR2owShcYAeQq3rsYlUD15lgMAcyh5DR
KPCCqlH2cwHoSIjMK9KhU+SWJZ7rcBcG4wIWKM2hWnfFZcaF/PpJUIs0GS53OsbF
9n+67RH4cwVjC/ponTJuedIvZDxJKcey+X35aHLpz1KPg0+JKRF9T24QXphNL8w0
hpdWtkoYhPwjVvQ4ekPQbjBMgv9UqBxPbFf0sEBtFyni07kKcKn9VfqWB7r18Loa
m4oDxEuTL1FQOkve0txb1e+oIKgkPSREZdYrUUqWaFUC4WkDJtgayclE0HoaOE57
VpT37oGSFvlsW2APta79rz5QCyftqRYL/vuPFv69K7uS1aAE5K/5zsVk1eeOGJ2p
s3VOODMmI8Q7Cx1tP7g6OKDU5oCmfd81zY9VMRrzvTMW0EVLybf9626ZxyC27J4T
mQui5uxI3xOQwD/925JumWQRQ9fkO6I0EF9VwMwYwfbg8L+ydfwUDXoZpakUOO6o
an0I8Ql8JAE3azdmdLB60TYPJBXGoA3I1Raljs+Wu//0cKjVHO+ROVL5WYJKLpr4
lBjvVypym+gjxew8EvD5xRqucOr4RdDXnd0YxkSKrWdJLu6DXFznnqt/K9wvN6Vs
WkSXUZNguXq9kqyve5BZLvTNQye4ywZOPTz1bGeAdMrU6xmNWGP/L3JPh0aYaNET
TsU6T8TLjT01vhppYzdClwuNpe8kdAcqKGmoG3gKI5gT1A/K0CwXvE+28kCauHjt
LkcLKdgIJJxV6XerprczGC9CPgnB6iTxa/fMXqhBU+KpeizPjrj0R5/CLpSxFPMd
B3rZCO6LatVfoEprdGHxG1+K6xlf5YUV0Fs9fqd96SR1E717XnGPZLVzJjCyU2dE
bcacE8+T7Dq3yZ3CLg5DKJSRa6xc5aiky6x72MBv5GzAMc8Q0p5GvWo9dJy5SLnG
i42HOkIlzqFVJI0dJcbxoKPooVY8HgXzsGhMHafNoIbi3ePyMjdNn+AlszodFvYd
tqMUQWUGsfG5e8p5Ip7Sa1dwTEK1OOFh41KxUfKMqlAiufJtj25tWJVEsk0MSGT6
R/lq4Fg2mPAnZ55VmbrmneexcNlX3wxuFtmns3JI3oc2eAl5pNHmI+8xz71lO/y1
Lmj9uqlDhADd6Iizf+NP7VdAvGt1EyDB+ceIzfx1ha5U/HqJe6/PA4RyfUxZoAIv
bnB0aV6B3rfLyQijoShqtwXeyuOBijlgD+WIGKGeNARDYuVXvcEmV8j36MA8G+Xy
lg4oSUSa8FvRKVMI9CTmvC9GS7E71uoU+ye1bF5L2MjtLeNMfFVvGKtC749Vw0QN
GMc84E6F2fdeLtvJvyWZxai2lNfxElLs27PdKmx89JZIhkOBhlA5Z8bAYhG/U1Yo
mfyu4KFE8/k8A8opXf+wP9PCKoEZAFAWYjfbKaZWfc8L6vQoZm25bD5Vat9MkPrz
RvEEXHN6qQJklUgnl1uY+aYKoTJc2u1HT22hGdI3ihwMoUHSNJaeGIU8IVjoLT/J
Vo3UExEbf8Qjmy9evH/TrWFqZhx5sQtcta6d3O0r/hYvSFkXLO1D5MzOsqFvaiz1
mcnYym6LkZiZeGK2mm2cUEm070ioayGVAEoHA4VNF/QyWXaDyOICJtzjHCrkSqeX
l0UW/hQwxVEfC9+JOxIubzNGLNKqLD12OrvjqssrI4wszgtxfqUXlQHv9uUdIvvM
VpB2UgFkmAduCl7I/vLAv2wVGYD3dEmSxqmkNiCAUmsmUX7lqA3XkUmWccJ9H1O7
GW5lsvEnvPQh96XmO0dxxpIfOTwnhtIfvHDQDG8nRxxiG91k3wuy5DmLCHTE7zIh
ZfR7QpOBSsBatPZhuVFgUXuBL5KAriL28muuAjbosjz1MWFvzjM4PePckzOeMV0u
FjnGbBdMcvFnqaYuE5Mh3EmNyu7lR9+9/jrMAcppN9q69fdYctmaXeTanjIfCv7Y
3YnoUEQaJUTXfGBSpP9ifM2908CzHWddBNMhxY2iQWZ0jTmFhKCtRXgXANb2tYXr
P1Z3uH6ss3CLNFqVL7hWSyhC+FPKWe4zXIikxjPuTfNYrgWNqLcXER7OxjKGzw3d
FKGrGZeDqSOlQHOF8v6TjPzCUV7rsXsq4acvk6oOeytyAi/Wc8+jINvumSYAq72Q
Txl4VxU39HTwiTW0ySluoxOv3qlHaQi3NSPr63q6et47ez9qoHGrOyzOsRmhwNas
Qyqzh9VYfyKJTFWLleS/pby1uwNavh27vfMrgD7yutgh5GuCQ5WVpDa4OOzDyF6z
7afRl8i5TnsENm984Cz1Hs0vfkmrxSTwE4zoPe7H2KSO+a84QjsQNyRUgQBP0Nzy
ykzFMfU61CmCbR9BUF5VK9skns9oqm5nS/PLa98oPt6ZA1sbbPrmu3vvKljVYUQ2
MbcpD6bf8jiFUerGLqz4s8EzLxVNPJMS+drZHw0T0v4PrmTlqyDy0q1NEre1vAxk
ewf/igMD1GJfEp2qi2uLLle6Huha4Vh4zQEweoXcQ1EZoFnrN4dSscFMXRi6W33I
Xq11+rtmNVbYxFuubJDwWWRNEgYrMeHDtOiiuCGFslAMct6hBSIpQT2n16jLFjgB
5D2OKtZJa4EfJBuZvKHUNCVe/AefHLlk1VaTcmzAryOuJ28ebJCReDB4j140RXWq
91K82WW60UeTjMUKqMcRc18JUAY4ET647w55q7qkgkezaN8AiHsuBSMxHUn38i8g
Kj9lq+/0m4dsOz9sYG+ncjK8LdVOCLxPwrQMRZHnFSXnPkajCTALBVRw7phtlvc5
W6ggmoL6V6WWtHchyVuu8wpdPGUBiDHrGkLnurZD5bF3kHWe6h51NWQzP9sFg4qK
DEVvzt0mc8mgsfqx5wJA8S3aY1nXTvpzUTLuDbwWbmV2VwOCYB0eUXSjZWwVkDP4
fw+LGgyeWrETLgGxFCLCipL0dztv2WpkGwvIvbEgc6k/z+2ZaBhzQdEkELESLBgE
gL4BBOyzZHkWRR6cl6q9tO5CpVJPSz3P6Wgw9jI0uvHkJgAAROvWg/QIk/uWC1Jr
OWe1ibY6bjCkKvMAry5MxU3pP9o3PUR94/0gB7F5q3Xc5E87oDPa8Bj0BQErDWM2
CIJa+oCbenm1e2exPl6rxZV2T3+zJlA6CejEf0lcX3HtpQ2QCJLpij0DKC4OZshI
H6T67BMZImeFW2hfJbVS0RlCIRRZ7dY9X+MS1vmlWMg5cGzOh5P4GtWvg+DHWOr8
LfKHwwXFbyNdOpweNBZ9uyY9mmflbyAajmCYwm2sEocn22xKxGf5wBLyqxazxxzV
aLUeu7Wxdths3Je4fB+naL51nsZahY4Hspdm+9upv4f4JROPRfvKlPnxvWfbGXmu
zIHSmmcohlz88Fu4uPiiKUMKAY7R0Frsv4ERL0p36Z4DeNmOOMxodpDkXO72tFLT
bkHSRuLc+KHfYJcOxt5AgQltWqSlEz8bJ0tALZqtWABsav63x2E5okSKQtbXtWee
0+7bbfTgMM2wvqviAeoTyLzVWdeasCbn1XJD9RyaJYHdQiLIq86vfGpR7wXEq8Xt
PPiX++g+3/VTDBmNJoMcNkw0CcUPd+BPT3+PgFGn75oH8MbXBr4oTzbYGc4vBFXM
POGdgt9DK06wV5L5kXwLoC2C2MxcDAbNLEtnfMEP3pHLRHc807pk1hhWHBe+TJwF
FuWly5GjibOyxS8Sq3+8l3rHiKn72vNvL5WL2X2JY9Qla+prD/qJzWkU6UySnUqE
dlV6hiZ+bJTIz08dMUsb4uxKqupwmVdpk7p9jk2e80LcHGWCr/2TGmyS//D+zMRw
f1NTObvfdwHzcnCXrWnY9f959cDbChluFPB6veVtotnYuWfDtL+IKs92jBzVNmzE
a0Um5kTzsoAy1I4kA5mTGfUq6G7ACearIe0TMIpjHifBZ1xKGR1DTwTxs1jVS5qS
Ih3504W7WV4DBm6/byX5D+JNcok349eS35sVMtxqpBCyqdIDME5LqBrrdYAbhA76
524BURFOrODX//X1vFlbvH0E14xaGWUdCCFT+kVBN5qTHkMSfDKcgVOELmjC44HS
nNQ2SsCFVm3MY+13AaqXRAI3gPmKxJ6hZ4uxcRTC2yOFotYfGZ4V3Mwq3Oai3GT6
wb7I+NT1z7xaCm+QeXP3xO3BghYxamM1Spv5v+UXqMKQOwaSo32Eul4Et9jGIZC8
O2++IKgNbOOkh5naCP2dU2+YdIFHB7wDMDbHgmw7Lx914WmSZKnlg4uAiR0uzZVW
bufLNaBx63TMGww+mhGG0APsHMvUmfuHBbDXsGPa0Q+G9GLZKoRPWhN0TpMWsNq6
lSIxKHOZgwUy3zMM8/7O0gHPI8GpRvVrOFZng06hW8vNVw2U2KFIF5mkfPJ01faK
RbAvrR5Ehs9pO5XyVIDK1sWL535y8BoY5+buxi3fSQzyjYWbtMUDcPr2/3cZfK9+
SNWUDtv3TAtk1wZ/V3/XMYEBhzla6cy6evqIdMAcYAKKt1SvUwNyXlhEdAXPTYHZ
j0Lqkd47CVEEX7gQIGR0nj94jOuSc4rdfgnjTqRTegXKOms84Fxo5EwjKPyLbH4j
0oxwA1rRlfbZBfN4MXQPh8IiK4JM2cOG6XK7RuOdfuahLWIkCGFm5cyxuaPMMenm
n52sP3OMlTsjmjCzQbeXT9ynx06XdCn9VgIC3IWJYcSs+ts/maCgj2OHT5DIjgJz
QBNqDIF/GIkvATxODJJAMgxIKgJWTM/toBjgQqw7RuRdiCqiQWBtEc+mtvHExn4i
iSeTfBi2btzQNNONVHkt4IZLNdABW7lBOMTSaQIlvIscOQjApKMRcLSSi4YJqqlz
siGH0WlSocoFbQ1viWWQdLcy4Ve9WCWhu5NY9bnla/UJOvS4Lqcc/+77eaaP/xQt
Z0/tquz8yoOn8uO97shRQsQwDXxMwZCTM7kl6t0YVsMw32Cl86nlnmGBZrs2d0yJ
Csm1GDFS5A4U9A/bYU3NxSHttQ9l8dAgN//RqbUlEhQo56kevRklPsbEcvEEQOs2
g6f8cPL40DP3QqNQjuIonH+q6jJOYpbE4mImKrx5Rq1+mxJo6fBYn3u7coevmNTi
ZCwRHf/ouRdNjhVEknX97oG8fz6aiRdwrFsVo5VvIJKRoJnzG3rpVGgnGC3HsG9C
fX9vhgfSd5WhFu5Nt5sG7AIs80HORzHkOu7k2n9MQiK8LvVJLv8WuIFBEHDpon3f
hcheTgMeZY2zXQc631OjFfjkZz7MD8erHPncm9Eak54/KJrMNm/qCE9Gy3E222qy
SVEaXHCGanDCZRFJAEva0mUQG8Tgwfgs0eevOO/3w7O4ZgSDXUQ677eNfz3jQZOE
ZuZCA+cQ2dUzXmGbZYzpL1xCNO/SXZJ525DIaqSgGpqWzONzQdPMP+mTt4mMGxBV
iRtbNUwXLF5SGUQ4zvbXjVf4bZO2N870sq/G8XBSjDpeB7b+OpK7iJIDrCgwctWv
Uh4rvJHNwSbIIiHeEOBzw+p5HarVJvlZQyZtF8WzVeHKkJzoWR0Wqt087Uetph0H
VyXcx7gJ52JiunyUz8VikCyX2Mj6XJLDsOZuOHJtxgZn0MALX7sgesiHZ+Q/A9wh
VwLuaTmJZJL2HTEe8GZPF6VhfQSaxrPiWNF+q4MfJ+u1/Xs/5l0aE77PPLFxke+x
I3ouR8nrxWVzQyViB0CGj+M39sehNM7nTl4fzeRMiFxHJpbuSvRLjoLoCYC7201S
ouQPTNe/tOlORZZwq0hRECQfzx9y0gXxoXazcFA+nSuTiWMOSmq+vbfp1s6y39ji
5LiTwZVAA+BBUmH41ARBAJ4nijkk0J77zLuIhk2nmdxLjqQnvAo65+nmazx4uDZk
Gzk3BVm1jjBPK5ilCV2t0reX9OCgUY6Yti2yOeIfxNIrVlTdquBKZtrukAb/5RGi
ENb8BqZe0AAfJRL4pkz9BuZDNJzZkOUNQnKNeOmMFxqMscMHeGsQW5VXycpHpuKB
h9OlSzo+CRhG0txAupKiGCdqLzmet0Qwis1IY7A17RNIFtD8bEc2rUdYx/dyYllA
VKab001knX23nI/Z03wM236ipigB91PNNsS/3yKkbgMizxF0UvAVSvKfFXlr5WyK
+0xluetU9TIksQ1jkewwLF+Fi3b6z4yCFWIn71D/iUuOpnB36oI49GqmuhhRinoY
2HKUbls0Sr+FQlNcTRnu5NskenfPkacSrSQoyd776VE5WtDhvhvbZlhDTQXfHuN+
0lXB0D6XQqCkpW1nzyXxmtqGgdkA60DLy4t851MYi7iQjZamTzrQ5NKv2MtBY2g0
npfrAUjCjHMJiXjdOanHMhg5AA/UBucADgIJU3evkN84aDKI7kVGatgJiujKHoWt
pxlbJpnNgaeOeitD6j7rK7N2hIYfsOYRp/hIQUs+zxPQ/MyLcWMUVc+Fa0NYkOAi
h9/Lu/6ejDzxvmx7YDM4eNYQIOMMFnuTdLFQooFm6ATt6MVjmvkFGO7ifaK8cLk0
a4+h6OsjKsgLvVQG5tn+yf/NaKomN7aNCJoKxgMo6GjDarZPqARB4K7UAvxQw9Wh
Vd6SaOxr3lOoZe9fRGs24B/hNTQWJLXegcY0BhVgRBVpOq2J/GGkePP8oNv+lbR6
7poNb8MKznNNp3PjTr62VfEYrjKAdTlOebjgxHSkufcbqOK9N6cXyRYcrL6am6h7
15zpbHm/a7qQFK/MJ7OCmAm4VMs8sAjzF1lNOPfyeEmOZKy1F/Sr9PpbOHAxDFqO
9ffFPiSAzvdKdclIlm45rug0h7bJ0aPMScGC/wKKRsGEoPRUjxED8Nz4zp2sAJTG
6XjEbDrz106Z1zINN9y/NMK73atFLunyv3zZ1zyDyJj3RRn0fTrYEYx78Wt9lxis
/CcQdJXQCywZGcWWH9e3WARQVhRz2W3QcypGdCWIjFEgASbGsgpBvPKOP9RlxOya
XOlQUbs4RZixrCLcuoJA058dlxyS/h/ZxUHvzB+K+Ri7MmTrV2kzjOjZAjtOhZ5Y
CKwqP56bJRmrYPcqh++Qb95nt+2yUhgio0GTR8C4g+mOibr9DvnucvXSamggx1qY
0XULodwGoAWJFDZEaENb/JkD+GYsAffXYb+W7M3t2nTysgWHA6EC7HSaNOqeEikK
nKoJE3aDHnf7j/nxGIDFljuD8e43F98rpYcpT4kgVnsUbxOzN/aYSaKppXmi2Ox2
bQNwKqlTUT9FqW/5w3CWxjOwJyWjKoRgGzga7+kcPgWkqmiFPNs8We0cCuNvDmJo
DNQkw4cuXshGEH6p61TSJtodN9UQxLsoxrF1sNAjSR+o2F+cb7HjaMigCMLKQkqF
FIQw5EA7O5kPusP4kEOe0nA6wCEFWiOEar2W2pTeB9dp1wtAUgMNYuBPXY8ZT9Nh
9mlgDXcVyDbs/94gpYkcVkfK7UHSxhyYEi+z2QN74Yeqz15VCAClphXm6nvguRYa
jIVrfsfCxeU7lBnCT2H2JEvkVqqRX4A/46DON9/xBYNglJ6sA2O2LGf117MEE6GS
Nw2yUZQt7fZDYYaYc1RFRk3Dh30a+74Ekx5140jjJ9aQP7nsY4Z6gFWoUyHomYNb
iAEbjI7j5Wjz38nO+QBXYedAH7g4KbjMdlYgWyWQaWWM1IDjLCCovKCArUoXFuqE
ntRXllgDmbxbdHyqMxNelphuODSL3qnZmteViihKShjz9/cCXAyWjcdAes1NnJNb
rdEHzs2Yr6fJSv7q/fRtOF3tiVQt2awoS1egVh4Bbnj4frHTFCkWv/LRQgO2QYJU
OY+H+t6qVJ/plYRB9HGRMPVTQKHCrVCw786ixgXyKXQNFlvO8YDsIaS7HULiHIuV
JHw5LJAUQFapPAvXT4L/XVRlaSmTIbP6PVvpMhfUtbjXuv040tpKymSPt8j+tNz9
tuh+beMEGBtx++CsSLg+QHV3VDApZNEtAzNYMDJiQ6PrLzLlXjzD1cCxzaxmoT8O
cgwS8m0kGpPq5mUFWN8CFCF4Xl9dIZT74BBtG7S8EfDoeWMGHWex5frt/WbQw5Aq
N0yQ2GE4Zk1oG8A+mtff/1IxuGu24do4433KTH3KjGV5YJOeXopRz+YPx6EP/fyi
aTLmuV90pzaFU0Pf0jm1oKWKs7tS18a32dlRdQ2tsh/uYTGS6o7eOG895hkF0AK4
MB8jaxOyEq90y2w7M+2A2gpoXbhpBiBSg81OY9fLMfQUqxfcj9EuyBQGsW9iNcP2
kVma7rbRpoooFHSnHCYHI3U+ViniTXaQVBdzCfGdqAnfbaXv5J5JHlkbq0xEbcip
PeW+W4uNl4GLpyvOlKiMUQhamw1K/fpnGEnkFfQ4J516TNn1Y/laRyO2pNe6urRr
of1HZC87YUJf3ZDkwQb6bNFDo8YqM4yxTtUVeG5FL/HJOBxel/24zo1YuK8w+gqs
EWlZfIxZmsP0sGi+Ubgwfwle6UbDkNlsC9beQDlUdLnvnAu1oIwaCR0ZBVVWpjUL
uCJsLZHPNBL/2GXlOL2sdb9yJRXl/CoxYz5oXx5yLnqgemxeM5v1UDL9ayGxzwwA
xyqZ6xBFVTn0sQKLmnhaRjMVkeZp7XKbx0n2yo93+eYnocIosbRlQdijG2TapuCz
GZwlThtVaDna1k0Rx5i30k7bwAB7GhPlfZibsHJ9qc57ZIBo6gHrmiYG8EkMktC9
Ig5Y2jA/NmIxUZM37KhqmJ6vd91gMgWw8sO1q56luRaQbGgrvCbbPPaqti8S+C7j
4OYGgrKxKkziawlwMf8obMEHYtyJcNQQEQ2BwoMQKyxZB2RuSEb+oySZkAWBIwvf
LnLqUeLqf8qGtxcqEs5+rbwaVH837bLJFd+uThxm90xs16YRDRQuH7OPjY+SAHBT
82nV1cnyQAmlyBZqjkwfi/kPzpgoaM1Tt2AKzHYR+3UDra/nLhoZhMdeqWEk3cyq
NTTN7K3luqwXvUm19Qjy4smTgdtBNbQ862Xf//cCMEXl9tCdmoRea3/Vof1PjDVS
Od18cbcJ4xQiKH2ygPLJwdpl4+DB7uaWN/hVFYslSm9pDyviOY4+Q8j4xT68ouii
U+4u9zBJdyGiW1YrFG8GgnmoU9rs4rMnmoIl7QqzS+qCRYaMyiM9+dBgdzwWIHBh
k8IJy8CvMbQe9c2kWOSocazYsfJdc1x0BAmgyURiuFubJoJ5T6uma7HFCQs7Oa/A
/zNo19tCXSo9eoIejmxJoXDb5kfkyMg2AiE6mUlPccMM9vcW20b6atkPRwRws0kz
cYa0dJTNXKv/jaS/Twp1HWT19GNmoqhjWcli3kUjPEwMenaBNVqNu88/Fl9htE8r
WdrVwxKFT+rousVvc5zrPiMwmFQ5ka4qGrzr88VTx00dTVovEegsMWnZDPF4g2Zg
BNfMGibPZZI7B0tmgLvKFCwzI1VWj8JFdo90xLJGjdEXh91+QqRIyk9rIBjdSXL0
U8hMXKVUcdPEEg1xQ4V+Egqwtmy/aVKPgFVnJLv8tfzSlgwIrGhRRTpjvkTP06rx
ijqBpbXLbi79q6XNMNPCSqADVduPDwECLKu0ceSf8jSwekHGQES6JurwcivY6qdY
RKHtdWVX7SJcn4Z7JRZE2nzb0WIyJDiHP+AFDuIMP6m2wxD0z9p1viTstAY2y644
bcY6x/Rl3gNfv8sCBJpV/2dmdyY9JbqKOL4vAFFKIUM8c84bCSUaYv5ncpJu205e
anldyuMxetLte225HSV0uZ8J8FroLI4DcuMePirvhV+qP+K75itv686F/RMSfy9C
a4/UEH/g1+eG3S4pNuI+Fb/peYozV8o39TpOufhdBecJwxKNjI+38QZwV3f/qv9S
4j8/2idpWXOcn7/zbWv1B7DWyeb46e4gVUsgSmMKafChuwJHZwaj4MbFQ3weYk7k
ID20qPd2B4qMqujLUNLaObycXxK9q1uaUlFFhnhiRj+bhi0keWSkejAV1OYAqju+
oeRv8mznMUTtRGJPx0ZTncv+U4nCGElQrg7tnKAgExZELvx7sJA2vwq1Gj/Dlb1S
qPx5iI8Ef97Q1VzfNK5akTTKJdfmJu8AO5w/pW/LQ8tLwZ6aQ2jNGsrg94OBZoGp
VdX3xHVwqXBmsQFQW+sedDjS7Rj+k3Xpok24Dv/hEC71uMw328KMNL9hMINP58f1
f3KVj/3T+tYnRS+I6h1O63LjPNmrDx+jBYxQM2RHNd5zGDsJaA/QinFXqD8fQxPA
wt4zk/Z6DbReEWNYvgxfMM0F1GSBon91GJ7RYTrQRSbeL82in803HtEeQK7/v7Jf
4Olu+q2cKuAnY2OdNlPPpRKcm9cbV033EHW768MhaspS3/2dEsJVqXmy6Ld+qlnN
1rpEKi4pA4tLbtrGHAVMBdYEp19lBrX83g3J61hXkCovWvEzi03Mwb7sdmIjT2U8
Bfv8H13ZCOxWHpUuDR3PETPDTHzx3bTaT+3dx3DZg4d8EzyAL0h4oCja7Mthbnfj
kiB7Vmk8iDxYbR1ARFPTPfTg0DLiMhNPX4BoPz6wp6dRhIVbMXy91obK3XayE4A1
audvmELmAeAbHBTMc/7g90HLf2Wunh6Slrn/e26TyZzreJ4s4lIq5vVOS+2JnSro
zTIFBEpuWQwxarZFf+XKYl8A0P5JgYSpZYjg0+10QUBJZWb8P6PlTAa1H0oV+DNy
vo5G84/ZS06p2jjo3nYt09e4/B1z5ikFjsvDl0M4r8M1eTnLU3Mc8l/uDqhf48Jk
6nuloSNpney4C1+A+Klxc9d4+qiFhs2buJtwuotdM4pZPSADpyru2MoU2nRRxYiS
E+MuYlnc/htFgS/JZ4sEg5sUkgKW0EONirqSBm5SsjbGXt9zqkr9+PwK9Uld71GQ
XPjyfFEXy6MRaXGjraoaamdibA0L//7dy9Tdn4EVckE4A8/zsJXwe7yCNtgM/xdi
8Zed4AQI5hF3gEfbLfFMqcyZIrPcu3eZyStGgDO7BI5MMSHm9W4nlLVgE4nHoLR/
BVDZLrWCj4W+F/DkXmkfXZl7Gna8H7h0Lx1SGGIdoQvNqxkqeMjZOWtp3CnbI1/E
i8Qcm3xhh35LfIruXbU9xUmTmSBLFNQmSwJJdLeeTvUZatuPnfhCIx+a54VbzHWp
A+GFfIPLVvA0dOHsuV5rjrAP2PT+vT6it+80X2HKrj5CUK2SchI0fCPrac3la385
tI6GRLZ8btmvJZPbY80aJIP+b8nUcsPR6s1SxH6571ekDR3XbB79wPb1134oFSqj
6g6wtMP+zfx/IRRVHkiQZ+VacmvJBMYyVNtdAhPHflODJIH0p4oLlGvnaVwortLS
X+0IX/mk/JpH0o7saCmx9K6PgyZHoJxclbziETcyvTtGIZQSilLoEowwzlFBuT35
pHzXXgxLAQICL9YoT3iv3IOLQY7Smk4rgR2B1ydjmOEF3j6h0kmqXlpRDxPpYsKJ
havqp6hkXQToghjEykr/ViKDW9c1LXWpb6z5ruLN1FPUjBB/D5tPVGYJAg+irq+q
7fZagx2+Fn9TTmXYjEAuf91a9RHByLBEPCJvhQYnikKqdqp9vhnssi21oD/OBFjU
SXagJlXm5y0U4c0NbD1E/wlzueTBSPcoADyHxHkX0GlxNZKz5Oe6fFnVumCOcLmQ
X8f3yZfg9GsFtV6VUxfmL8jFnGMNJ7miCwJyEMrkv52dZ57BQQeAjuuHS01smpW5
9+ap98O02iXJOsj5bQUhvFH2toU7VaZBsSpWgPpe2Yn4Szgv4Q376McbzSzZjNxD
GNm9XfcIfL9p41aRI/ehF4zg+7trJGlYy5g31PdSrIwy/O5q/iBtgloCg7GrJ8MY
kaEzzXP0PrF3d+iRqvyWF3WqcDJMMlPglxvV+CxgVjoQa8NOB7XiNTyiZ+aa/Ffk
AbXAWv3I8augwZfsE27cRkRUbWzfxIAheEU7ZnzZufSaMowgoFVd+qZROV4YHZK6
Wb/4VroiCrJmvX7otv/wje66VUcpsQ93ZwRKlRJkMW0PTC5lWw+MJ+dqQEh37kzi
7y+cf1lAxaMSFb3sTO63/oD9801lOUiDwpnktqnZPDBgaQGK16YmSIz/vXxLs3UL
tOB074ExUx9FQqRKvssPZvAypZvS6y9OPDutApieWSjoIYfSLUuDwq7FQfdadBES
5lHGiOqCgdeeBfShgNcGXngnJh9VeeKPR9g/+9+b80v5/LiyNTFz3R4dJOaD7Viq
ZeK972+52JwCpGlW360E5ODY7JJYIOtDhwthLBW8zpjCWhMyNKrjSsWpgMPOeamk
ugGbXPrXYxHrAR7/Wm2c/7lYQqAOoybs+bR3ZSPci+2PbpGj2ckqygix2xIv3Jx6
J/Jt4tjL85ZedigSqrJsh61UwxtOlBgqsw+Fh/V0pRAFkWBVidGNtNzLVFGhwaQw
PeSsFMNKKUmSv2brdgT47Q6bkIQyN3kGIHUvOO3Qj587GSfmbHIKIlRu/3xnf1UM
hnFQprtyag2Z7hRnmo23UupbXx8wAshIBEFdkejKs6ro3tZuip0Qq/nPtnya7tvo
+NyJf3TG2N7WoBMynY0MI7MUnGkIIoqJqyiBYlHAGzVPow1wRkJwxUPxk0ejxGjk
sZGrHY/BBq6ygAfcv3tWmw42iVPu6Y/qk9xjPF5BkOLaBIr7YEsXKV2oaS4BoD4K
Q4kpL1/OylF8q/GqRdGol/nlrEjtUhA7R6Y7ZH5S25CGf/gxKSiG4xlt6c3CHKmF
d558kMPQcFP8Bu1Ew3GgI+M0QTZ5R32+q/lY6V2TAfte8BhiYEIqIr206uxNM5gZ
+u6VFQ2WpmhWSGe2g6mB++jJYsD9toESp4Que959WWZPgTkWRoEfPzuI8Ug4YhAf
5RwPwHpL9VJhXOYCxQ7vlW7UIZjqlsXGB0Qq56DEVtDDeVGrsUr4RPkZZH0t2/KL
GHqPkLp5RPiOu52ZXN9E4piWWkhVS2AcjmvsZxpAoeKqiN+Gc1rJ2nSisKtgi8+B
Fw1436mz7n/xx8OC46b/XTHEQiGBSdHX2TdDHSWTUmkOxIJ3zef+jKNDQDKg+OVY
qdmbLiuLYuOicUnnZVL4AsfQ+RLSLVIQrIIVRGmNbL3uu0gpTEmWy/BuvK3FNGl7
JQgdv/GG6EVKxvNzDBY8GLbdv7sk6DWvBm8IFOo1ErGvELlLCqPNfCx3himNSk1m
Tf4cIv4p42cP4tUfgsADB2eosCBfS1JyDRgn1ttoU93tCIZ9KFlDPiRGb1/wHBAq
L1CFJG5QKX/23mdxnq7/jFz4wvbIQBvrTvvaMPqRtEvsp5t+YxfM5lAx+lb4TMZy
Qn2E1amZMYQ/epdfudFClTW0V1iRINFA19lm4eKAdGoxGmvkufyChW6d1Zzb88v2
V7loDkLRQAp7f2xuThOv/1MHJj+y5tVKHPaIDCiIy7Y4haeiAEwOk1IVJsZcf8EJ
E3M90b5uRzX63hzUM0Tn+GvcADlhwCLvRzQJV3LuN0Q3HrqLHwc5zDYDutMan60y
J+HYVSYEPrj8ei1zLd2a9TRrtzm5r+KJCZ23VwGUNx/1e65XWekZ8Eh+qqAtueCs
gNh/v5KfjQE/PmlxlKSQoaDjl3c2Zz3pPOI1eMYIbXGQ+xwcUxcU4vlZS+lbbK5G
53ZVsZcXuTvY4KH0XiUmSYQwHN8zNrzk+Xed0h8vCdSENat6uhR2W539bMQ2Enoc
N8T9BjNHEf5t6VmJN7Nld54RKSljKoGwJINWDvCvESxnQ2hO2ftI8ePxE2oXNv4w
2vxK7mNeKWZoOWPYoLfCXzkicvOOyxiKYp3mxT6lKWQEY0vYsEmaCv/fWtMsjxeP
4lzuzZcTfYbZysok/d0lsbFKsTo9e3yi6dZBI6sIhxUH/eCQtNHuKjSHnE4JChIE
KYf6fSDDBjVMerjoYNeedLqPmWw77Ng1l6KzXdbRxK+RLJWpNynVYh5pDengMisU
qJ5NznZ0skVI2fZqQ+/i04bJBUZMGv8/oQwrsANfZxOfyHGGhtvEEv6i15GRZKIq
42iVb0Uqgf7YjuhiX62qijHPcICrIrO1plGRmabE1T76lCaT/R3jj+e0+lknP2IT
QknGeKxdqUgk04vCnb38qfEn6D3HOmaypav3ezAI5t4jD0ilL/i6GyjVZGS0ttos
c2fA/xY7qXC2KVMVi3P+qVaxtdnWp3DAR69fxRtbYXU4QAhw9fUxdg5ChjodV8gR
NbzuSwmamOU/yEGqMHwFvMgyPCqmrBvVtfMxtSRqa7n0yMsR11TgwC8UriXdyK0B
luVtjF/DkAanvhDRxXKXsG3kw6VWlmXtTVO7XPS2ZXuiCHXZuVrd2fqbZVn/+OWy
ooaAYucdolEJa3Gi/5VJT+C+jlFP8N8v2qXKPWx8hrWPAB/WxZMM6aRs0jr/+bl1
F1NOXz3BWuHnKioF8x7VY/dvhAMU3hwv+GXmOgwXgrSRKKAhpnCOkscNM8ysBwY4
dzqAMEua7oo6dkQ3Y7g4TUx9BcciYhtqgoLSXx8dVeRhscoulZt78DSUubCbH1T1
txaSKjvj3z6PKkrNiW7oQlUfVzKWcc7ejESm5UOmkSFSeUnNeFQn9Bb4I78VBjq0
FOVMsUk+JbX9sjVU4F2Z9V5d+7SNhl2M1oCipf3foczPOYc2K+JbRRw1q24t2MsC
Zt6T9ohSxoXVpQQFyd0A72ewQf+sjIyYUCKqi6G2bOGRYiX/eiEaEHJs8twC+r1a
Dgbfl05CFSCYbTF3nickjAU+RfOgnii9N0PjvZh2Tu+Ay3AtI6jC0S8KYXRqnqmY
Bui7AmmMleD5dMStyCwZyvT05mDPV24mlrRWX9R+Bg7yo5e+KNx666PLO2oZNlRY
ie2yWgK4N53l1/5ZEpN6amn0Dky4+V+YrOl2aDghkPi0R4D4t0fxEztCAU1kshCE
pNk16x6PHdnp766greyxYhEC6qZEiVLkroUFTcV1UApOrrx1GU7UfgZNlimrn9e+
yFZNSln7P5yhkZ19EA34wt9ac+O3oxv52owYUuN7CRouWdMRLz31G0K6kgURLgQE
K2dqlH7F8JCz/FULqMbxIMGyKTwM013M0sz2X75WYI33THPbxdjiUPy8Y6HVl33B
DmHrVkO3qk/d2B/r0l/e80OkzK3gohc9W3zDSNzd+yJf4KRgMlXpzeZF81VZcgPs
IPxXog3h/MZcpauApBHgXxkBaiy34qWbahW+kuyi6BCYT6R0/xE25s6p3Tl/8Q8C
gUISAutYMKqkP8+g7jmBG8VTZ0zMp08mvPvOS9tJsTnz94HSOv5IV5FoCtSEzbQ0
B5tzH5mBQggYPq3PveERCDwaX8OZM2yqWhXiPuNw9fTP86bYraZel1j1mv8D8vK9
98t4ucg2FahwYR3wmsZG8zr4clTiMl7q6LdnO0yUCC0itUA3bZf4BhOT57q15xa+
9IDPjQRwT/9V1PU09M4MpWtsqgCQFfrtejFFSKXmkMbRgVWp0MmXqZt0tGuRoz8M
gZz+1d474sPgukYDU+TqE9P9T6dBCe3atsC1AZnKFLTao4DLX9yaxBuMyQ/oiHFp
bhsjTyYQPSKMIufTVzMohSY9ieuPwsnrWMm0WI/KM6N/q7O2sLKGMR3SHDn5jNca
Y6iJdUSLZeXCT65aVD+bpb2Km67dPEIVXIgVA/+uAdOJZHlZDv/HuwixD4GSP8Jq
YtN0nNpiptxYfFKcgFDLH05i4kWLBrlU5CD4Gon4oiyChyCyPkyPJp/OtSsk74fF
FXLtQNHbXFcV764t/7mHh/DgcmUKd8VE0dXSUPWbPeEAz5yie0pTkI4MFczRRpxi
/3FEs8lmpEwUpB3wYVBuU9KX+Vk/REFbtqyRpHOPmXEYDUeVRZhl8WYu7ULTnI1E
Ule8ND9UWcgXC8fATcG8YzsAXxzOs/v1HXxIJasTpIluIH4cMLWEWpjvUjCYVAjb
I0Cflk7MykYFaAyLoRC9jU1NDnKFkBl1yqGH3rgOxHyK+mXlm3goEEXEeeKpHZ4W
bZ8fQ31zBreXz7bdJaiR7SqkU6PgHUOKYwpMNUMBJc56TX5WdIdm7T1Q3dwvx3LC
tqqulxOc5fEaw2+CM4AaHulhM59Okz02Q8/npWDN2JMgbTBbKI7nJ+S1scOxe12O
m+mdsKmsASS5hjzj8nzPKIDRYUmQ5H6nRvNzbhynErj0rzMUGVxdeNb/6yRJIjOw
Zgo+swxpXU6yiC9lvKq+6arcopP8P59usqj2kqA0yemmfvAGVqMbr+cEnxF1dHhS
tD37U9JXs84Twsc5Xrsx6V0zUmTHVV8no/oZEcn6He8gFDMuiQRpFZBslGUXCLWQ
jRM37n4YukaNRYW/Imog/fraG7o4LZkuxM1TsgBOo4yYvKp0vr6CGCl3xsVp94dy
/5W7IV0NUyVJKUGn6heT4jvu69AAetwWQdDj+FIKTwgjqaSXdOeiKZ3QExstunoC
UbBVjUka1S5h+zxma2bxG5NHMabZU5jOFKSwzeMKdPb0gI6thcQOCRaUlrbQ6bOF
jjthLYArA6LamnisKEFP8rnUJDCE0Vjd27VzY3eFGGNybIKQSZOImoQ/hqPwbXg5
KzOm9jKrGjDKCVp1KjiVZVEOWaOuisz0H2iL+RWB49pvAFXiEMvEIZ3HdFfB3O2S
7z5YwB/DvuCS6/SWs+liLJxCXXuSidMkIvMnJvPBdtg9jgHISXrLr5y9uoPrKMrR
Lq8rZxPTAMd51dHaTLDqXePLo79xN3nKAQCx7rd+FZUr6lR3tOi9h1aaEb6r/QK+
mUy75ytO5L3UpJ8VWwfwlv/tiT6QnxOnRvLwaMGyyxx0mSvMN1LZf0H8Ue38h30f
RBWrICFWfoipN9Ze9cQVMHMG+dKQHEJ4zjr8o2xRp1JHAHMKfTq8TC3KvQq6LHKn
Oy8wSbshLIs007b4Hrt8cER0VjMSE0p85mcvl5qqv26aPAGSIOwokVHfgXaDa6XT
s604jJChedOk74qeyMLEln/odLeUam1Ta97k5E6Vj8YafBgU6+eQYlolgFJ/jwye
SsRXAymSfQqGjUXbdt+ZV+Q7sGJlYGXAmBHvGGZ4pzaCWiCcgybDrdjq109AaNpy
/mAopsydOlNBqT7BcxYnx7w/DSK9WZusAigF8i5dOCjfrL0gnBRXx9gjMEoCNonm
iqENjRmyHArZRPkdPbvC2s0DNAP1bqEmL33We0PzPwg44YCnf+Xem0DjUY7WYsHb
Oqe83MshHm98QvpeslBVw9Rmmexb8xfKa92U5BD3w6cPWFp5TUmSvHgF3L7VwsXN
LBiYWoW/cnfrcxG+CWTsSFImGbPpQeZctYBlGRSQr8cklWTf1vfomwEA/eBm6xXr
3y/4uqJr9oM/1sG4a+ywnAWFQ4wCJNfBKflGq+eRJr++VxK76Vlm4tv0OrpIPEOo
wYBx0qAxBBQ3Zi1GXUBlAS74c9b4uofqYmMV+OYBVsTe3YABigOnqomNmm4Aof1k
HAfqZH1ISm2e5olvikZAoX9e9whfUXGxeJPISL4wRDO3MyeGtlzm7hNKlixK+T8U
gCbDgd9AtnqXP/hXRrCqt3d4NfW5rvXyzmx2y6MSxahNnKjiwSpo7EEegwv7IkpL
91vCzR2W2+JKAQI30rqPkVAZl99lOD2NpwsnhAeuqRuI54ej8sOqXhJzRJBn3eH+
kLMDek1JMSkizP7F8/+6UICSmZmw59wq/jSt++KTxaFf5zx1m5sDg09SN5ILBxd+
wiUACMDTtqARmSUIWVDXQO4ZHAdF4I5xGz79Bl/uv5DCJ8loPvEGsZssJmWVaoZd
9palXPEHroJD2CLaeV/w8KECW1j+yvVfAfqP5UPvBC3pnQKhg2lftY41Vl9H3+70
KLRLZCS6fFQRuEPKl/Bdyg+WASThc5OzM/UT5rIrxVI8uIX1w7nTjz5dnCoG2pfW
S1O5BiYOG+bAQz5cZSXLsDDMS4RiBuPn1Rx74ENlYD81Jd2z3vW7SJ8vYMrtJrK9
ksBU+HR0X2KdkbnrVHyS2dhUysG4sJRhnQXUjaDUPZvVy8GFf7+jRsH8WBHGf1yz
HYjAE9HGb3rF3ZRYAoP/z7LXIxI9yBgARJoPFJqV2xxadCG5lKSrLiurgmU7jhor
PRjp/gZ+UVUPFfzpEdyVwvz7JHx6AvDo6wUA9e+ZGFE/xiIoUNwiW944KAoObY5D
fEAFdIBSLcvSgUju2XLj3veD+5kVmAdm0v5Wbv/ooSYTfo6smWatRcxd4cxwg1Ac
sSCvPeEZX3cdc9Jf5BMcPAU+3Mw5zL/pmSKK9KlaMSpZi3iLTksCPifSx+4K9py3
Itgy/Gw2Kx8lpnp4IzrNkAWPzVSvFO79FwhMWA4A+Eruf3pWPLW5AqHmu2L3dNHq
opW9RXsiN9aP0HIiOQHNfmZi5codkrHWxSBuSM9r9R074cYsWmMhAJzqKiy32nIn
YkPHKiGaNL2AbNAwVZ/72a4nT8xhNawvZS+30ZvPVNukuCILTTDTsJA4sIUdts0b
S94krbWsZbHoHAwCb2OkQQjOPnq2dDfMHUQBx8U3qeJF72H5snrvlVic04bBhHH0
q4Z3wTIeYfXBZR90hKRY5KlMNI/mv3nEHUnF8FGWdrV9QQNLenEFeV+0qUmbgOO5
MLtJimfpTCxkXD9vIbPb5u19dmUAwN1o/h6bRqUy/uAN1kCqbg7di74v8H+dPgLC
WDZeP45drP0beJT4feYw9LRycUu48KkIiM26e5FR6y7uMYmkQMizdCaqWixNLpjP
J/7ERd+07kTZwgUlAHxoXGA9Y6BTdJLI98k6eS49urqbX9QgiGjWS+zXfSYwoc12
VQNHXOZTHng/T5pcHCnOYanPy5MySaCzuDWwi+C36RejsmhUQ693nVcwUP2BHdcl
Nzis6UzLvduW8Ui/TaFvJhVgonfkT0dYIYrdH/kbzm4SJZjiBDI7ks1auOuH0npd
7Ixyct07tUSuelNjy3HJLQkulBp+NdtshFb7ioTVyySwcNAdfqtRRLx6tnsIwJMY
yfC4I57tRhtxCBAVVX+ieThvfVTMp8tfHfRG+WoxqM+rSdbymuonOHdji65Bk7G3
NpplHTqqVpObtDuSdZAiqmu8+qvdsEaspUsNKNEaypPRZ4GxNqAPGwhwzVyHMklp
vB8vq9uTwIygFFKOD+GcLeYF0jFUhHb8HAPltpWv5zYhSeIMKaOdIJ6aiZHdH58B
U86TBpBU1hPafW1otQnUVUowSj/xSIeMa8ZUKsIAJJFWraRXupo7Nud2dCf8AoHQ
eyjVqAIJYXzsc0Lupt3wCrLsdjcbyhfQGnk1AyEtH97FSNO4hXZ2sRU+vp/89dGi
qKGQot1QJaPXEw4sujH0ZGBL8JbjOc8paXHl3XSTm6sC0EoOLIOf/R8A7t6a9Gt6
bjNhGrCgqX78BWesSgukehMI19U4rT9ehdIzbQ8OqhUChoYDPcm+Lc/sIGlNlWKK
5hQqAaXRxSkNwPdzz8e8/IeEGR2ncrZEdkwP7DcO7kYVnyChaAwOANjaxQqGLpOC
1RZP2TV/pG//UfAIibtVovXgS/kc58hL6cvoPIrUhJaO7d+oTIjQihkAE/zVqoQ9
icamIy7ibwXtw4ogiFv06TTFGp7MTjksYDXpF+rtpIBpIEKrFK8/utQJ7mJldRt3
oUt7hs832Xuy0NzWXt2VEYw+FWCbfMi5N8B59NLts4t3FpB3ImNoYyH/wFXuUBHQ
43j5DF91BCwOVUM9vg7cS6vArzgnaQz8QaZDztV2I2ye4PQWA/GgvtLFFF0AGd0Y
HyPJLBzvMX1hRm+keHx1UhDLx3sIytfAwezqEX378A4Nuav5ujQfVyNEPCPk2HVi
QzokzTuvpkr1iA/7nDKkWqAuQXfAxch5K2lEsoSVHlnycFEjnkfYWDd/MGLPifIf
ep3nZ+aPWWb2u9xxzgtqyl6QzOEtZYH6b80c+gX/sjThs1Nbg8stbicoK5F1YZZt
J73MyPAPx8DeCTpRGzYuC94CVDWeFERd2m1SJNUDYMGuUAaOSp0RIt/RMmCaopvB
EUdc/k5X3xTxgnoarfFxxvuJt8O4tDGq0cHobRdPfvyCyfmq0hWcdL7CzMDZUFET
F8mGw9BEBOc6a2JCQhjAIBdVolvoiOaAbUCwZlbaQ/MHF6o55hG1Md2YogEIe2kj
b+x/Gvx70tdxUtedxWoPonUNr4+T82S3W6+HrfSpNlvAIH/T//Io963h+MirZclo
aXCtIV7NVWNADg4g+b3jje2vFph46Vj+5Bc+KhGq5Bw2WU8LdGfyFIu7FFyvPB7p
RDiUfa6ZF21G/faNRRERTEHO2iVv8GUYN50KqlTxeKWOTRCFKYHzZsIb/Rb81mXb
1ACbMhlW3zJpd8QiONuKonifIwuyc7OsFtEqDuuH7DnI6mq/7TReXRO8+Emk4IHq
ZDEk75UuP4HaAGJiuOCtTcEVYStqq04Wtwyc8gIzlhikpwdfbJJG1AqrPJCoEVxZ
xMxIXTJYagpMTPZ3RNBlCjiWNE6dPII5ZzvNw4UfM6e0AvW4SycgpOLob1IYDg3v
VaSNxNpgqVAX9aJq1fDBAgVtsRfyezs3hR7K4WPTOcJrRpAtZSTq5R2g1ql8Vyjq
uLCvcNxzZdd9vw1wUgpbUEdNHsfhsHwJJ8jK1fw8cIyDVor0FWU9ygOzlIoqsiaq
vYjLS4V/rqEHI3dqalZjA9jAfeYHhJfY/rg4Q0gZ89pPMTU7hMe9rSGnB8iEsQYP
GqrgYGWNxtfJuYJsf62NY7th9O/z7PgsztAD0tlJ5XQMJTI3gU6CiRxCATFGrZvn
7k3VowHHucBfc7wMNlBG9g9Spp8YnUJxJLsSEHzkAw9SVJqTv/WAtu2Lf1/Ii5qW
akfP+aOd8c1h+FWjjJsSqNsjDUegZhr3zehZjFSCLzD1H7S6DM0GM1/j1ze+bUEk
p+NItZOhI7mPra3xm9U+8vjiAePx+FnpoqzNX1fUPXUKJhvF04jX4JB9hCNHISZf
tfYpxBjUCateOBQNRzlChNisANzP4BQhx+JYKlrHQKnPY9CpG5+meyp305ExW3Iq
ImuqX40FiYaoZatlVDzy6EMSUt2ZRObn8FqDCZcJZY27rVPpY72+PYgQmsSUBwMc
j19i17ZVOskryH5JAkV81ty84/ALt6FVMnRERV1l8rKF7JJX2sX1d1xVxvEii6C8
37QlrBOoU917JFnm7kgASTXR3TLDaD3b/hlqyO8C4f2Md5+Huq9urTUnd3iqJ2qU
7KEH2xlZp+kpFDw17WTQ9ulzI81lkIJ7/TgMtwvZL/SQS+nFXMOquNsw4jSrAodU
YvPkO8c2zzwecxSxKLIDeWkPlAhb78VqDU70AcLZZ9lfE69ai7CKXWoQe8vzN+8S
veaF3bxknpF3l/PqNHPUEJeLTI6JBvp9hJkZ5x0QEuvoVUZ1D7ck7jH6R3Yo5R8Q
5Tyj7L0N2/nNg14R/eQHkL50Wy3gPsgQ6GlorgkRfFLVJ7SuaQ0quXIS38Ope2UA
1OXl5an86CMOE+6A/1rkaqwXAcdR6NxB3Y4Z98z6bNP4yumwGfms8ZRBdSyYs34X
ZU2bXRsQXAuiRcrcWrttxbkCZnrGmS4POdBEbn74IfxgKEF1Hn09B37r2fvRW/K0
NwPo88zXRtHQZrsscYvAd8eAflcVWfwnqjnoxci494tUDHPUNyiE36lYoYKYk1lk
+4oqhUWeOXUeIOyVrLblO351ZEI9z2CMgfCTnIlRqN6XwsSxETEEIBBCXz/373BF
qhnMePoej9Q9Wmh5FgWa97j0wMtCpzpUraFLhRZm7mTN8PZj9DULQ6591wPaoEUT
TWRGvMMAok4jcAy8sF4YuLXtxzlC2lm5AUFACZYKCXUcEqTOc/xEY2yn9mH2GXIr
ML3PAVZMhRrvANiX7SPSrteDuY/HtgYXvzgl2VlVCZi/Sh0p9kZyW/NKplDZRBs7
JGaZrSHRKCSQzhNMej8SWruFyr2Q4m8I813Ou4Q14/p1/4KjNG4sfpZ0V2Bsmdkd
yLvw8ydI7y8lSxWcqEIs6/W1LAr3VANp2t79FK8PMA8ivEyLQo/9W3wIT8xArdi1
AuUrW0GeRfLKJkdWWCDWbLTIci8Z7Mm3BYw9INFvKf/ZS7+vG9RJ5I5vsG6kX3n8
Z0aEM+rJaLJpviH2jB1DypMUSSPQwlxBtzAFCVOm8kPgCbElv+rUoREgNVOKOwpd
GyUW3JoCyRurHElCxvbKRaapONdHn3TqGUULuzl3Yi2vCONYz3sGD+zo5vMh9TzK
TDgNQSWFzGYYCKO4joIdPr8bfvixlWYtH3PXTQAqahV9q5ckNBHwvQE3vMvP5sdI
NiPJqbiFcVR5krDIhgN1cVO6qmP/IMocYG5VHFi03aU0swKr8vmFMWfZDnmOzTQT
CSsBOLaUppYP+zGOroGJomeA9YmtVhqXs0eG4k7dhs7HuMrQYtuTsoKhBf3fWemn
dRIUuvbJdRryy8c6rhMyL6XQj0q7bjsMZ97cf1uEwlPOKyeV8UlrqaGrg6+mkGma
lkLu7DkcTmsGRmC6pgrGrjFqpgRuboavbJmBa1vJaPB19OH9pWjt0AD84nfK8j2v
kuqiCBeB7gMLMvPDSBWdrvt8ViomvEMh8IkrkRA4iFoCUxQrtZZVrOEplwP3+ahc
Ib/RiB46jrfXJjJjgkXt5kXy692CxdEVGgOlkT0+tUZGjxtcYLWFis6aDsASCr4+
I43QDJSttVeR0ylCCJ65IBtruC7rR+j41yRuJdDdh9XfzvQRICBFw4EONEDenNVc
XwvqeBI2zjoHyeqYa+p1vnWWxgtatJCtYgqgADpnoD1ANt/CU82vDLlUF3jbVseZ
vYaX7CTe9L6eJOUMgq3HnyVdUuSa0fQ13RWOWpEhodnkZs6pBTD74yYe8sQfVQg2
EMpDfhiszwoHiHJEcs+54MTT+YXaGnityTLJivEFJXOs25jE2bUO3B+iYtGZ3zSE
jSL4wsy7HfIAAtBY4KZe20i/Z3N2AwerWcgDOSfhQv7xdIiL+yAtP7pYOkwULBz1
5zQtYY+HyVMNZ3qu7NWsE6+xhBTX/xBssluyu5WUVCzxL39ypjgUNlxMtzF3fc3q
xLTYwfHdPpDvEQsTPxfTFO8LIsEzSHaNZumaFB50yCKIH2CDRkeQ1u4tOM6qgXXK
e84V7C5yZy2FPrWrjLp1540vficT5bGegUXEesf69dnl8qYw7I0MeECiCq2zmTZq
BrYXCgUheRds5DGVr8zgtqGnTgAKuzHg7mRIC3LZAZhbxWG3PNx+KRJwJKlz81XR
q1JKRKH6F+gF/afPtF+FSWBqCpcGQ5jPIYRpO9bybJm4nigbYcHbekugjqtANdKA
SA9Xy+9qgBG8+/WFoZjOQoN5W2MgqxTlPRF4RP2PV9798goHfuHY+UtQk/FFTg8Z
d7COsx3IhzYL385UQDMAW4ri9iWhEVNKt3+vvQsk368IVs2oKVfpB3GPKa/ZHJF9
tTEqN3de/x1mBF4oZ8+hB3DNsWeXXIP9109ZQnRSgER0exJT2LEziPxyEseiSMCo
tBKtwmliX0Ju9Q1OIHM+5O5K6dC/v4qYkx1xwsR3K1uVi0Dopi9uqcHr5GsBZ2QN
/GEOwI70yH6N1N3FF7JNq9YCgUGOAesVVBTRMXoYc5nq0q2eBHplWZAH0n2yT5iM
yyRQrFwo1cvq/alsk/PmdqTszsoMQ2NY811L3qXFjLbqz7INlu7Y+eWjDODjDat6
M7eNMeLyrUiNp1OehN3EYlg52zdZo0om2gOyJ0wNLMSNs+Tk5smL7NWFE4FjyNQl
qPPAwKMFBN96kigD/J/DWixePvHbJm26B3aeU7CJTZghrlfrbISuq/QTOHnhl0hO
uxiFOUK6LhE0RrcLM+4Fy9RcL1I76I+p2HtyknkB3vQ9ol6kLyeFzXFXihd+sG8P
NwQnpaKOJJMOKs50A8cneK3tR389J5de0ddH3mk+DZ2OFrc/lnkbpvthy8vgZb9i
4zI5ywRRpRx7fPuPzlbh8N+lyCkElqY87skztwOaRXO4vUNJIQvNxF0qbzICmW9k
2lqGsxDsWHsdKomUqq/ne7MX8+v18L1Dk3i8xPwRG5Dp6RhnDEOxW5vyP1aWtSE2
JUEAw+so+coNQGKgO45uW3nFpNy5MjUt9Z/Jx7Aw4zdnzM3qdnDctY6BQZGGYgo5
LLYDZgRN1xB6yJpvVBuGGJ2yaZDR8m7Hglnv1K/VkN4ix0U+EMHGsSxQqwyELGl1
NlLFLT+TkYZKtfLU1zQFViIs+ERgAktdlip8w1VlffmDeka7X8OP/QayXa6DTB4z
RmPF7iSQgVn7q6XsopBgT5CxnS7s83WGxT1Fr7KeKx2LKpx2OVciPaI0qtENsGG+
Q2BjyNoU8/17MHpLOMEbwfOhmcKAIFGvOoPvsGIlIC0rlHesIJgNC5DoaeisD2ZB
jhybVJQlTtV2pTV/GAF9QnRkQt+4EJX7AnwKyHYLPATUZAPpl5Kx9odfUXgyZpKb
sethjArgPSm+Wnl1fuak8LYwRsarPAsjRJXDW1lQPTHKr/emgsOY+4xXCtv7c12l
MuST9wexA0BxFwJl/BqahtYPI3/cwvVj91jGoDQdIbosbh6ALjkIGGHzk7wBASex
9QTsUgvDD7QEdSU1b5nQM+96kPmP4hpP1xjTmvJeUn7ZZrXTdec9mdg5QVvU5mRa
8BdIeCfJm1AfoOW5xo6tSJRjt4lb64AaEIWI6dJC5TX0tYgRDrYBTy9NHXm72/kq
s6DykBvOZdm/dROqk8ntYTWzjT3JePjYYmnGU/gkokqJeaIqXyRQnibWwo3Q4TLM
sUcyhr5rFvbhChZsjMwJ0lZ0DYsBA0NswQ4UgcoJtDZ8Yl4mZ7XfbuzzrNBCaSb0
Di2VJE1n+SbGYsy/nnMTwMgARlFZiPyipT6CNmtMA87fAVtVjbEizjc1x6tfv76b
rq6Sln03bKAlOH6jZ48Cv3JthMYRcQUGS2VkahbKcmIlTIAVlOlp839e6aKDcgnT
5w3NRkjr4w3xiVcJp5RHrNSlILAPrh8ZbkL5Jm4PTf+v+SQh70Y0jH/fGsw9LCEu
2tx5wtLLv5mjHVR16B+kWHXF8q/WmqKf477H6dKNiN2WDcbCw0UyTMuSbnSLwRRc
L7QkWoaGervSQXVMDTdaol0mI7vvKYsPXxiBim08GcC1EGyb0pyz2MKWjheJHhAN
ou6Ew9x2sW2ZObiCzqSGfvGmlTc8OgWRMGG+Uho1t/GewLc+H3y9g3mrM5y5p6U3
sWzcqw0TCvhOwcATTKJGNaAlw+NZD0ICtCf21TJamfDtaac+GbDnmIfqATIjY6FJ
LN+VCKoSGyjw+/RhyLhThMqN163rZFpvaiXqhrxj+4TguNcYs382JogwSv3t4mqQ
TLVCZZ8JejZLcnBB4iSoiI+hpsXLHmR4iX9c6U8fuDc4vBgDkv5ypnrIW05AqrSc
TuALiCOhBiHIyBjRNN6AAcjjwgoj8O9RHIkf9MWoqIDOfubCsmsg2Eq7Myigst9x
IEu38lZqsdKsO1CZGtLybxFYQmTYqyilQ/ZYPXX9HpoKAI1GEsq9vTmaQR8p5ofG
cRjy4FR/hMlDDHzpBezVZxvRjGJtwWN3yx7ldOvuDbSEupL3exMSKph6AsgiabGH
1w0wuE3KQHGDgJJJvA+1QkwwNEhkgAxxDqHwly5stOKKNTWVMnLHk4VfwKDd3o56
Savy2l2qYL7lGivu1ZkHPIrAvEVyKjSpfLGJp0woa/N8YxqKvs/5AdbYBkERReWX
G1W8tDHHX3oKjVcSUuk2vy3qk+inBhm8LH1ONwMmsV8ikbdXqpJ/vjwfjomeKNRl
sQi/oYUTpxE/kwKFNO503oFfnwvBYYxw9U5hUFIzJu/5G8O6zCGEUgWAFdRICOW+
Azbmv8WAkb9+oqRl546Muui0MWJzeqog19ioFwm6xU2QT9hLkDlCqyHvis7WdqsE
iNIZlv35TyG6HHaOL6M+u4tu/hEoXFdkzFgF8aYtoa+ZTqHhfObkJ6WrcDDRdkwX
TRFs4I4i7ZITyGZfSgsoLMygXbvlPsxWJ+JzaNLX8ogMXxo8cCyavbyXWCnx8gVG
2b+kV6qOmPRdQPT2ZC8T3WvQori3eMFXeUCPxiafhcNXqzzspWR1H95EooiZ3tea
vm+nQhZg1wvI+7ZusxdDzIXgrt0Ojhmp+Fnf/UZiK+H25Of6k6Tb16iEAD97T94/
95R9iXjGRLtzBLxfjjS8eOPTlKoio6MsXxTl87dr7FSWfLqZynPFosTH3tPDqiun
xcsTBl4ihC+PT1PPuVLlNFMFL9ASU//jpBRrDpHKykHDv/KVf2avknpJ6n0jwvKH
10wxvJvl0iCOavmYMl0892l9oCEeBMEwRSZj4MuGCnXheITkUD6Ls8yLrwAod2Vx
WdTwnusSrrpcPuQqnDdeQKaEnWEfX44pw3Wnbnl7+NInTlCK6mUu/aesKuvn3GUI
pfjdg+5LaFygzVZiKFF/MN0YqM1nDrmW1UUu9M2m00y9+KPDuwcILhMosGyg1ThV
9twmbt8FPXiUPRZAcWRKjW9JSDbcbmlRRCYDJzq6/Keu83iJ/uB4WEll6Z1KP2dK
rQHndnmELNXyXtIgdJpnqFjIYB1wwxtGl4b9eIFHXorARpfT/8ipADOPmOc3eo6G
NR6wSS2T7KheQEQSFETHrsqQBM+2zxbtWQURtBQ3J7xqRujJst1o9DCQmtRaXlZI
ekQsh4SMweuaFMK1twNuisxP4a1AtikALkFafYsDoiJK9lvOfxjtATYXQ/8DRJJt
VI02OB4O/vEEbMtLFeDJ5r0V1sI93Qc8os2QAJ4Q12yhVBYi87EQyxxO37k+2+/U
3NVzugvQGOoY3E+A/z2wiaHz6FJ2j7W711rjzdDVUozwh3kwgAgR7MF75gYpSg7u
XGWgxZIYHJC6ESv7tYcMTeuVhqBL7iHB85lZ97/67rMgrMiY1ckjxCxaNPvE8Gwf
6DC4Gaxfww5UYABFz2tXULnWmSRupS1CXrklrUDwiQa2HrDa/EOOs6M0bBy91qbA
kjCQ9M7MlWsF0BuNKw55E2cdaLuowJdZSo8euRwpFvolMJoHmTzUKIWuk71x+Yiy
YLR3snyk/KB0oH07j8bTH/2cn5/fr3ZHmkX6juKW0Zq4ij+9BuJ3ILv3bh9GwNT/
iYL20IaMdWiJs8YdXWZC/tI4zhZvH6pHi4iFif6zYbAGwOpDmSbOUeHOwJQ4WluI
rZ+GTLTs2lrcxkME+svxTYfBOeVflD+tjBwb4seLuegVTWAocEc0MsRkuZjvdkit
DjDyfHQEzptheSBRWPfwRFxo24zx3st6lEdzMU/coepH4KNtHFnSCX6Sd6P9XUhJ
6uiMktwRTK013WFKPeu8E4tArB/xBXjM0OwwQEq9iuUIV0UXJ7ne+Yv78tDj7MxR
LCrYvxfcdLtcpqbQAtE4P/+9GtwP3x1ESBZDpvzqMJ/3nl8J3YCKQdVWgkdTq3EM
9LzRo0Nhq/H+K7SncW1o76yYJx2AwoGEM5t1+i+7FfOwiZR1YgG5apamcnA2p1Wi
yc6x97JqfZcJkCQ+MJZsfnoyfHSGr2U7O2JW0OArPOv45hPVAtYk4Sxgh1MlMSBp
Dklt5wNxoWSsAOBg22UHDJA0MfjgM4lVLLyp973G8s/qAvXTsb9NSzppc0ApfmcU
HCQrUmBjZAW6mX5PnhnyLY5IusAdntkvqGxGWr/IhoCbBhjvhR5Ee8btVqqPqMx/
4RgSwiqgvARTU7V7T7n+jBMFJqM5luHi2pm2kYezsQDEsQV8siT3BlovA4/m0mko
WuiqZ6fgktA+rSD/IVlMzBeB0XgkBzhfJoTmUWciLV9KkP7qhI791+bEj6Y6Yu/R
jXdCTIgtyujdY6XjPjFBqbEYuOEsON4ubmJc3ut4GQ1rIxKcfX181V3uOnyrZXLp
/1Oc36cx04BISCAffJtRNEIG6RN09SuHGmQHihqfCAaMRqh7emDUIeRFvM9R3uVJ
Kl+B+ix215v5BFxLc0M5gnJhg74BHcJRYCLEwfR9NQtPwW9hytxnmL6PuqLNU621
1EwwvSLYrgiZQnk7JnOTITveD31PMEMnTfofbaQzI5GXexCRxNVg9lJgdZLNqi5d
mY1N9tAEsZ9hTO2wFc/sA8jzydDgGj0mhi5b5HnOcbwOf00hhRamIWKqX2ToZsWS
czhtMDP46NBQcsrFCXi3+J48jl7vGuyjDaEIPpr21/jFFy7G6EoUVwF4o16/DPtD
LGJktkywIIdcheQ1q5vNsBxVJ7riqjNg9SDU39s+Kw5+P1rJT9PzRo7luDCBbVCR
8/rl+IqKA2wrKTaGqHBUNZsnsH5DLkJ2hfmtcU7AuZ/9a6HUkkl15kwR0AJcxX04
bVq1GmV/+hsAELZV9S6LqhdenIFr+hpR9hrN5OIz7+CF2Die+THqLF6WUXGYCQty
FP6fen8S2wNVffEA59LN4seyag3dXWrqSIaVZPngR+A9kytOT/J1ZH1g+9hs5M65
U/gzZ5BVgNyBR9+VgnAtGhBSCJxDreFDl4JTOqsspMg77cgHF/4nDdE+a3Y77tdv
LPXhqBDBg187bYqJIrN8q8MwA5nxjbP6kJY2q42pgMWxzpAxukuKRk7h6TvtyyOO
uTECjBZrd8JUTYap/ByY1q4vumtRIuGCdz38AAItO5LzwJyzXm8CKUCkMaeYnT5r
GthtYQSI7UnDaR0+unTrpM97dVbeIdmo9Qlw6dOwNXTBUhsB+NLNSKRavVoW8A3f
/0XwZHOrDumD2zRFX3VJHcVBXep4W321E0fxob3E7+CAV0Uu9oBenI9UJfqfnlFA
OwqwgyT3zgN+yoBtoHkqHNd5IR5C7eVg8bxM4ezRWpgYU5kAFADqF9jFlfy0dHs6
REGTLlJ4MRTHxbxmT+vnB5jCHWd5Y3NpuOl0AfE+23rHxZ8zCvACOqGkI+W6VmKF
7qhISGEgICijrarLTfdjrfCrsLKMlpxbVjlYtxpzQR9DlOLgntzzuufyrbV5B5ye
E7TqOUvqvyuLt5JfqiOeJti2F/fd3SL+sL8B05By+UVE6IPQlES639zYhU21JtBA
h0SzxBCf23y6gm18DEGE10WbKMPwjPLGE/MLy7Lk1SQma0WJ/MOwHVDVe7dK7uKv
8ZlkQ9NqNWMHHhXJU+AtAl5JIEXnuLikaMRPoSkIsIyF5h1QEOH3GjY7qm8VkZu0
/zB5/xqqBXeXegrBwFoLvBEUjdMnIuJPbYxrgERtOzc/QQnlPU0MEUoPsWu6v/ya
6i2GWvEHKMdLYnz8nPyMflU5tURkxxlnmY894KyXDwm4KcEyf81/8c3Xfex2f53Z
F47AoB+D+IkY+pqVbSsUZZdXJjoNKcSdY5x/IFnBwJplO40fvs+A4v9Z6upvlaZv
nRgSuKtSOzXsiER8Cjve53Kxct4/jLjJfIY7RsOXGD7tP6co4ZEpFOtw9s/Wj0B+
FlA3tblj5rVEJw46m1IIqdzecHMfBaOSig7coIutTAZIgdJ0z+DqmiL61Oz2LUlM
OjY7BWVg0FPdBpMLzzpUwTGu+9wDCHqNTPFEGqYN+9XQkpmYd6/gHwIc6ZafCjly
IbuaD0I5ZUV26MIyrKUwNVGZT9ZH8x9xvPCpvngQPfTGSapeKQ0/wvrpwFD1WPr9
UmurPmupa7ViYWOTMaivwhVnIO+cYhuzvUsCUrpaiSc7nO+wsysk3XrBg0q/nrFv
Mv2U+JlQRHXO+/zMbSiUu9ZGnUwFuVB/RNzkQHmU+kSzlXrHwoU76ZivOB8pfugS
ZpCczHoS2v+5/PBxeWlvAf2Mz1u2N2UcJzgizrUKLG09342qFLrojN/zGxQ4oUK7
r0o3FuFIngvSWJh53c7YBwzCyY1FQuotjfGWeBtTxCJ5+WVyoCZPXRqWuAaXsUzL
qbHGuoyJ3bUw1sJy79jtCLFppLfQOedPn5EsIt0rlhPNP1xG+UzeDZWzAqOnKytG
LxU5mvlG1D4T3K6P7+k+sda+2vjzqJwT2bqgWMN+I8eaBPZeLc3apDwYPzw82BPF
xr7dGWaXkwHFKdKRwQNnVjJwfmLdFJ4fGt4Ypjik71UpxqWQOx9DFHyb9yzz9k4w
DJjeZTYpiEUXKNS3JQLFoY71DtKoLAjZf/cJgy0TbxrUCNv/btAPhBEglt9jdtqZ
X1IMyPTRe/Rrqx3TYt6MdfpBvaqYzPHw7vSK3amL/5OpJfJnf8EcrNAfWnMYClVf
Rvbynm23D124jjvh1liEbZL6La2ShC3at9ifk3DeXGlcFsJD9693CFDXPZIpau0S
uRFP0UZ8ToH3z+/gLMEQUjjlXxfT9NqA2XRlIbt3f8MsA6HKQyijGqQANyXrHTSV
yebg8g4vmChR/5jMEUejIvuaxR/t5I8tr+hkUwM7NPApdYyDGyqmuDpJ/cnz/X1A
gdSeSDAACtRJthxMHBctIVfTAAq1SrNx8Z3YVF1nDWJthPhO90Vv9bog4SLJnjeV
/f9nqxkhduQ372r3/9S9HuU8Pg9zOw0GAkSnNciC22n+2sYdhdxvubNmddbk9Dbj
Jf8OikllMteBvCpAwkN6JGa5tx55RAwR5xEonWihQj68diQe21Hk6Us9gq2n5AoV
JPylD78jpuD6glgCHZgxIemCFLG8e1qD62pxMqkjglkdvmvC9C+vpqOW5NFK7vDS
7B5cmzP3KpaqaPCwKGeRSOztHyWrs1rCDXpeK7CgjxWIgnIj2pdUZdqMLCzzePKl
Her32/aPbPYyyO+1xfB3ioYjbBI9mo7U04uZMFjKsJfUmrroYO6HlfyqsHTaY5PN
VMyExqXarpF6xk+auUV9kYYr8zibk7468GBJtVBsj3J1iVHqm+EXTU95TmyBHFYn
HzWxH0n6+CMB0xQzDNzjYlK1Vhw/BbN4cXFLNXg57XZbmXPU4zROANMJHAwbwSnS
ZRcS34GF/0+XNoUEuEKTDOFOBIIjhcijRekZ7J6VNPozI3q2nAk82HlUa2TzPRLZ
R6h9XuKCXawl7LIVPTjUvjsQSQXtief6J1EvXNCcKGmhsptbrREFRP+jlK+YV5IF
t9LogqSz9DE9/5tORLkjbf1AfSJt4U1BXWUaTM33X8/IQNIJdFQ622yFg+tvK2qE
ntr0REblRfTttQ9fOl/YQ3YAwAx922iba5e3nodRT0lNH0LnkK0X8PzR/s4fzeNU
y78cqKoojCHjsujnQhd2HSY9gM+GVKVJubLegyDUKZc9PuHonTSpD+XdQbKsOX2G
mV6hs6oh1qL5Lk1YcVSjSb5XxO4U8FhYYa4EouWKloXW7J/EkDsbxftlDYBFjnxd
YjQtqQfnDJyAlsYbVLonS95ImVY9RudKfHFsL/vVyRJcgVKcnOQLAb28kC4CdEFH
c/0uoZgATaqrJN/6kZSGFNv+0RcANtfVrUdEvfBgYOZ8fqihjmVP8efs6tiznP0F
tAZAc0Hb3sTekUnR9d+YMIUIvSXgXUtednO0ntmTD7oWhpygiIC7J7INCWZekVEW
igxh9AkR7D9Da/aXCKcxGv21GD3Ks2HUbGaMDtdfjjhbbN787QaSxkQ5RGAjuyEN
JRv0ruRxyn1iRTcWzTnKyaqKY30DQX0qWMojcFDqHaqm7tN22Ilq/psd7Hk5V/sS
fLAmkrfWCF/ax+mqtHfGnfdYL2T5Iyca6FfmOILLtEpo+Hw0Yn0csitNcGQR8drl
kegcZetK8PwenrmXEpFvfXkmR5CYn7rBCtjRqd/RLoV2VUUrdk4QlgtvPtt/SBIr
YuDY9eBkN+Qnr++xbeZn+Vj+NmOm2Q/es55qyfyWg0AdxY8J0Yw6iS22d+hwq8Pa
0iL9ystBbdwSxuXdh1nTYos+avjwoPluaAVswgDgdEABrrkYJLjVeI7vWy+IyCqU
DeLlqc+Z5bu6anE3/yEJ4ys5DhQp3+ZP4TMmdof+esdGwAaj/zoipFHt6jdzJ9VZ
wyfZZfdkJQ5X+DCVb5V0bh6HcbIoQY19axoRsjUT2qI8xk126KROYvr8tU9ZlsEe
j+cnA9ndTYdQazSGoR+apd+dahd/C8ZVSY9m7gcXE1YdYcTOlChPODvmWe6GgYr5
NFQuV6nF4Laxbzscxaj+8Ef4pVO6nD6S0OLoY5Dm0wanM6YRzq6y7p6fVa9Tk2vt
QnLZkt6ANhdK+2RJNWGEFSDZQHBZCSBra+kZfsP2FD/fFQIo47+1X8NcAhkMBGT5
MJxpjvy8yhumEy6kRKbE0JkA7uhm0CgvYUICyrUoDc0g9VDCST3tO0HPwT6yvHgg
zxEPs4LIPmDWFLH/4qkZTR8xh7Wz/kD+ZRktBjXtiGqDBLxZiE2LeIiUJjK4saGm
qq6KlaIyP6dfLDnHqX51L463CmmTNWI9PDZ31wdguuSqQukHyikkT3KMToIIlkH9
+Fq55flwOhPoVwS6Mh9OenKL0UNHqTvgwSN0JsgIwEJkoeEEehZOepCx65si1zm+
wbf140yRA2x+lfi4sYWRZr0pwdj3l1jnlGhs+IOpIpEA7sZ63VGdQ+jsdUrvXHoj
ftVTBFRDLwosSBYu0YbGcLsDe0JG4xJzyl26/JsG6YuyXYTKe6wv8oSG+I7FzftI
5A9KFLktKTA3OCO19p0FRoG4f5BALARMopGYuFDicqcePN+/G/uEZvPHpuAh5MU4
zkix6xOOmgujabzd1XTLUOaXLlHkrDX/kwtKk6Al+EVLbRUBrhVU835OeuLo9Bcg
c80qfzhLBoE+CIuUt+Uc22z1JrjIKSuDG821T3LVSVyFQ4aHdrC6VfTwhgPnYlbM
vfw/LVvFFgsYUu21TQvbZN85o62YJayU3ek4hyieKXA=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kShqfVjiXbmzl3wFp2hDJaA24VEG0g6LK+wqWPsgVC4H/QAFDZ00AQxe2uCrQZi2
c3HJfGghMUMLCOaxGtQ3K37JiwPfLliJUlTPOA/Xob5UGbo2vNuZTo8CLYbPvVfa
SWL3MDVK//dlZGw2F2/dRDhoRyfkLuwKdZexT86t0V+eQIoZbYPrRWp+chZ1CHg4
eibUprKo1xpeGBNn9kHXN4V4kYOrvIZ4Iz0mjhYUD6o/YWr7+7J7uAdPsXqJrb0l
oFYHb+tIxcXWNAmsaQCqtrTL5PD2iqNSTFlMzf7U0clL0atgX9ZejnugUNRS1Y4d
dlQmlheBBLMT0WCQgo2LAELd31mTLoDHPD0kAR2epuGo/yYVtpww8fMBpfOtcmDJ
Wu/bdcpUNODvKYLXLA9T2kqeSY7WR6HyMxjiPuhfFxzeR9eDcN4uufkUBW5ffDDC
MFjRo3NqDHoofPxHmKIf6TzqBJ0tU28eCXpIOW5Sjfe2EksS8fK1UuA+0VgwYH20
ZMtC75xR4prAXTkiz5/RBaz4bKMUVXiZ2GlQp543v8K8Pg6qR9U8HbbGe+yObcFd
7rE6PF0+Nqzv6AcIQ4zH1MtMff70wpztwpf03aJPn0Fx9GrUzO87wU5z+U9dHeG8
pesWDpjmk7963OEVnk3jj7EnofhVRbjelWZkydldMMl5q4596D6Rm/wdoJAMitcS
+omAtTKFviXCIhJ8AVY9F4/xMDEmNIyFqYTy/eDEW1ydCaFv8o4zRpOlJ9eHf9OR
+szDGxjXLsAlyQYIK5taAWUSkl94oT5h+WHC9jDRMHFQGmnDUgScYa/cNaE/MNDW
DbPtCq3rChYaLA+YWI3DBoI4TtWqWr0aadB3Rjk4Ns+btJAZ57u6fZ8YE9Orb/rF
NHoC2o8cdtEM7Clj5gOAIF2ufpPSh4ABkoORY5hf4lDsuNYw8M9gNaLBq35smPi0
OI+JwhO8EfAwGjrT8KAFgw2etIVqE89s47aPk/Ld0mEI2CSdP9CpqXrAxXnZQp3m
LYh7JHV+kwChUC/4ab6DkqHaPNpmCSlx7H9XimJhu6uGYLX/JtBvyz7VqGB07NY9
ug+w/m9cC0hO8kjnJbgwU3VUl2Zvkqq5P9ZFjp9ecZYI9S8/Vad1clhEGrkfNkB9
F9h1mpEuiiLHYRVYLURQmCdjFUiMPh9ZD/kdVyZ8i3ume/4Ce+CIYWqhTEvCbhi/
7C/awfuqki7SHPU29CoVzwnvQ5QGiyc2IF/d2J/b8h9Kfiy99lvcxs9b0cHC/pVi
tlXZhxse+vopf19CTVA6lqA5495aOcJ8FzGwbCZw0k29WP8pqdOgd0+hyXY41TNW
LidZpUUj4CarVXkhqC4+8mg6TmxSZQtuViFY5yNzEtTX6767NdXQu+H+sZGKrOph
iyfS5s3Se+VWP3DRuilTnWH/EC1vlqHIZ1HgEZB7HVI3Up5eReX7vuNlGZ08rNQ+
405BIdgFXnVnDSqDN+7BlmOOAggvAwqAg/2T1qvRMHkabiW+BaViq97lsRXy+UNN
pstCgMsvuOdbR3+Hyhmgf366r8ig6qULh8nyVnUcTJOGudRwoBmdbiuObPrHgiGS
5h0IKN6mVC5bFCrnPsf+CgyR0FnoaZmJcAvfBqnUzWZ+YcQ0BRfgKln+Wrxmhltt
ySclYMRDyTI92FlIKwzvqe9oR11+VYQ6ajYC53AMBQQJXQJIo0VoPgNGdEm3Pnbo
A3FhvbLgip4WFnn5bnwpEMvF3eZ+vsXgCUucyIuTRhPf7omrkHKSXeUdvihJh4qc
MwEl914Ilxl49vLijc6YUsc+jsCu/KirSzhq9oOilFXhGVvUuTRXPAw5kDp5/J1u
LWK2EsdLy0nmLsSGAdLQsM8fd3PRxdfK7cXiF7/Epyw6BSu0qW7V/uoYYFyh8Yxk
3BoFnKMP95G1XxRjvaqGe10wpDnQga8wafP/nvf+zbLXvl8K/MWc7dZBGKwc9cU/
HI+s+hpXzHx005GrLygKLi9xK97MfIVn8XQyuhRrd4Z93oLIj9Zf4olCy8N3VWR+
I7g7yXqJM7EeciNrtveNsWoevhRktQyqCWuGIrhwt5isJdhGx7iwNg7T0GVM8TxX
Sq7qZPJSvH6H/xXZRZnLLLyiwWcgyKEqGXq6UpH8s59ZrMc5jSft1tWzUu1Tm03E
gV6K6EVcmnuGgRQM1Kl1rb/wvWhmAOSebJIJZ92rBOzrnRd/NS3uikUlgzPGdzgI
pD06zMpU416ZGA6z2bEUB3pk46Hz5SVzxJvjLkGp8L2CNpo/eToAoFzDvYwTa8RH
bOZKHtRNek2jGeAWaBQUTBWkNIOHZccAm1tE0ms60O9W2Ilb5QdOhs/Z8lFiHjUU
gz9oFCf/CeICXoa6fVfNTioU8SuDcKAfLcoTBfzshxNE5fBQt41VH9S3j9uoZd+k
SqjUsoMzfV34+wNQQUX1xW7BWcQgCvg8s6cije4QPmKgdV8d7sAY9rhVo/vzWjZ9
eiJMmxI6SK27kL46jlL1YElq+nS9B44X3vRAxntbZsDjtOOn9kGB+FBL0nS2OMdW
n4jEngre/MU5zmzOciin1xxjBuJh34naE9GMwDhwDru4/lYxeVrTY7udvuv9Uu3a
lJheb93AW5W1qb0YEKBjmZE6AmbdSQtIYhkHgxQJjs/vLapewIcFA9SIvnZdwdXy
bEfTRsVEgYJBr98nJcUIeqe4e6VFtYRsMeuM8XzU76a206xIplmDVZnNCiLB/xy4
7gB+3cgE8bhtCZa1On+oNsySWbYXpVKSmI5AcBP7tk68AczG8wNxPSuNZrtdiBdR
UMk888JG5pcuuv1fULkyq0FVhPbIxsUfXdMiMU3o9sWnlNGZEDBYs7vhGdSVGXX4
vGnVAbWOPjdBAYmKdjG2bE1kcbe2QclrwYlvDGppvdIjDGdminFH9Keq9Dq0+AdV
wADFuGR7tNLYE6Oec6mH1wnutfp2CaCFdtx8bd/KCRrjc1W6WMOKE6tpcD53zrS+
k19Zd3OoEiafiWNwEpjmZGuwI5f6unGYwqrn4pEvNhYz5q00ujt914sBs7TZwRod
4/2Z5qeqRWr+a/hrwF/tE0R1UBvpLveHu4oAPnrVJpAjsC1kpLxtxAnadTme5nzH
h72X+bsRmrILRs/L7ncmBT8Ees7hH9kEUGjNtTN6bblCWwGyyugrThxthIu4ShVJ
Qtl2IXX429GnYxtC5uyNGZH7gVY5kqWf5SztP1EAlvlJgcDsTuurnFu5kDTAqXDr
CqYnZ2FmuS06nmgHDHzIZg2V1oX7lGcLx9X7Xxiaa20PMLyNm3TYNlx8TWfcE3up
CDH3zj/EGhrREzvQ532VSTbdq5tdxAFw6FJwIo6tb39ShCVEMqiTekAZ9/4nGjsa
4413L1Ew4q2YtRO8VxVNZNpXKIMeNjGRoSUDoAL+3vuNhHzkfNCod2HKZhdva5D+
elO+UlsZUXJ5L+GYgzQ7+KM2HRy3g0O1A8dFfwSXBUCvMfzjeBkK1hMrevx6M/zw
oqu1dLwVPZS18WCVNvFsgFJN9PhxLNjXfj6fz/YCkWD9+FcW1tWNXJUjAXWFkPft
zkVa3reEY8qdyUK9eL8WrkqUVdy0Y/vvgkqdAgLc+MzBGQRglG2ExsuNvQpU3Xoz
GGgkpR5h8+smEMXRE3A5cx6OecFpVzfc6aPoaCoLV3RfN1SfuT9Ydi9e/Nz2Xsc3
CFi6GNABDxBTCz88a0O9S+JoitePv79GoaOFb3kjxETDTEiucZ24KT6lpJKRHxJg
lPAZ8o4MrtPWBoFYNNwmsqx00nRzD0R6i9W6lS/PhwYlQJmqw/fdTnRbIG7vhoYq
u/8W1sc1I1NU5j8zf6WWBvMkaVL2hK/EWmVZ74Ix4//NzFqoS0lAeg19cwGc7vfW
276+p54V0e4TBGhhD36vcbZreHdvVHZN2I3TM9P2q5LqGIn3eLBCGAMW2dqS5NJx
n4PFXE9BlgnrMTwAL4yAK5bc0B61EqtKD756PacTc4zPT6+A8GBW1FHSR4I2MfsV
C7dTomoJ6yyGj4wLN/MnOUQcuGtKYiPUfyeDCvrMq/t7qjK+rS0UWsEckOymT9rr
aSQBs4oeZvN3/0LPAFYMVV3rvA839BOuJrit+TjRNO0d72gG9A47SowmcRMvfbAh
yZJXNKXloDp0UjEHos+pTKZeWMOEXlbFBu2t0wqKSiJQAB7vkQjOUXfE1M49+yxE
imkySR7PMBCLcyGXe4XVFIFn+JD7+qmEE236tT5CUijFnDvnhSV0l356fc+G+ijy
IawniuT6KFu+Q4rRabzHIUL6r9WJZJCOcJSQ1lap6grI2lpGlT4cgumcXzgMACkc
QalpCasdruzm8z1ifLw2z8WAc71NoWy2ccREYdGTUHUA7PKNHgVcnYfEMLxlyT8N
iFP/2y6bAz/pnNEjZjxrEK8YPL6wTP/m6gMCrJhOlo3txwWAqbZT4cSRdvipXNKC
xSSJTY+vp43/h/+iWt3D1KVrk6s9fB/VmPGvqc3RC2NDdKjbA8du1Zi1mjNPfsur
v1/oAUNF5tf4xRGTGvSh2HMTzFJAqbtYnlb9s/U3hSOIiwqwzXZM5PkHXcxv31w2
h2+LqDytEGT39/MASPcrBz9rGkyd3Ti34tEtkEbe1AQci+qJLQjuVOXe40W7AvBe
I/LBzNcUIX4os8dBITjjI6J3p/2TlUb79aDaj5m9u+FW84bxmSgjQ9ukgAtnb/bU
xJ3E3Pe0hLWPLXnbLbGwr59OOwaJRfMbmAYYXETojYqrP44lYW/HEUJPOvFIlYJD
E418BmKtvMfMI38E7kO+v4aDXgOPLkRWMp9l6hkUxuYs3j30kT+8SRPIQDG1KlX2
GkcGtzEGhMOLLnoFF2FOGcB7fuumIfr/vnmiyj1yjWPNFzc5iy0lo+pn2GYW0dQq
syxrh1yT/xfgCK4hZSG2mC/hivS//OdtYgBxkSurtgCzw153N+nzYqw56wtP4dup
2gc96ZRgQjpHtzH3GWjicEHSLeRNx0QZ8kiZfIu2qsvJ9cDM4X9KUUZkPtBTSHs4
AMhrPgwPt35tMi8AQgCXbhKt1tbGiAsOESntYAYjU7BAsOLHp77XP7liy26I9b28
wNixoOxGLFruNlX+cMkSOE7lijUPKJ25lsNKWuXZ4+GpFBlwm2Xl41Cz4kLQdhD0
Cl36Mb1hF7SqzKssSv1YRNeA/6n+Zd872pgbydS6MuIEmwzgYADST0EdLXj7eJ7c
nwkOqZUcdjb/mlCsL98y1sBqP/V6VDZG7JirAdHzzhXiPdWqNuYKIduQexcX1uq2
oKynVZW2Iflx3eYSXHtnsMWtf5BVPrbOeXgRXoLqFb5lSWYBgK49B3nWjNDbv5Rz
e4XquX0f73Pl/YRtFB9VG6DBNrOxhSQXHscgIc6OGgEYkWj18yJ2foK3Ugdfm196
B1WdVkXWEoaFyrs7o0DNsVa9nU01v6qepTnFhtW9YEENIjPuL72T1vx4yCRQrGTd
05UxK/J4ygMnCY8hegDqY1ngEchvqu49ANKElbhFN995z/l4Sd/eHSfPrxY9eK1B
VE8zmRq3mLsIy5MGiroLuElUobdOSzZE6yCv8CIROpqdaY0mDu4J787pGnWG/res
5sTrXiRgrjms6HBJPVJ35AFCaGJ5WNLNGR2t9cEIK76Hc6rNaaRCKw57aSa8aJ1Q
vh8GY4pAPF3wdbkQr4gmdqadw2LuLtkcnL9zPZd9N8RsgQIXm/prBI/1PSN8okgz
D3TFSoT25bJO8RA4k/bfTols31ciPvFCZM/c5NADyOb2dYGwP9hizi8aQMOGAvNY
LUMmRLkudDrT38ZZ9kViGjq8aAW76hi/XATHa+KLRMVpx8RaFajxrKAcwBZzvp+G
RqWXFvR20I0ATbGLnnM1s8mXabToCRiRQK8ICpSKYeQD2GGa2SIIGrW8fJYLk1RX
LdohHwtBKIeENVa8UE+0bQsUSC6ps43dG4u3GueKfU9Tr/pCNDh2BptdVpAnh3AJ
KFLHB8jtivjEX9Wlr2G6huCWjAr8I+aavdAPdRJtJGzX8rtWwqAB82kYUFJBc5zz
qyhV62neCWMXLnCBprm3j/Za4/85xCfEgy8Tk2BNujdy8Bbd3JdeuSSA53BvIAnH
RDxhSp6AS4+4/yfsdU3DWsZCfQwsOxJien0Wujfvc8QRAgh2Oslwi+CVfSwVYTOY
dUwdkclbGLEDUldJIfVW2Wx2PYOitWiXiGc2Z/zKYw9W+snG/AKp3LZHJ4PooHd7
2t68IcdRjBwewDf3gKnFIS/uzaSk2HK1H/Zi+GU2Yn7cE6zgsICvWv6VZyjXtcJU
1nQpTtIpyS6Qd75jVx386Jal1ar+j1LHSSu/x67l5P6zOdJIGJ7CqKiGdBSAzUfx
4rfZpNBETnIMmaESnX7fqyBABY7LoUewhZYvYVnr1AK1qQS+lBGm9cvyGxUJSGjO
+LkOoYNf3962sZFIZ4PO2Zz9xk9M+OD5NFXnXkWhOyaWUXXHNgcVl77/vMXgvOXh
jE0YvD2OLHLhEu+3/7D0Fv37iQWotK/6bxruoEgYStTkYZVX1sxP1a9cxvhkshTa
s6X91ZxIg5M7tihFbcT3c1KmI3NTC7RkWUgSrns7RW4obJLgtRPCzeZLldRkflZP
ea6i2+Kiyw/EsE7E95MIYylSrDJ0DRN3dC3T5Yyb1D+e0n5AT0Ail89CsDkyJaig
lFNf6CevJsUM7pprh9U/Wjd51eyi9W2bDt3G92ap8FjLDxzhjxPCflZc3kv7Otzi
CVOElppg6CuoMzXOMcgcY2DfkCm0RrNR0a1ntkNzOk8sUkVzFQpM+hIaG+0RXyVT
JZ/sv6kImO5IiErVSY9CbDhd+QSLZh1/fOLzG4JSO5/leIhB0vmfiEqTkRycvRD3
gZt5zDrPm5N3i++B4jxZskSG9HWYjNoWOsqWDSehAN8ABwJvtQf1039LtDv4BeGj
38BPGRidIR+oDmxgL740U5Z61i+lryFHuF1QNvC43KALfubBG86F/C6d1vc4NASn
AWRMxaMsMrYvrRF1tO+fuJTCT6AGHGbKog6rRx4ZOIk6tOY1aj+ZXMno1L+JVXBC
VmsvGXCZhJ8Qpa4vBhMlqF8sKf9cxN8eNPvbFwjpfoCUqHe2718zGMvH+14oYwIR
Kgwjmdowq72TfJMIm2ifUFN8wMC7GbFfUeoZZIOu1//ryDMGd3J9b0L0DQL+r19r
vfiJOzCCPFssP8gWhQHXwv7Kw5ED5Raf1NWNfte4xo5m+k03q/IHERI25nJZ7zXp
d/6zETXLGG3ckHWCG2O/mLfwLkLIOLY8a4hqJnOAVragSjh9hV1aTFS9cHSJ03QJ
2pzHJwqs1glmfwSHe2WziXIq+GzwtcdNV+H5y0rGBHaTTIsaIjxQMA1N2kFfV93T
P8tPqaeItfd9ETefC5B/NsEiE/OnTiXsFUg1jC3J78BDMf2DksK35Okju4RF4kIJ
zy+UzgxXRF/TafLKG8sD/l7XzCFSSO7yDVsDkcyjfKfXaiWVjdmiDCJiYetd+bm3
8YapD9KWtpDyGWmUrgT6dA1wsPj+rup7VC5qUrJxQOJRXpfC8+Mol2SvaaOzvXsP
e9Blf6ajVfl8D2N9HpfC5E+tFS/Oz1CwjKtNoeEsCT45Plnxqe6/1gHByF8XrQXE
qLyL0j+N7EPuzAPu7lQKnbYonE8rqVrivwfg/mr7ci6llnyk3XxT2mxzqoV0nTUX
W4DAfzA22UoDRTT4+jA0BigfCL2rp8qyfDmvsgPnyXOgKg2NQTOB/5vQ20qYxlBx
r7p52vvbIN48LLnZYYBWjjYI5az6qJMULwYtLCPHLZGFArhpgej29tGpB4r1dbi8
WoAioAO+BwIA9nlW9acM7AIudvLhoy8mN/QYIHfuRxJPLEHyNtF1s+mNvudpk0yB
W0PjbrvJJ6DSjWO//zXr4xveNPM2v/BAN3V75CeG8qwgEy9U4IYX5RpqnmhrEaHQ
QgZk1mAmAx8DsoErU7UEiCHCiMBM0kOmViLyFVe7EJ7jye8xl9QMGNJ2IAGJCIoj
0cxga9cJDq57mrDc5k8D5V3pYBxZ5X0QjdH2VXGXXHuJ1AigfPzDGJoHUgWBpbVO
BuoG9LdWDdbFbhZu7xkJfoPQ27xLZC/eRgSNj1JJ9mghXYJVKvcFjeWodmHWW4QB
sGaV/fqOad+WEmmMHpmY4pTJ6kRibMLGTuT29KOdlqY=
`protect END_PROTECTED

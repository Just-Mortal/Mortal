`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDSGaaHZv5hNs2tE1xFwxXrwbPyx6qtyk7H5jgHykbSY9lDIjhC7johOahS9bUPx
l89TWnPfym756GqfU1RAtHZEMOLiudW4vyHvAKClrTzvwiDghSm86RFTBsdaCHi9
Cubwluoqq/dL18Yfm3UGKlN8zCSwnjkAfOAaBquOXWNl5XP79SEZ1mTjdeprgR9B
e9FYBZi4vqkIfN27kpIcdkZugsvVuUsm5z4W2sT6OSSmQTfxAb5mnH3SPj+ss44a
MazzQrMj0SdfVMQZahIuE/ixVDDLRFcRSJpmksxf5qauiAAhrjccXA46EbthzPG8
MCjI57QcIZBEjZObQ/xklbzEgXa+fgipIms9fs1YY8SweeZ9eD+6dr+reBQNAgQy
JwL+C0y/gkm2J6Jju9qTOX3Fn6u7BEizggPCOrXMLxNPa0bmo5Rj1/1g7tpGbx2m
CteHsL/G1IcGmIfps0J7Mn02bytLbAO3YDsj1u4l3KoAzS1pihgvuUdiNTqk7i93
O+ZAftFLNc4Hb/iaJzYXN8SOmIRGGa3KMBjfzjXqpJ5/YM48PBfD63ppYsargUE3
kyQkTGRx3ZnsRUHQVMOWb7Uvh+N5m9af0GogbjSeuo9M7v4BvrkI5brflcjfBL7X
6oWCR981+D70kRjqedlNANgI43A+cN8B+bkubOShdqojkAywNpdnVUPiBGooQrlY
cKVf/gm870w89h2RzMgfBWTK5zndQ5KFYr5aItTiy4EXlMHYgKN6EbTvHev2H7jE
xtP1042KFq26Ijd5rv12O6FMprKJN9aGFNtBOYzB3nFdDETBaQ6dhPZ61ep1KHnE
xHeRTeJfFGQRGVE3CTpB2rXUcu2QOm4enMVHzoStw+j6sklu4yycZIVEEtAi7EkK
i77KfA6wQfe4FNnijFPHFadjEX+iGcaX7POe0QWH+xA/WuipoiTKk/P1ZoJxzgje
yB0VnILv9HFjhoDPAOlcjUUq8Kj6KpphZcEG21O7k41237pgV6MZeCQ09KPezuZJ
E6LaFBdKO2OFl+HP2f7zu6b7wfB/k2asi5+BN73DnMDbvJJ2EwCzsTFYsGpNtLrQ
WL53UYgsfKyMc0EZQ5E4tadKbWqrsujgtnBFNO7ULgs3Ca1tBmLQBtqpPiBrhGx8
gj1J4KD2ddLZ+LDON8sBnUKvQHcanwp5wAStsxE/SuEZcWaX3D8MheeYOLv3cwcC
j+nq/EV5BE+Zu1YQe1ySOZX7L26UyCUKb0AyvTFasqbeyW4Idw2FA/nGcIgrp5pF
kuAacowJeCq8d0F9DKSizjH6qLBtT71R+ulTiRH+JbTykT1PSjO7+QOgayiwihfg
SGPQTM9oIzh/SqA1uAxM940tveyzCyPz/MaUx4EidKRSGSqPx9/+IwCrEUaLfico
k+AeeV7l3VwsymPitJPpCMrLRzunG7OKqiI5GnP4Ck9zm5sQ6elIXlqf8/6Ny0uM
htcQtORHo6pUFlXv9gzCFWlRLIWnmXl1EbeHdRxgzPownSr5MzgjE1tdmvNilezm
vyF9NYv1a449mgMsys1o4Ule5laIFTGmO9lNQ3lbSpmNRRRFqIpIJUFfnj2it0jt
ncV2Tub+6wgHAhQh+0fbqlyYK3C8MN68IUFYNGGoGwhqF2XV0HiYk/F3oIbspjql
v/BAHa4+Q3K6VoS39P6TBbU6tBezq2bdI3ouIZsxRQS4KJC4kgW6TGYBIU/MXwEJ
RqkWTTRg9qx0KMGo3+8WHY1cH8I8Z5aYKJQptcs3mA7t9Yn+82ox4bXWm426Kj2x
VcRvYrdGs4UTVLS+k9qugAWzFtwTbPb5YCuA8rhP82OnuKupbymvRMnIHSiv2BUA
C7ee6kCSyNUAbKdi7DcfMlME4nnnNjQqh5Lw4HTbhhcsA5/BoNoSrllpWcDtfXun
uNTiro2t0uWh7hiCHJfI8Jr7N0MWd3wrLNamakz6b0LO49OFvwteGLUT/69WWdzy
bO2h6fhFB0pctPMy22nuxPX3VrDdNf3XltAFoGqgu6IpqWewEeSHgZpTT0Xl3FkR
USeRSmAX05R7U78JRAUszJen6pBFhmfPiL3Zu8DV8igH7FdA2xm9V+4CrNHayiSW
01AwymeAdtx3C9V+b++BI1kXT1wsN/ynoCREy8aUC6EEzBIjtUCioBOtRMZEuPJB
Nhi5ElKfWuUbZIxdu8Sjfo5Yy+bCycIEAYfmpJtIxgghU+IDGUq/fddWosz4kmVI
9uQHD0wsgQZi+lrzl2fbGm5B7KSMuPNKD/kONZiqh+A5LmpYr377tSM2ihXXufQb
8UIy12Xi+y1+QcGylBgJCaMZTO2QLUxOQa0lFcdrPUkU0+g6FlJGi+jhrjKXDTZo
EbWunneqElqEceP2Hk8WcCnz7malYWCURY7d9pRanALELrjj9EJMc5pzgvTKmcjr
y0JlzAeOKPi5o/Zwu9JhmTOC0t/nfMYmLov05fLD6w4Rz8ohR9IcbXQ7TR8SUKQD
St4gcFogmBW+NUuhBePIUVktZrmM4KpMnDP9W4XYyeIC1ACgB0/bIO5kSCfpOhyy
yEtSaZ8qttzX5UqSHVe42fSxwPXYhp25SMlXoQJXjOd+mN2Xuk5EURNcTXiFnZCU
rP7gK5J8Hl9LdSFoJy4YUEerpKyGnUJhOpGbBBTY//yHJG/Kx0eIyduAulKDAyN/
WHiAk5EDIicMH/BfG9JIPB6hnVOpKI2Pylbf9PoyLh8zE2Xffpy/boxh0fN6SQ0M
KqC/LvoTuotXhtmTRIDcSsqCP3f4lKAq1PB0+vhSOsHDgbFn0al6wttIECyIGdgz
LfgBNEPazz/IE78quR0wRiCrZghXzokA9RRxmhOxY3r8HESK2tZkAy7G6LBGi5oJ
BdyO77daCCOZEkOf9IWfeQLVdDxwd5mioqHFF2nSeJ+QmZq+Vv4KCmh+ODshJaZW
cRtZ9h3qd1IAgRZRN1yggqUCNPfkGGs3I4Nxc5637rk5S2JiOk6uxiN/skQu9Eg5
/TLbmQh6kzwTGPBej23Js7Z8NFUbCaYbm3SSuc4jJv6oTlZa8KF6SZy4/WLwDTPc
nw8Ge0tCnzfxdfaH1r9rtmT8r1YfpOBAfPeQxUVQYexCq30Fsze7wOJfcElslrqK
2UNggNb19C0ZCgzz7vwWK8/iix6xYLUnOxfQtbKrIehqqNyrUM1FI7alyZ5eO8BI
8JB+ebaU+cithHN2AZDsJlLkv7jbVf4Vf+2eEoCHueB6NI/x6xkaWBMZozoWQ+mo
huNbYL/w0c77awJiCC7NNnS5tpxM84m6AsBgogZPokrH92JnJq5moipKX1q0nDHr
VhpUk00dTdZgDukMp7mAMxzdD2Yo7bJKQs7LBwoBeStvRNrHizkCbACfp8/UdvoG
T808l7Sc9bY+Ir311TJb4fwwfN/JQpBEUokUCsMCQRkQyjHuJjmUEovoAtof1ZRm
xFauLoerjptGWApnOIliy/V2sm8KNwdDoa2pNRT1M1YZazVGioiPUACaTjZ8Zgfi
y6sm+yflZ/ElCi+eiNWaS9wi01i5ayxMZd4xtWG55A/Bx6sMkkSmKGZH6ClJCH0i
P/DxX7shTmma8l1Y7fSdLFA3Av2iFb6OGqYDvKidPvfs8FV+/kF1rOb9LuGHSHII
8berMUxBnK25kO0lw8E9FzmKwNkuvi0G5rGSLhqfNQTxjMdcS5LdOCv/ZsKTwyIX
vmPy2rTroNquMDwW2ESCwUyGdjh4Fi6tOcS7Gbhdo37W3ts5pSG75zdcyAr3nHww
rYbPiQoUq+wQD7w9w/4Pd/5d3vYJDkMa3Nlx5e8INEz37ZbdUwR8WW6NHCAALawP
X/XZDMDYsh6mAaGcIIyY0CBsoQb+r2roxnFAqKlZqh0fupVj7BLYc8eyNaqSfi5Z
Dx1nTQFG1kbrQaklWX4OZtpAAQ1OkMbtevfBFb9RxZwduls1Begp1aHKlljJIIvx
PAwQwE3UiM2mJ81q6gdBeoQJjtRJt0tVWVtHSy/jwTha6vss2yN852oTBgp+wmVC
U5E5teeVAFD+qxG0XJGOLH+UoURG2+oogkj24LJM2zKky4X1ERqHMHw9l6NUt1jo
sbL3FHxXvUBNHgR7u3UxdBP/3d5btHk7rnt/0FeA/eks0b/5T1lJWHpJ2oR139M3
CWE8phJa6YfDMP7ukUt+wetGvK/TCIQmBaaoSPktowYeiG2wbdt4VH/Z3bLC4g8L
O8WW3/mHPVIqESaSHbO1cNXn2ZrJRm7ScoVbZLCrpwBjQEb3B/zhN7Wl8XntK7x6
6CNdV6gTkCiFN2SBr8fYf7mXJrl4RMNeCNCLNPoKYC5n22zN5XzUBrw3G+FEUZTg
Uizwd+snShRomLGjFq/e7uRd/Y6xoqAjBfkDf2lGzTgnpcP1DPnOYw7G9RDgGe0r
GoXLf4TDD8Loj/bQiRj79OtAsISQDQS4OALOxHSMgQVnKtDdfdO3s4bC65qRBcCk
OJBZanDZw1bcgGrG4kyu48bgs9VhjCqTsVTOMf0xVZB6qBMn4mQq/yXoB6Myg3bQ
hCbScR+S4prbLUbMErvwAPhbbWP5T6ADuIfHERJZTbCrqOFcXU2w9IB0W8mpmCWy
OZsheyR4JC1p/0UHjk+LPzZQwxUhh+rXpY1L2e9Kkuyy9bx5jUL4a9HOpRgS41tN
IRJCQOl0NG1ovJFukSe/CD+cDNhTkIexZekjeRF0eUczZWM+vb+ooBQzeGDq75EG
/kIOeWkSbQg4eUY9naDUN5YfNR2EwDYroXxR+nZcNZBXVpw6YNZn5d6HFb1c3tAK
rFJ0cpQR8wJZ0Tg9qjJK9p8Vr2zS63F3nE1eYYhhiRnMjDZwdrWqlImS74FM98lj
XNRGsada+hx0XfvNu3yDrtc0Tl8ecwufS6HCuKHaTtHkfmsyxB/VcXEkxoLu0OVG
exUHQqwhOcjlxvxnvJmfarV2BbQsuguN23EXBfGQphN5YHMFO4e1ulcwlA81pvTH
IH4iy3JI9EEOVjnxQ3Amzfw6/an/h91/GhcR4SiWcUxcMe6GQBBQ+SjndPCX3Q1R
xsF1hNdzyo+AmcMpoZKascvKaj2bVkPEYIJtnV8g9Cf2I66mgKWhJg7WcjOxwrhH
5aD94jPmzPU6YXrtKfRvw3ZMQ8KMDG2T0rqY5DC6H8G7prOI46mP++kTRX8ot67Y
S5wMGBIfJEjnawZuNN+J2uHQXSrbLERlqGdR1rZLSSo3hXgIP4pwBmNheIPrB3Ov
AWKrMpdRkjLSe6dZ2QAoxSbwq1qK+XNwW/RTHSYssirX88SvZSRDK7XGZVx+bGwK
nHz9lrLJApQkf86eU3VugQRLMkZPFVqmNni4uYrqQwcYC6lgrLDO8a+OW4OjtVHs
hAStZYl/z2F77hPlVsvxoDADwuj3BsFa9yI2EzU0sqjohfh65aLHgoDCfnBPwGIz
45uv0lPfpBlz6lG9ymtRGGnLQ2NpJq7FH7DL9SWH7x4HkmUsf+hVy8c916dmRO9b
xthr9qDUrVFgLxMT2bZ9z+A6cIMP99A4s0QpWU1Wv0XMGgxrjxQvuyrWxNVXqIwP
xf8vCYXfaJ8f70RVwgjRMzO/DU8sWeMdcPBD0hAPeqf0rxQdq4Ccy8QbqLTCMkV2
4z3TGYL0O2Q3TMROeAGAqpeqkwLMotHWFkeO1OVR5ll0BkVs/TVugFNVtXj2h5z7
LePHTe4e33K4sQEiJPUl2/gMrRa+DDXrMjk99rcXRORQDdVh/zbarOi9ZKEObzyF
iu6sCNAqr8SMgrD1aaiLhV+Ga5wC8GBk+W2SUukKC0LRbK7yZFT+DZr9F28zMklm
4fuLfsP3Y/U3KNNwf6eUxx5FI6+K1lti5jXYguy/GTlHxH8TGjobWTD0oa/7JMao
ksaj37+Mn8uH5y9dDrxMNb5GlHznJ93jSlfmOj5ny64qOMzn1KByckMgf5kF5Vok
5NXlIZALVIP42riJS6QCkO3zZg34ZZtTw3IEhIxyHqHfqj/FJpYXCxkiS2XxO03E
nx8URniUH1FDiXBzyktYXKvutkhq305LZkDfhtn6StzUPoEsomvFqtGvj6XM0VjM
p5h4JdJbehPk/1uh2noCTLD+t0bIPskzQrHtexj8WyITXpxLdcEaZJy853tnn8Px
u+PvBS15KW0nh/2y5Hb2blAub8v2V4aUCjsdHHwacod3tnXwAtDdd33XBYp4JTJI
BvS24dHr0qUvBntU9lOQVC6nsaWsJod1AZoj/394dxBGfD21gOgstmt5cnk7y9Pc
k6sAUsbT4PnWG3It4PRbrNkqIreyL1yu7RnANsKm59lNm7GCitM5FwRhGBoeohLU
snxxs4KisCdy/SaWvDKDpY0m0NGL3rkrolUj9UaTNVsY5I+WXOzxzKmXHmGd827o
rpRauLmkXAUHuKqnH9sfHwYWpcrAemV3TehbSud0ONSNbTPNmsoOQSEofns0fuDm
K0faUkh1y9Y0n/3ePB5Z9oDgHp5vs9dqQXspGBOUqrhUKFpjLVXgewCgK3gYCTTy
x2hOmCuh9qigooymIp8SdN2QJ0LmBh57Vr+f4GjH9SqAHfLQ2rHiFGGtR2CGWgYp
pXuTWravHy51Yoi6ngw0A5Vd9+Yw+wNMguN2gf4n1AFE8DfoA8uOSLMYVZPzKDQp
/oXRbnWdTvujViPEss/Vl9GBxI7+HUT2b1qtlM4Vj16V7AaDESEljE3MX2DHZSsu
wdNGh0OaPGlfLVJSsq4ciGegK75wZiazmkU2UOkCryORsCgQVpy/2oSUNJVNLdvn
b/gx/YRZPoCOnVKwQTSpO2EKiV9iZIk9Hx6zXrDN1i/LS9OfqHVez7LHF1ieY+Z2
RiELPBLV5PhTMRyAm54TzwL40eKHJacrd3SAxj9yGf0ZpyNK9LYKU2XXMuC/LaXF
SdaGY4bcoTLo8IGQ3Uithd10zNHzqKLQ/OSf1G92yBOR/iLCp/RWSbUIFgidvL4M
7DcKCTZV057HxlReJh1JEsliDryTp9jbpMZA8PZVfyyzvIqAIDGn+jkAhTO4Mp7g
2kjh1BjXObe3VN3lfAWWPY0FPMrOVvnfmSFf6+juciiseXO0le2NvSc4xk2b5m0W
2VhIq1DhM4pxhk391QH+3JwO/xl5oD4ZithvB6+WYqMZvUC9gL/DKzk+x6jv0QEn
PT039jzGO54UIBgm7hi9onuLR0oW7HANYcCmR7jjFwTrOkl1PKYL8WnlRU406Zdp
8I4qSKS4CqslzoRX5Z8i5MnZDzCJUQZihrRiCecT2DWyqIX6hJend7g2zdjrmVRZ
nCDfpEYxuTV/th5OvUscQwwgViSziz7j55saX47rB1sf/n3+ALSciHgKcSlSj408
iKNruaHjAat3zsoyid3nOvE84lYs42A09gVkE1g+Eg8ITNpjJ/1H34kVVfraZEqw
MXlVqYkn8LQqfxl/PwuzOQ==
`protect END_PROTECTED

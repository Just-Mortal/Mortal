`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lk5Ju1S/rz6nnhq8ha9CljtkPMyHG6W/0uuSJ1mW+zSqTh2DAw3l/S81/+IQ5sv9
imw7It4Gj11PbxH0oNwLwOy0V8Nb/+ZWi6MP3zG5oJM7dd4kFYvIVb2xnB2LD1X0
gUZVzUmByNi9jQiK75uYha6WG1BQEBsasmsToDzGAnLAV0igNJhiBXSFFi7xYy+v
sMYe2zNcvbjLBeugSbpkiKUIr6kn1WRPGljQocmbG6jwJEZGTF3KADHSIQ+/5crY
Q/KFpCo1MpefeGRORdmS4HnefIYJXunzAEqsxlCbJ4/kjGIBUDXQuD7LS2vwN2T0
qv2H7C5y0+VI0nTtmqI6uhpx2g/DXdd0I7Cm8s6AXwijm1cCxY6Wc0tlH8aw2iUv
XE5dAqIzJ4pw3INXUfEZ1O9MoUgq32knlmNXgx+U89qRsv/fTVG/cIG1X2ArMjMg
cX/VP5JzpULpRYh0dZbLgU3p4ubUjjnxHI2mfwZ/itO5++YYNu+2lb3uwachgq+L
Y9+edJA/zNf32cgjVs7+N/+ci1OiqHZCGmBYUQTU3hVrsow3XIo6Yx5sawagzSyY
NLI1BJs3EkxAixdt1EMoIUWtY5PK9uQQ50Z3EXepSEreLt3otb6MLtjRi3QpMn80
qv2PThUMbeJdlMoW31VjUJ2I2CnCSggqNJo2Micm/gYFOb9DiXzm/f/s3+9nx4WM
albAUo1zQ8C73N9lICLgUy9AsvongVMZ4w4tLZn8RnsDPNDnzZGjHmRhAjyKTWcs
n73FMWrUnSE1RetHW34EJAEhMUhVgv9uTswllBvhDbZPpGTmCyPtrjpFUXvMQ5Gz
lIKswWI9rWUcMdq1oFn9/a2ATNJ+vJ+reKW+VIhzeFMyvJYQpy9Kz/RvlDxRgP8U
86swIBIcvMaRNvdSCtEjWKttVH8eZ4uxiAHy1I1H9hdkU2hdHhMOzYi6EyRFrT5p
CUq/Ul316ROmfyluOpfxsejkWYwGRWdLGoQqJ38+fkloUKnLWSKlzQ0Tflm8rg4c
Unv2GAVaOnv2OZSrYxiOs9+Ly8VjF3Z6oVrDoBSFAFgRb8YfQ8YCKotGbE3/KNz6
u4itl4ZR8w7cpvaz4nMi9PZaAvEEznNJRRlMnvFQE8nDNZFrmMuOGpS+kSqbbtei
eK+CgjtSHcZ/sTf4QC7fO3PaTGktvyzPyIN9w5mqRxQTcvVuyorzcXtS6aqRBNL/
LOlrs+yUwCvTOmhNPfBNri/wneHjA1plw/6yk6GvoIwQ/hKqmJ896HkBvf7DbVhh
OAtETHv34IN2GETxTCUORu2RSEVyA1nABNEnKbeso96hfxMo/M8hGWh0p/K0/Yrd
bMnQ8fhDPnXUeuB8k54g6GpmWEzVLEOtDbO6O9shGPIMn7P/AK7XDR+7goHkjpFH
KrtSGSBL1fjys/FumJgcLy2NyZ791DQw6BYLlTjKprEKO6uLIz0bmmSW9rA6Jghq
grBSKqfhm1SizrtKlNBVCsNut35k3XEFlWclQmOjAFRI47Qlc+z1SeYe6HEwVWG9
NSi4/rIIbA49GfwzgEE5hW69UI9omZROLtNjzGcMm3aIT7vRF11vvkal+B2nF7yH
F3AQxGABLIE2cuuZRZo4s/J3hsUH6LNnqUC2hPXUvEIeEK30mpYfsM0ZOZE59Ctk
gR1Xmvgl25gkllvyZvG0Pk9yECNH6ILOjT2SLo+1X9GRvlp+kf3/PL82kxDlA3zt
L6ZXhDHz8ewvE39fZN1GUW28Yca3rhkdePqGZIdV0srYFx/i/c8Vt/C3I+27Ptap
RTVGLwNoblpwr4YQcGlnHoqJnRQVEJhlXSkKvcRqDkbthNI0TSrWvgpevjJYW+Zm
x3j9q6uW9GcCqFfCLN2yx5hwyXO3dbu11X8waLvo4UOBJHIHBVHl8B26Vi+HvxXq
ZNUfUhkP9qfqikMocgK0tdYF0p0EqgMNr7+DbAl6oL+5Qd/1EUdzOz5pjk30VtrF
lpd7oCWco3dq046q15axDZVeKnrGVGIbtj1Jy3HnQoPSqa+tMieIaUal1zy17soU
Jm15CV6Tt9gnOksFV/3K/3PLEHnnoq7HcLSCAtzpFr4MgyYjVAbGhCnuNoPvz60E
aVGFeQi8eBj9ca+tomblZU4UeFa4AJNUiMMWSTPpI5K7WhjwF2gzPT8myugpDUKF
2EPAVJkkUf2SsV1DEOuEX9jMDM5N/ZWV0K6IczjHRzqG5FIHniZMr/7X1Nd8Pg9l
js/DwM/9jS6pIh+WIVAfVgX8ais785QpZ10L40FeXODcbvqV3qlnnnlgXqjHbhDi
NsY7iZGv9qJ2gmU6Qf8Ju/D9TZ8QKm3Afi5FIODaEAKRCu4ByWHOta/u5dGl4+tR
l52b179fdFYhbk0JST4ozYT4jxrUBlv9FA26fxGIDu4g4xjaa9zXLI8jx5ROlTwF
aIrY1+DfshG9b/IozOKObgKJNWMmAeFAN0OdiEs+I+6Sg80HuqkM/EgrDL2CUK8b
HUYLPasfTYZAcxYpK7iGDkHC3Uj0PNtrOE4Qvl4ko3guhfbBJqwsmotJ4IHJcZ9q
V45U8109FZ/RhlO7m3bBMTw3cWqMJgd+EsNYfB72MfENH5ZzjfuB9CB9kDGHmN0Y
1YI786g6unK/4a9c5lUfI2PPjkBx9CmR3x+uOTn3HyL2MnWP/3AizwmybeTqtVYS
ATD6Rf0L3Dj6nUg3WQg5LnwgB54jYdIHix66h56iWSYhega6ANaRBrK9XdSdik5M
Ixn/upE3aC8hz64hkot5nHZMyzppKGwQbF1vACAOZwGLolxkLPbcJNEm7Gy7tYpE
voyfifi0uhDgdJg4JTeYtBwktVIxKyC55mUVoPEQEypNkaWySiEzQjFg7R+2h8L+
p0/zPo7FJgpboeRMOVHJQquHVArho/8tGskMyGkaRkROKpgXqjIRbYbzAXiMKT0R
ff3BbN1M95bqjSYZNY23fOTaYPGBpHdtrkh2ttHIU+PxwzEICpRvdx4m/8yiWftd
DynwYMGHiPwbQ0g83Fbr/UDr2p3SQDB1M1Ied9NAI0xHCus3c2UMTLTptk5blGLO
MQeSqVQQBqqprefzk5RpXIe0295Roa7AF2E00kA6m6eSOsdRAsUF7CP8fRCZfSVO
qkO5Ug2R5PkC//o2SDoTD6B7DD9DxE3lvdMKRGAC2X6rEQWyqSEOMWF5o1vmHPfK
c8/oO0RN2kKoFc+9Yc6dElmTDnNBoJCzrFHO4bv0ow0uJW9Ry1mheQr+s6Q9cD2X
TDjgdnM39I3yMWmu1OLly/7kS+nTLu25TXUZ08/y/K8t1eynC8H1fjC1SetxxH0z
DNBSSJO0fNb0IAIlqLFRrwDj0eKcWxuhjsEoWiHDOOZDm77yrbILZHfHjQTEjbN9
cqUR2mVHsn5ClnI9c1QEnWGvXnULzHShJbZQ8OQ+NUUVQ7aNrlj6SIs5lMFE5YWl
5PkzkNDqYUyuhif5p8Q6q2YGR00SjYLGJMKy4tFedKiePc/Y3XpWDFras+eAnKai
pma0JJz9Rac3/UPptnmEbXlhh3HNZyfZHp0jJofV3lTfpUVWboIXy8HU9mwh4gOO
M8k/Mri7ArUuObj3SVwBM/r5D2VloHOpeohHd9EkYYFm8+VH8AUcL4BS7LS92jhq
f/QWNLSoFVbpizuG4P6TZa5jUeFwH8hiViH7fw3Eq1viyWFvjjN5/EJrbdfiRW6K
DNJcQp8O67OkA6nOzHnAs/NK+obJ2OtYyRjyDk3kJZgaARYD1/CNyR2p0oy7YGXc
/mPXttQDFckX7xYAp3vQg5VCZBkteHPe6kcA+Ut9Dr3tKUksu0pEIl1ZjiGC184o
cv9zVD8bze51KZs4jyvqREWEl+Qan/jQPagih+QLpUSwrnUhvruYd7KwDPp9zVtK
1pbvBx9r7NWxH1ORkXmWOe1npMzruUGN8oR+xRfsRoQ9JMa6c/td+4zgaenEQlcy
urn1jrTUFt1JhEI4ThqrHWrzq+PKfEf4o2E4otGrpytTJJyoH3Lr751cwoyXlD4g
v2yJM6Rg9CLOMnacaIO9BLNO2FzBwrbfyns0+YloG0gCiupTG1iKOH6kC5gNgaYN
TMLeJUo3DfkA++ZURxMwmLcDZmox2E4iJi7TUkIJ1bAWeT8MZEp6VRXSlNbPrH88
wP1DOTi1RWw+kM2ie78/AsVWlQRfD7zKCimEc6rktvcA7uFchgPrjsT6E1t7kl6c
NSikZhkQCZwXP/zer1sNfpXhJ+VeP+t4EJ3VUdffvryg8aE6vS4PlCI+pzsrnJ/2
FOPqfV7Ul0+OAnPkQbC8rwiJSaB91MKM4MXU/hftMqknfGMS7AQDI32XhJbBwyrC
b4D8UPb/mFeTBmVANtkJXcAibelv2zwyiKjZSrhZrularTNaQb2JeJSs4D1tqQRZ
lKK6SoEJqzXvtTY+ijvd+t2IyKiVzcRA28bzAQAJuCdeo5AzYPGipOCJhVXJ0LWk
j2gGTPZhXqUL2LG9NXTv4gcw13QVRl69/tNG85/Ypyfjlont+1SjwjzpxwjuSkMX
A30XTt2Cu2PVJ7abyflf7nBkJqKV1dGQErgW/1ltAUz+Udy2GUlESy5YJ+oPaQek
ogyMfMzdnuBYa1+CQdTIxjKcIt4AmHXLvAY8+rNKaDctwo6xoidiY6KAvC0nvRAH
rkkW2uMVvZu7eYdSqqd7Et/L8k4YsV+xQL0UdEVDh6/otC5mw0tJDxt7NZwRUT6i
iCtsl7ZmvrcmVNca3EFjR5w0U8z0I1P9wQ7xK+li9XTnz2klNOTQVkxCtSFT4MQN
0I2UtL9wEmaUCwqY123ngIfKlipodODtw6cKYmkw6JIRDJVVEKl8YX8xx2FaObEf
8+T0M+XW/UNNPSFuHNGHk59UnToKnJsOOryAo5I6Uxx00/TA5q/63ttL5SBMxQFC
8yBn884rL6TnoCJzB/KIsnXeQk21fTfVSZohZmopp4gpVm5gTMLEtgGS6mpS2wZ8
9prfv3SFb4XLqGbNA2fBzdEkJ4mCjIodKN/ZJjD9+ewzb5fvSPlSE4kCESKxr9iG
wNvtZkodyG1kfmzLS2baBOJ3DC92Y0oapbti/cxhPgsbpNNAd7TKCUPead3EIRtc
0p/PKx6GaH/MqHHvbTlef6lO+8l//jg3B/KvF0viLDmSGIl5x53kPgyHLD9qB/+x
WqtrgLbMkThkwhi4bt/8sekXg89Y2lbi+/PwGQsBbEEQrrBdQGlwObffvGnBLiD0
9rlqJTl04acwrNqM1e5dLo7Leiq2zO6zdW7cp+yyymJPnC0XmbopXv8tcEBc6R7D
tLpP+EkeekzbSPOlOn4EUJx4HMPMCHYNBeBXC4StdguOUyg8OUqbiJNUuuIYAh37
oeAKP61v2xDtlDE4L69dcoFt1BmLdvC9SqAaYCqU3W8y34VSBOYfOxcylqACWmq6
fN8x2XXCmdIeqO+otrVYSedl/mM58U+WODyDxxqGHRzILPyumCXBOJBLCpu7ueZm
7Agt1rkEk9DOutIbsHP0ZhumQMn1ZvXiEbAkfDA5mW0VQre9smV9ULPMqKXmtqjJ
1+K1B9O6/inCutTyIPQSM7TBxLaLfNhEIIWY+jE678JOcGbuAT6D+ycCEW+SCp0g
qfiwfRhFNezyafewkczWvGk/g6vDX+Z4qrfUtzEm9q5ZxcKd9iAeZpLOf/55gzFo
qPSgGPa0xFybZj8FbrNkoSn6uO32vs69/wvsyP2t4V+KXiTQi+0impOmDiXJ8fDI
KNgQPUfvgiazHf3AApF4lpTHg2m8MAz6uepTCstIe2ilwlKgErkNrB2V17ZMLf3U
S93Bg6MMTcSlyklJW5aYt48F0LC48+tSoOH2fy9fyAMUUJjRY0UPycN/jCdkyVpv
bxmM4pyNraDCYc+cyz6AqVBggERe/hx1tgOgk/09kRvv/TFgyhl7AEZcb+fi8K+D
3z9TeiEWa4P4Hysbk80oCQQOYzSDdrLs5uAXz2zejpoRvLijOlLco1dbnNCu97Vm
LKYYMXtKaLU+yCT0xxQBeaNTfrSkPqnaH7SRISrx1Yxhc54wrljlnkcYuqBQGhUH
+Z8wGxOM20hqj9HDrvfkI/PqHI7r+kvw4+BNLYx/51+QIqoEl8EN3VGSYfIu8uXP
OsDLAwL59kI5gi9F0LP0g/1FIQLm/r5rWiJR3D/ERCBsuAzgiT/XBmEXosQWjZnJ
d7lZqqeo/Oupo4ABWHPfbi2P5ZeQ8dS/zADeeoMtPmg6YC/uBcn8fSBDFwFJEwYk
uSNqaOspTqxKyWrNsHkbvNLOnT9aamf3hhaHZ3af3n50WC9dA4KSaRZsJN3662pI
oVd0lvqob9IZcdOUbO3HxXZ3iJjqsmATZE/pSy4BdIJAUVGNa+QG32b+w4s34+h6
Gh8hJnhNijIp+YghKyQvw7WhY3V1yWjn0sLs37VNaIzqsA95UDftTmu6Lx24RHdM
ZY/ZH1xwt4HwuD932WgUp0vlCV68MRy2wjmLzWYpBwyjgQ0Trx1UE9UdDsfhwqQ1
rT5V+B6nEsunasaSbPqaGrw8VU31cAxfo5OoyLtaBhMX1c9rx9fWNKQWF42fBZIm
OBsWf+4USyOJDrCcV/j89IlXrILWbwVDW/AFA0qNSqXg9u+kZ6rjB/qhl24JOWbF
8iEdAgsCwcCHISw/ElsPvk2OBcpAOH/ZKpOTAUH89DCWium/FD8YOm0fDC9YXoj6
/nHN/K7ybWiU+0MmQdjfo0Reqj8YanHPkMn2sUtefIjWZ6WvMwEa6h4TwyTghFsE
oNZzyELtu8t9w/pH16mjjrsOs39QrR4pCNlYzUVaZQD8jLA+wLdB25LRBHNV5G3V
LED57daDXRzDgCIZlihblHRpacnJvGZ32SGOR606440Due7RG6YDG8V6vnHH2LHn
DocggfzQKXVIeqjswFTFcO+OIE/dIySRKlpKJMo9oWaSglFNFEHrFPmQuNqrCihM
wMDXiu/MqBTzqW0sUUrMYS9H1y8ST3ASppR2dxc54uJv+CjbAo0FN9+WQAqG3e1x
pNbW+JgVAkHVFBdBk9L3WNfGdYM74pB417titNXcTvOLvn1Lj9FRrgxXfe3/TN+j
420pE5Jr9qf/OvQ/+ehls3CLc1eTAuLkxhZEy5vN4waXS/UKO1FYzufGojJ2yjyE
fSepG9VDC1bTaf7AP1+0XwbTnUWPIi3JEOm7pEXuT8FIjWIoHsNcNOWL95qkTioi
W+Ls8mIoI2dIV7ZKRcxu7SzVRu6AMjxdE/g4wtIWAZ0+lqAvjI1PcVxdRUFeoKLO
H7z4wOjjTA9fOs0LnlFW7DfjRnSry5zGVHNTZDz+9Y21S9BfXHSVMYFX40uDa0za
Q5B0kYg4i19NHWi9czlAUeJKL0q+1lDHc1ekgqVmNo3+SBwyvm00Gd6gPx47JQ76
GrfbiYQaqOCz+dQNEpqPTQw332ydJRfPbNCglgcGY/JZ8riCipvdPysleYEoxZ56
z8P2tXrymDACTRYK0OPQeO657R4xzrBQa2eRoD5biUWiGfZAckTOQj3ltuK4S8eO
KW7W8mrElYrr0Ww9r6hIImTEUQoQDwG5c/1qPuqGioJmiew6Tq9X0i8RMNjlnVG3
ousAM1lzikvKFOHMoKamYK6R8rIbCC940N/OIwBxN/P58ky3NyqYcLFmy5pnbYEA
TJfHIXCgK65vxtQ8eCR4wfCQB/NZ7BO9eEkECrE3LjDClJse9iOBUCcHHOFD8ykU
iESfZUFuUfvKJyF3ffpqO/lSjMo+K+Wz0xJniANvgPHeh/z3v4Xkvzze4cuTN+WI
g0eNQXw6l8X1mh/hwXSJvP7IB6MYXrxplxt4/0FK3tW6i0EuuzH34oAZtHjY9u14
T+aItn8lUjWd1FouTotm6mu1k5ZbOUNCyU7nGgjKL+sCOOdBhUwy6A1vAKb+AlUn
E5CMwbiYYvSq1CnmZTtCOc5XEZTRH54mRXG0nqoMQFOroamZ5hYqoQfpF+bliZj6
xW+gzEPFJEFRkZYeHp0LW0ASwJfbrAvNNDqYPk2S4d9EiNQGjSYqf3lh70/0v6ot
kKxVeOAqelLRurzGZX5HUVSUvoUvyR70yZzqvNswwkA4Kfve/GlHrOdXwaejk8eC
ydlxGnK2ox+D2B6PuRwNiCxL3I4ut0ajFik22ywa823TSKaj2GpBaor7VdGwEFHx
rEbrLlv+K2a9aUozYYePCG4uJrFj73WJ4+W5IkAmFHm9lCDSDL1C88j8aSw47wQw
VW2eAe+Iu/qJaSvoBhcSNEAoTIFBeJom5AN/DmmXFcSWJVESkGF77D5ramn3cu44
PohPhnff9rOmtjoBirkOeZOWP8fBBF7X3r2pUViC5FEwoMyudgwR7PtYgNNJ9whq
O29+TUIY4ATcbJllBfq43GUjvN/QCwhDquw1kuMr7QUgZAbuFo/xHqABhA3eN+/q
DAm3CexwseT5YTH6S2Rv9LX3MuthDK5dRczBppZgiLMTkadkByaVeiob9PqhaLFU
PmVF2jtvySwCrX328ccVpVYcfghgt0pde4SuhLXZoNzbTdK0y6U0c5izpf2uTYw1
L3Ox/LRSeUB/bZbeWcgHy/jQR0Pn8pRMJXNepwG6KObALTH6AEctx5JZZbMF74nj
AwKL/2DGy3m4mynznUzK48/kk/CfP1UbphArTG09cBSSlDiksfRZbDabQG2gJFs8
GrNbqovctKUEiKZ46W5U4HeRX0iO8pT3wmqHj6oEHpj8H629ctsorDc2DoQXXGLJ
hd//pa+VLedyiovxxqowKUr95iaH4cgsZeTYNCY1wWbuura62trNnE3GMk5Gc0X3
pn4TyWHYGz+Jw5UdbjEKERZhRnkAX6ScMeVGW2v4FAo/fxDTXqFyIdo66GVj2ztp
qXml7I6IhdxyeE7JsVKeIP6A/dtimK9troDXZK7UdV20D8+0ri6UmS+/xvYK+iCe
HjTGgA7F4HDD4yR/sL7XUx04KeK3kWiT/xi0zicBdBicuGiKPhn2Fg7WhlsBQC0q
93NUgKa5qYlGyi5NQR5C5quiU6IoJxiL+XAy0myNjc/P1fIC7+YiNlcrRYSLuVWb
cp8mV/y39F50KghspRo1/4slLLxURvem8YvRHDn3W/3PCCrmPzWEjyJW3YQZK3ak
l0YfJlxY7TVIapdgd5ZHxV7i+GwRzJAkRPniVo46CSU9N/3YQPnPYaNkLczCI1Ph
jnW8bLQ3dj/d7PEJjmEkOlNV74TXqp1ae7rM02V+p5DGXpoNaHbVMaTI9026zjl4
SyZUCPYfgWDQwfKFPpxqjliCNAo7ZvkIIYvd3efIw0YXLvMP5BYZhPRtvYQEs4PR
XW5SPkQePuIhWlnTj66cvJbGEjXfSGXWedJwmfd4qsI/E21hG/JkRQFMcg4sKcYX
mTG3csFWcI77Wi1TsBWfVyNl5AOQUYSqFbxSO/dw/O3PV7ZCa6ZTXyGqdh9stY1a
vHNUgZuFkp9uh6oV2f7t4D4XyxPDV7p6NwtYDqIG6PuqqNKMkGcQhcxp+IHOPK4e
t0JyMQSm81TjgfvURBRXIKbMIEtjkITBmHWwl942nYn/1RhheJvsLxOYgFcYEnI3
n9FMAFgGYQssoK42QFmejdKNWKr/P5JosZLJ+FTFfDxsJhXxyN/uLTalGOV0JErz
MWPDarDyU5Lf54tTgJfT/2QVYfo7Kt157deSxLVxpDu/dhmK1CzX8Ddzbh9M6jcM
rGL/CiKBMA5BG/gf+uCRlYsyYvrXfeIJh/fskryWNevP4lD9xkaLSQbVx0lxKWxz
ISjaw29c8lsCPr/wdwNJ4uRho1A1s9mLImAWaQZybO657i3M0LQUywhFzwxblcZu
7/vMnldY1RzfVJDK6NCp3IV9q5h+GLMzLKTC7iSI0kYsEHOQ+/raRAaJgPRma++3
xWoiPZjrD8jKN9MAUpzSKsA5jcEkQOCPqxMPOPswLLFsBmlS+SCIe5KjFBevjt92
0ecWI6RpnZosgVfUxCkh26xFnn/aCFybuneqtfk16gMm7DeGV3XRK351WSLRWvDg
iTXilVtsOhjCMrAoQ9lqXNvxn31d3/s7RlQdmfDfxMymfnNnPwjkvpS4XpErAyi2
pusq8IBRl8kkjbt2ZEZnNIjctcfyltK9Vpl9xGkOoYqsrPYsW3MRAOJn8cc2pGUj
fwcE7RUnbIAnJFAxg1thODuhPNyPamfPE0e2WDPk/u8addiD64AYeAqPEKdrOVNG
XWE50v37W5k9kT6Yg/+PkiZy8q2Jg8Ou2b964FHWf3mjgZ8i0a5YdRBfcppjdbU+
/hNatsZuJl0HP+0ZmvltJ6KriCYWDyF6uRlBijn3ZU7c3gY+QCnbosLxRrOGZH2F
uD1A62wySTCq6HJUSN5PR3GeNHVt0fSE32Cpcrq8Ztc10kIFgPWQqo2ubyZ2GbWN
k5rekxOC5MgxvjnDxKcU5jIc12NC5u2x23/wn2EKCLTpCmVmUANid33d7qwEzT1l
NcP5W+VzcDBOtE/cmPoQyzH+81UAZJkzAC2txvNAdAJY/qaI+VfgSKKDd8oDw2mP
gkaFXrwBSE+AsnTVfD7mn5+hb3sEBEH1tdUegqMqx21a9QJr3J7jF6f0bTN19qrA
Mgja2SdKZLTQMU9unyi+KZUV/SBsGnzCbT+aW2hdChDRg/PEXDJybJtYtbMb9Lqy
jGs/XDYy1UpL/x7j8wfRgKH8JkhzV/3/6eUtJZ8CTQNJy1PmUu+wqoViEa0bmmdq
FUpEu5xbaFj87PnoZN1S3aIlKOqUhFHOiPC5u6/Gl0IiUeKO5hajoMIsuiPdRYsc
22j55iw/rj6rOzQBLNTMZHZYuSL1wqkp3lf6EhZO57qUnVYw3odCxzUmGsZYPDB0
J7yZnitU62+mPh4xCNIDBaKkukrOBPYJN8A7myd/Zd2vGOm+Q3fEVYKuWk/vi1fx
CpPFJ8YthFWktWZoajP3zZbymJoBGqIL2ty3Rve3dNTnpQhNfnNMcFh5maujkAy/
ZOAxn1YPPoaze4QL+7/NcH8qj78PiVaIhVtDJRTrbMgs2aOljPWOQDKDIpkaipRP
bJjkRI4fBsa0U9REcMTSM9JD3J/lRzt8+Tsq8QkMLVvB/hJb8+AD389s375JHKnO
Xotf8IqSXv+Avs3qGkOd/C8I8QWi5Bw4x52cGTMyjN5eZ3XoJ+5KQ/L8j9WSOz0w
SX6/jsKUzZh72S6xNjIaLRCH7YeHzfpmZsEz2OCMgVnX26eYKqR/SPxb/HEkHb8p
JIWgHO+lQdbK3ZgUkqhy4IurIuC/0dYB6ZosNQ7xHNYRW6BfEsgjSpbYtFqfWF/x
I05ok9keNl3XO4ioqkajEgJeYC59G+ryWq6FdK7w6JN1mNro65sdLJpLXPJDaAXn
zBM3Uqxv2LNuHLUgDJ4VBFkbhvnFQQtRAb8+TJ00uFsCgMH7u1RI3/kmF43dnhxq
vnozILLr2FtmW/jC0ZZDNn3sYRai4GOMqiGu6SQ3A2VhySCdYpd1+J+mLDsDBPEZ
ib2js7C3NVfP0R8KExFgTIYibQXzzRnLfi6Hlyu/WiRGpbnBA1tB5jUN26Sb0Ulx
nNgy1C/whDJ+P1qUQbriHGm4WisLmcll0O1qjrmNAqzWI5hyquZaBDB8DiB7GDql
N3pXLW0osRjQd+f6Ee5+ouQzxLZAM3Z357tMoHs6P1pLBCpKKA20tshuxsYf8K+4
s3MjjUX0oBrLXxD9+0B+iJXl3TzKbSIU1e2hWGihOUcyfGMVixtkOQY7Mvb9bxWa
jcZWAJ0HxQfLj27ZJZ4jzPEGkd0nQlimIB8gLwN09I8jbOPNPHS1YcKy2uB47j2z
8AOcekf85n53IzUu7ZAyEO7+3p3jMAkLDf1W9p1P997AZYoD1YVgBjdGt/nQ7siJ
/qs5OVLEh1w6rN4NqMVvEHQp1Zf3nGeYE6OJf6bxt1Y4dbL3QJbPs+X0vCQCEt+7
Gifc6AhpbsLkuC/3gS61iXkpIUmGObI1wZGzieBC+0LnENieHth6f8NtD49d50DU
ipNnzOWVFX7zRW+4Eu2b+E1BgfL7fLhfSBFVIzgZh2QgJzDbxmJ0uEsZDroJ5QJq
TrdoXB889TqHWqvh3aHbgGR5jHTsEscAq2Yh14bu9xi+WDYN8miRHt/mP3ZwgriW
j0SQp0pHd7o+e25gl9EcVhEzf51KRLlp3hC+wMzXNdu/9Q+KyQnCFfUTeNv8zWtx
f6JdMFLeYdRLcaj/zwmg+c/0gVJDWQlhHYKMd3Woka770qVitNzQogn/s+eULPIq
0Jasi0iOcnJNc5Cnn5OYjL/DrnE/GlsET0h3MC3E40UFcEcULWg2cHoqhs8hz6M2
CQjS0kEi7zacXBgATCUsRvoCUnRL9fqUoMOYFD4dWLlXWM66zXtz4jOF5BmHvift
MW0GTFtgjz4Bt9IlDJbI53YWiDRn+LeIcASjaR2YHBQ2RQJbCXMofuo+RgOxdb8N
mLZmjHcI36kqJk5pCiWUo2j5CmwNlNhjNYSuK07MFZGg0pwIc8nXkAvck4LNg+Cf
Mnpgo82xV5/FoSTXdi9wUphe1lmlgiGR9E5uj4+7mmtwqHcUaQhG1ibjcydXZUS4
/AATU5mirZXSOlxf1Ygf3FH8UWJWXanOA8O+XMnGtVAAw6HLMXbPpjgShX9mdj17
NqR0mtJOUq2Ksi7khFGCW6Daj/Ao6QwBPtyS9awVgmCUYzNRPNXKe35l0sVr85Pp
6QzQwBahGETr99NvPNsZ/zkhvRo/V8fOUm02BAFnbVkykmDwIemDilabakp1BPFy
6Jkdn44pmAxd/5JOnaCMZJOIOYzZrQDU+O/Ymqjl911vKSNcxabu6y8RUL90kS30
9exiaSRE/x5ftjP5N0gYwATeIQUpwqqIZDInS2Y+xAeRy1pZYxGUlJods3JMaxP9
U/DvrFs7WxhoAZ2oeRu7vLQx7SgIdi2FAJuI+/ecZSuG3laZ0+0ZG1vbV7brPyim
NcF+WKSsSvXTCeHwlA2GhmEpLJoRZLze5Me+1d2ybKUI61jHLXBYzdezsbzpZh4I
dhvUvqUnGEAfRs1vOBUypKnqgSrQpysUW//utY+ehZ5hXZnzOJvFoi/MllXFutzY
XTS4nBLAkyLuqH/kMh/PiuY8F2kDZf8ObPDvs6iM9zws6A00HBRBKBth9VJDwd49
7CPlRFeD79/plXvPeATSPQvp+K2sWtSFtkeasZVzksiYmqrilo30sby3C22tAXFM
XST1xG4p58f+wgNi9YAKdDtW37DBf77e9ZClpT4gxwHjLOWNQ9H67T+8AZ5j7zx2
rmBXQvIBoE0DRRL0+935MLa6lDByOExXzLIau2Od7190aqXAz6VHbflIhZUtScod
/IXmJEu2w6F3ROfACbPwX9LJ3mg1DaLWNQN4+FbiIiV9uQ5RSLeqPxIe2RZVS521
mELL0v8mbcfoZY/qP0Fnf8lL2TxQMvFpV9HbF+9xzcdMmGJhTOP8jfUeoTQMhOh7
7wt6nhEosOCtmG/LMDWEm2+tTkqeJ231EMsGeRyGDd4nQlMEm0HfbGpN4JYv9+9Y
5w86kcDk8ygu9C2uDORfnTzg2sCI34ZgSJm2thtK9ZIuQyDaJqLzgBdrElkcgSeG
b6NLTzbbyKJq+LwZDG+cUfqSUeyNGnxvj+yzQiE7f37/FmGDiHBOxo49SpPPQTmH
I80PwMYe3sPSgZF0gDKBnVtGD9ySqgprV/vpGkpIJXyPA3SVCZgEwLu3ArcTA+93
nXpKOYtJytenWTYzTaxQUwkIGEksEsxjiJnkPVKGWC4zpDJdxsJlPL4UR0+EOwn0
eOH5DdF6CLtD/IwPmsiN1KvRdb0eDV5CI1s4EsB96RGZ/cT1Ssr+wsfS5mX/KhDT
ngnRhbA1R2FOd92vRRg4rrw/tInmlBw+QS+bdAgxuqIXTHJSbWoTiepi18o2SHhJ
4P/9e1w0aw9Zc/wyQXHxg1UaY1biFgQcyejVbFBBRkPhErL7cUpUicsrUnIoE+sP
eUZ0VNfnhb8PO1TB2mu6kTMs9nEnuS7hYkiXNMR/6PqZBofysaC4JcERK4WSTu9M
o5LwKYP9oHP1qeF/yzfc+6Pr1LaiE8PXF0OD2LMR5hoN3C4jN0UvZ5AwhCJQGaeQ
sJN82FNSHZuv5KDp2e9jZEztQioi5c0taU/M8hz4EzJZq6iJ86OTcI32I/3lP/a2
IjVlhNUEMdjwfyIPm9HLfEI66o0wfiKPAQKJ8myBlbw2GRefjn569RD+VXOz6voc
MTWZX8Nu6xJZ4JFR51Ng0n1ju3Rwl8/qwsC3l0G/LYmMeU4K4xOjGQdlq4WZu9TE
E1lNjalG4bhUsP/s0ukCNo8x9d/SAlU3PhBaWECYsT4zsAq/NWpfNDvN2JclUr1D
Uysnm14pJWkA3HgfD8+7zp/yYgkINxNTc+GBp8v8/yLvOXoxAkG5zCoqlMMfEnXh
RFDRnUabce3C6+UUS2mb7ZpUfD7Q0gU960mzvkfgnpXfRxX8gGa6EM/84hs3ePOu
uBfUWVu0jJGKRvyOF3XfJK7kTz1wVklTvuIrGJZBUXPII9wTpqFSRvue60K9GEvD
KM7X9ruk8FYgiFaJkr5eUB0rwFIl/KTDmFCMMCRglQiF79v4Bhpu+QqXkbvOScHb
6GtkKHVAp8zyBUzidytIua9lzVDt0fJ/x5/KTPOYvptlq5Fm3EXVqDrgywbodQMp
a+b6KmAoYBexS+2fegH7jFk7WgUCl0N+4gNB8iRAMyuZ7pfSJAydBJ5BPcE/ttGb
GdFLXxiPctd20yxN5woj89nw5Tm6fQjsZBJ/fbb4QU91+Z9gSIS9sXWuoLvVKndY
JxdXtwGTHMEk+Uuf+DL2gmZ9sbYtzqUik6uDx6kdq9TOk/VyVWSGCaRIk0yzPQXC
ZCltMfeiTTWhlmSUS9yzQEtMDpeb9N1INMYS//2nIxa2S0+xQttvH47e3lmmqHPq
6WPiXtx5771iUV2lPik8F4blY/gtvFmUc0QE1qkzui6Z3LG+2X1VCEpJvy9KQ+7Y
VNfO0/1DvuH1MllQJqYwt4dR6Por3BZi132nspTDVVP9JL/eG4z5zK7NFhOwupnT
j4bmf+wb9czU8bS8Q5gy3S2o/IgZzwTxHY+RvTEQehHwNsov3tvy/VjqtW+bbOco
hUTIP+IYh9yjDZqrcAzBkn2prBIG1Tc1pGCzLvXXPoZkDiSJMGY5xfTQ7bezJNU5
dbp4Wo4xUqZEQHCPqclraHz6EVvhg1TWt7XuAq5zNCk68yheMg3DFt9Y09hPgDrQ
0rbYbSGUt77uPShKA/u2U2dyTgX/YZDrcSlv/VSlZWgwCgVHXm+23+cdJAlBHNDf
QmwLhetczI2q2d07IS5JCcz3RhOGa9X8nuwkiz8VELXzyt6Kvr7y6gNLZePcdn0F
SBdAkA9rInvV4I6nIw7UCI2TQ/Azswjm3aYX2C4uWp2aZgjLzT9mN//sQw+MBExL
40PEVHHmcBC5R5IMFSTYxi6KwVe80+xZ9zpewPNbAxxUnWBaNQyKkhzRxVMre/I0
iNHRJ4j0+u1pl2k4wfEBllWvPAwQLozz7vaXIDRS3SbH2EgUCsz40OiFASQCraXV
iz2VswbGzUJHQbSXwP6hU/ivTa6kX2RbeecbGoKEfJVYdyHhF4lw1N9V2C3ERzXR
CHE0xs/LWCe4fYOUVnziD3d1svhpm95twpD4W6ZJF0wWFe3gPgQcQrF13Z/KxF1P
C+HuAKeLPmfHpj30mXTfrCCDDzaZiTckWLnh8Hzyrifjibw381Qpo4JnQZ6lMtbr
5UgON18GBj50YD/wUk22A0DeXITVdPR8p4UJglmNTVJK4z2jfwW3tzSvRJg7Rds5
X+E2nTE+UPubXE558T1Zd/JHleQp4R+MbeVsV/2WVYLJqnRRYlfaM355GkfHrkoS
dohD3oFwgzCBbv15KJBL0UheVQQtssg9wMW4/Mp6UuGGhZAvwZWcdlp9wSGXExMg
5TlCoKss07uU2XN/wia7Fy0WHx4kdD6WsLbP0grpb5v+/iku2Yc1arPNbacVBF4B
FidDn/BONZ18a3wrWJ0dbEb7oBjpwUrQkEYXRJyMA8sy/YxLbvM/jVNj0KF3BXpN
LG3Fua5t3PNVAZ4X9FwrwdQy4GsC3T/sXPE0bSjVouanStsBq7SGUi0Lb1bc3p8N
sPvvWgT0QFb1pYBG7Vm28eiarjptmn6uVytpabKonuas/IBgo08QEAmwd+CeRbWx
9K5sGOQ7opr6LQAFSrofLIAhbCMA3CYXjNylGDrBZqL8IBIPEJTZ6ZlHkp14mE1I
/ACWRh/yqKMfQr5YQe4wkAy75gwgy4v1qR8k4ZX4VLff53G7l4ELILFytGuqPoro
qSBudMG1bfNVmFaSplMlJUoKYHCWmucf2FBJAbXNtfZjlwKnyfjZ50Q4hzpB4cEE
xw4hQGeu6sTPVWlzaK3mP5duxQhYWKEPCmU9uFgDm+q0SgH/l9eHoYBCc7HiMaYK
92RMByRhIaZE9jf8DAV8W+uQ9SnE+ngJlYFzLHA5qarTI088d7X6PSkUGqJlphan
jBDVmS1jt26W17bB9/QdrRhVpTbPAGoLM3bmrMzxZVPimVYKa/BVvMHj3k1IC0RR
XL1TwGJOeSz3+Mg8ybplUc2kTdZs7vIKoMoOL3eaUfqs9/gxt3PO7rVOz2mPcpZF
n/2omt559KfhVDAKSa6knSbGY08nrOeM7Cp00f1IUmG5MuLserGBycqc2jQstVgR
cHJRNilKvJsrxwJLUe3AK/EoS76HDKd2xz+B1+pu0jVBs5vtfhTq0dtlLEYLYlN1
k+tMG9bMJHNYchm1tVV02Z/U5GINduu6S1D5M6wIbcG+nE4JAIlRue7ecQczcRIw
Lx3lpOknADo+stBjtkrGEJ84lIxRTkjEiXPnChwDfRP8Svo3uGESGQVcWkHz1Ujm
le+YTaVkA6+9E/is0JD0oVE4gc5aL8jdMbbobAo+LutUkfbSlvSKwe/rNz+VCz8Z
51FeB/5Gw0kTM3fTm52kqkSwkcAiqJ4a8PqAhT1TKmwOtRGHk3eDzFMvXpRuT6Ua
qBVqYn+SZT1IuDrkpHqhmZ7OqF97uUWBh3bHhH6t1j9qItwWQVTZwaciZpsDGaJR
QklwQFGmuAP9F3DnkjBHKVxT7VsOz1JJrpANU94u6jx38UKgz7w2dyAzgscO8vB6
EIiu0HPmJm3TwVbGjtKvqWp84kK3dd4i4ZUMK/+6HpmAdymNj/iasOSKa9H2Vn9w
/HFy2lWeZrukIJF23DDBa9HHx2Xsp3PBMPdEVBW27veKOpEDydImltDVLqCET4qf
1QahY0wkLM+r1F/RhAVvS9iewQvpBvDn91+bYiZimXmHtztV0FyrCegCIW7p9SFZ
qpIW+AeCHbZVqJUrvU39IrImSzItxPgPh3fdqIPc2c3Citx85iGNPsabstoEQwEh
F3FIeyjZBfZ3MDfCDrkG917nh57sV1lN3j8i4QuT2KstNdqfNOPELIHZXaaCLTQm
Bn2D5PIKOUGRhbUhCel1cJxn2nCm6TpnDuMwZ+2dx8+Wo5PsfyBBNlcwH1zzd+RG
JKVd+40vVnp8hDGh8ZQ/zgZGuOEmF8A48aBxcZYIR3yHT4qaMM6TXVuMgJ8MQ8KO
ZIpLQu7f/UXSE6vNDItdZYI8fXuanoVuRMmUhh+UZgKE98NAF27B1wknZrIDv6IF
gaObT26rfXDe+kLYhQz0yDq35BckcsIdVQPaudg4lu5x/LPRDnRwSVZMqo9Ll2KL
x/F3zV2cP05NBcqSrh93DNnKuqCjYMP9H+ugPGQ3MW9vbiRZafXj6UY4VybJoSVZ
jYw085pL2f5Qy/IJbLhOCFGody5hG9uwKxao5D2gYaH65JTw4xFwsJ1fpXdoeWI6
UbIUNej/Awxb8s/AeeYsYLAMSanyNtnSZEH6Vojrtn9TwlDsuLcYH+DgYLJRH1Gy
kaN/OPDX5IB/mRq7lgaHcLsNpr/Oitwv/8a8vc2T7PT6kxW/XAUd3svcYoHfeDbl
vvbUS/MOqi1kdOoM19vrwM0j/1RcrtkKSbJfrmKV7elvmlaWf5o7UZdnIhw8XwuD
IkvLgoebuHMVjerv78AQrvLEC2xmMPlZr9O4cHHua7LnxDQSUFA1C5QIws3DV9AI
jEmogmegfEmhjDfq3z6Gb3AXo4TbEaiC/rH2iUAbj7zAYhCrC6gCNRuZrzAmcwTh
3cugidu5xGmT5IyxE5ZTk6MVh80X6uXeE5TlhOrXyH8FqowVQPHqkwLPaOmjlsW4
jL3bLb35ubU4jPxVLcTiEafAyIlTypshpPwERyGFlPrCdQHUkGqvzHd/vqQQY0pP
+hCCLAu1lLDFYtVOcWxSkfbIt9EXWx6ya7kk9Mnc+ysbb1q6s94I0qSGH8kJd75v
9wuCGwIIq9vRTvTsPGzqYetVuzQefeTP+KBMVij2cpBla4SDR0068e18xEowbBHx
ccXPpIeLaJ3ri11qHfAMukx7/AIsw2b3qByhZ1j9c/Zxr4plwx3333Rycvj3oGkV
v1FtagXCdFOAjdRFVSt/PLoTWVTlz0UqyeUepQM2X4c2o870/f+NpYKoP6GPqPFj
JIB2uyMdfQL5c4CZqm7GXh26Aly1/hrvEz6FJvm/EqwsF1BI1nEzzDlV/qqMKgYh
qDif/3Q4TZYsS9UEYN1mEDTIonZxIFH5ovf5ORXiLDzWyEwy0yTgqgCS7gVPAO3V
n/lNlhIXDSAo2AAafLia2/egGrZP/w2mZTLaNtUvTVB32Pj5i496W2W9K1h18yXv
01jp5RW6sQFLwDF/zaGIJiqs2oiScN+ShKPYxZMeLBStbbGGYZ8YHRm5QfuUYSPL
mWuk/XN0u9ZFpogRH9JZ1WBj/03Pi2zzUVc3ofihMAD2k60YTd4wWZA5tT6zUWyr
ATePmKalozGie1qeVW24HFb3fHbAHrhHu/PxOxYJWP8Fur8MMfV2zueiPpU6NygM
ZqHOqnmZVdNR/jxJQ0sW6gPaZkZVQXE23ZZ1dmaq1c7OizMhjewrEyMogrk2xZ8k
fUBi5PXLyDfsD6vfvbOP7AZL3cjQCFco9FtsRuVTopxhkmfe+m0JNXAK1MUEGA9V
nO6sfRfxxe9SYShefzG1BL3xqvfVjxuIE82dUg0f0LSWW/z6fZdpuA22DTg73pVO
67HE8ZTbtEPSo5LifMM7/ETR0TzGkmzws9EEkjzlgpyGhLKcxoaEt0DGKELwl4GI
Lx52kYjcOxyvxbqIymA2iD0X34igwp62lTUMceUgF56acsun6VRmDn00T/aR7SfH
VtlL2taCxewKh4AXPpqD73AH7zQmQDIaUqhtw9WkkuTKNiPPaWuSXrJinMbcs/UU
gx7dXmK8zs4I1F8z9erRw8SxZKCQGgrxfZV+0VbmukVqA9TLks0Ky8tgQyHnTFRV
Y9HcjYMNAD0cym0UmDqduZLmJ8/WNxxMjKL/Qk292s3ekyG6fUSfBH8yCmzyR4D6
F030lcdw+a7FtL8IMvyuCSwMRZcdXZHwtu5vVRYTCNiZlZDyHG7lobEDTERTIXGt
hBAFSU6JQx/ZW259yNtygohjw0c0Yc5LURHsOTzDFIoR5HC4Dzqi8hBqwYD9imFD
NI/yIgaGCE4+2T9SNdvIHFNoi16Upzxmrq14T4UiBriLaYjc/Vz8kQ5633nXPsqA
svx75VacmcX7oxiVGOn+Mz/NyXy2jWIDV9QqM1ufqh1CqoplxIgixFs2OksRvAiq
rwAxkaHo6iAx4ShibLHcmspTwXIM0+0KYzhnbh6aNHlXwJIMlRKmgOFuyhjR32DJ
SEnNLQ/iG3lzU0Jk/I/Hasn9JIdDTQ4t8Luo+7VyzFw+Wms9l21F9qF8O/zGaHp9
nD0l2bxNMtkhMYf4JpEEh2gVw9SYCee3iVNS21LU9hKJc7+CQNmylYbk1+JSY3QE
I+mPX53dS7mPdl7UDfck5qbZRwnv4qm+bTr9Zm+wE8MOsBxbpwOiHTXeDRgieFHQ
/Mb//79bwlZrFV7pnCxrBkIot4f17ZhaTBUoETE0cuH9hFtmzJdcAvrIomuKL53j
NB2wE57rvvg1k5BD7ncepKIqg2uoBOCN8IaHtc3yZhX0dUB1Of1rEd/w9Ud6hcTg
0bmfl2tVJZHxLHMrACG2syArdhA4JD9q9yJiORPIcTYWQiQzrWY0DodMsHAbv5cH
XNN5QI2RoK5PAo+ODAtyIZaFHJmSh3L7NLV/o2LTEfhX7q0ISN+dVcEM3zSU7a39
Sf8KxHtyAov+YhNtidNvgiHd4T9Xl8TFl2WGVEKa5E5LVXPNINQ9QJ1cmWLCNBdg
HyQUL1bvwS5Tnsq32xHMyr/s0LeAmCTlLF3jFK8wv1o6XRKZufN7UMF/LljizR1U
HJEIy48XUAbikMyuuTGdgafpam3mFLhgx4c9uyEGdsIjPmTE1W+P1kDojAcjpu1y
ccSXUbC6XNaXdhdWQSjyz2Img4ErC72/JCYuwwTIrB4VdsYYgmGAP7SWKj81GPNV
Dp7HJlBbccOTFeJu/55UqwqEKhmjj2bqbtSHxHbBJGcQt7XnX83ZNkKIp1XUk4LY
VDkJmuqXa2+ph/U663hu36+/DbrGrdloO308lS6qcnasskIZb/9CyKKh0uXU3/Qv
TIFokoZUILweJL61IGCMxJOHJuXrlcDZPLLYmLlLZ1WiGDwK3J3pF+UKRYwUcmGR
AR0QDa4DFIn17rnmNQZ8ioEYvNsfWo3aPv4AEWajuJui8n9PMP/6IOzmrMKPhVFV
zzAeh2hnR0SaFdZP+r/G5s1RKDlVhu+c0kKEwt51jzJqVscaAcZlOOhhyTky2VKC
H4GEM+HXwKPLPNnwtaz60jKXsouGKJFNhAj8E7lQq7FYgu4Xfd3SOmNa49aaa0PQ
OGZhFcsPXGalFtFPJH4jstOAIRH2Fr8xoIvyk0BGRyQ62m28tJhrUyJ3dtZBnJxY
BFF9vwP8uPsZ6u/3aIgb8I1rm35mSv9heSpBNhAEJ75F8SUPdQ1J9vnCgj5j0guX
j+ovdL1iSQQjNNs5s9IUMXQXfGr0foqXO6WkWdtOMYkP1BsNT6G1ad7XpyBejj6D
K1X4ymPWMJi3MtmYFX3YJfaKwOUKp5EN9LxpyzQOi+lskj70wY1yXkczLlGjgvN0
Yg3SHjSOL9V+PIm5gVTTIKbRjrzuW/BBXnTD+CvYvoXZFMX3eW3xDIQA6Bd8FqeS
aajLaQu9xxg6W5jJgGZ6yBdGxJhxRLibLlho7FKNICybrAMNowBYYE0Wa7e6U969
Q73oS9dTUnLaNE3GCG42mEo6lgC/95CYiufW/gX3RJV1unyAwn/pvjn/4VG7KCQb
/r1AFLJhLEDqz6wcZmsu1TQJ+jGP0Qc5rQ6TQE+tL6tLJmkA7O/c3oMkxClASUAO
Y5Vf3jAJkKT7hPJpBiB5jbcRg4Z3fdYfgyciPbVrgNsU3P1Z2/559r+a0xVcDKFt
ILwGTjBwUkRRa5mig66fZ4JjwlS/djUVnxuVcz14Zir5F94GHf64DSKs/iDVNvUd
Vng1JpnF/oueTOQ9zPPv53Lp3le44kWIHTjgHHHzLyi9zTQlEmi7YBqHfjk3ZVnv
h0h/Mn8wArsLJf4UTEJRWdW5AEHRIVtb+SZDnX6N/QPotm1QVrKjeSMz36i+tpTA
4QzGgK4VwtFP49LOzffcFl6EO0touoZplVjnpEp/mwT9YGq60Nz7xLsEVZZdltxq
Z5Kb/9KHmejwuz/ApRANvkXlXhw6Qi/xkKZIW2Bdr2/q/+Jf2JJeJctsdYKgl5qx
9PvcHCe3MEcxNav6C7XSykGSEFV7T2ewOAMpiWFznoCVL2JHF/F02YOOPnVm4onY
a9YZFbxIuhSRXDDqqgKHvD9ri2cmXdm6V1S1vvNmDzahdw+4DMDpAt4AeuCYUfLV
nmZcU3lS84qHPKGiiQIyTecvO0JsBi2KacTPafNmQIQR1BmBWqC0Pv934+SKJjKM
+VhbAA9cfUl7CHM+iQQgPsEtsvWUdP4NVDTLXEtRVdgbK5SInEPschHrztSP43C0
WwaNXTC+gLqLMOEbfRomKVJshKhWZ/aND+dFkAAOgnBk6W+uvbgUpzF9+q3SwTwv
N0YNuhdBAcrDfdjHFdhYG2SUYlfAJOrf9GuVsCOVbxgpUQz5ImAb6fZ9JEX+WMWE
UyIXfyZSeAiOLFP+vYC1Vy4umVpIqPy+wG/CBHCuaJrUafEiO4W7z1W5XBZz6Eg0
ggPNRnIaFo8gxmjqoeqor5KH41bW7DIgkHBS900dA69cC0gcItV0bTDzmP72NV0R
qoSS7mfisyvZGicLLgD3Ghw+eTVHZb2XLmbczKL6o1nQAbfLIjYqDatqQ5Gv5HJ0
vcMgsXAE6EAFMJs68GWTB1VBg/M3yK7a5aCaGBOjn3pmCm0OPeMGnN8z9f8tQCEr
iD3XhxTIlLmS4J4yXXz4ktDJmtZCc8HB1gth/QNCxHCmEL2kNOPgOs392F2wvYBu
pUvfwxy72D9b1m1D4E/hohcyK0hS92/q38a+D2JOxzSwqyiAA37LBuiC1LoNRR+W
d4LYnCQdMNySBFqpLzl0cRBtcuPwx9bTf2MKyDQJzyGy5DNiqwUl0BxVgiX4n9cc
ObbXuU2RwNRJEx/rYWcsUW40rYvr1Dyn8cr6/jsQgiwrArKrFDLy4Yw2ozJBUadv
7KdDU9L/2fGxa/1ExcmDct9sVLv9DYDZrgJct+f4lj66lLTLMVIW6mBRakoILF3v
XBfGlYYgfs5EgAR4xu3KfC8TevFrwdDhoiNDgp1jSdcjtV2dD4w57JVwoZsAug2x
6mzfIuxMZMl8+5Xc9EC6pRxqnvy4djJdcsOKapQ7oOBZhMSEq6AQrCyGY4d14tli
waTFyvCPfQ2KTG1cnaXElXjHNXu1YaQ3ZD+hPzo/6rSTTwEy+R7P1Y6ljzs0Py2d
fnVg3KS3fSNJItX/DJkc/dGF3NrYCv5rr9i5cq5hncxgEHTXh4uhlJLzofuHgPuo
KvBz0npbWcwzcrXWvATWjZeMZ3vVLPZDBtB4fchAeevBESlf1BnrDccxnYFGTfz1
sgw2NkdYqJX6DWjTBPfUxXPiF932pZdrj8yIb7MZmV6cs0541AATKA/vo9kbzp5/
ZDfgkuZdA7YbBd+xxsXZVH1E3IhDOdr7fc4323DZ9KeraQvUJZCglD0ldwBwycoa
Q5XGWmmSUffUBom7FKh3Gmkfc26RsdZEDwBQ7qGwhQNFUj+ZCLfMgZ2vKt5CFaAM
dQkhc5AMgGE3jSjY75g5wDub/sKJB0mV8a4Kz+LnlBLNi52BOC1MUM4TbR/Gcp4Z
KJRWmsGi3PqXyMorKEaT4INqeBbIJYtXZ+5gUQpA5D2ILbLzUI8YRNyu+EAbWnxC
fUFRPQJHv+X2f8/n1lEvCbBqI47Vezj3Iwz/SaLDxRTDbhGec0qzFs+JtAMK0MAM
1SyCZbXt6FB2Sqy6zrnmZWKh2HoHysvRjzhDHzsO8rvu85jdE+YagZkg9JKgclvn
TGxUDKylu8ByHx+W5gbRT6VbA2YKruz8Qu1DmSS2x/wZSn7EGUQ6YN3sUZJEurbi
cMUKI2hwQzwfXkU0VmrDvYPOf/U1X8f4oJBmMCaXT0JaX8VhTmA5S/0oFeFztb/o
/NUfxisAyxNh60Btbs1Il2QnDE7/G2V1tM8RZTVCMCzmA99mKw9IBZj0fNEPkqqw
BBEPoTPyZs0rJ0jU3ULn8oKmXkLzSiacSO4e1oA3piqMRoTvKrssHyr6lsow4X0j
LqBSl7hanPeXA+5CMOTC0vt6koTRXkf1Y/QE7X+e55olfesMkRbKKPOgfV/ggW31
oevi3G1qL8sDnLoKauftAe0XZoZxEY+ikPoQ765E8Jp+tpYBxC6Tj80R9aNcSrHB
/aLjI3QkxFjTStaiTiKzJ/q0z1ye3pcU5KQmcySRpKpidN+sS/q71McMpPz7v5O/
RVOvPPkPJKOEByvpb/dtC7kQ0UhbTP4yPgmDKX1KVrnp6xo6rtSyYJdhjLxuuiLK
qI/0wvRZ7bl2v2xLNdt+gOoNttGBGYA2UC5nlHYC9NuzEspPhKKuf9JaeMQdTIqh
Hs976+Ksx6v41YXiEzSiguCTKMWte4D1nhmx/UPPFC1mSjB4LwrJsKm390Wry8iq
hzyh44vehNMUCQO6qKn0PVTjrF+B3kSwXAHZ6ul9GDXF0Tv508DK/Mez3J8UG+r8
fOLAdqDucB91xEOSSu0A5ggUQYgMSjTxXFcYR2p3IhGxEaGI1AyyYTZMhvZsENnj
fqWJtPEREybjyNV5EoySrLaUeLxyjzRKqri53lq1FOWoF/RZaOcpUKYjfOus7jb/
0pHjhMqNlMosYJBN3XWFH7wxSKPpbcdhpb8CSfXATrnp1XRlpdEMuGYHMoFTAHhD
RjtFtmmxB0R4EPrBi7qhrKt4CXEtMrWUIhw1TJgzuhRvGIEDnCT+Fep+OQf0E105
ObIDH08IoyePpez0kXmz4rF0hKuzxnjdRLOHJRTsUwSuKXcA89mopx779RDqoBA4
04VQl8eIC4Ci/asekJpoAxCieHBpV1YGGqyQOhQwj9lXF/WflezxmDXxnHTDcMAj
WtiI/GiWjcCOMOi7oUkQ47Q/v8AOwcNPi/BsVjY8ThPbJNoUs7s8gNtvJDLyUW/e
nS/VziEEIWqLBpPlv7vv0x+EU/UupH3cj5FrKDqsidbemwcYYT4SsGCGdoSrrdHi
Mg2jFf8IX8o4feSm7WFh1OMp17EQowmmiWY3p5PCpWWbIXR6OOY4guiIjSu1YCNu
x70+WjlI6hCPWOnbo2qNGYP7q7pk0lRoTRbskVGD2C+n3J8Kmb7iwwThDmvkza4/
Z70CZAVWTTzrPer56MY38VQh5vTRVwAe2DrUJ1pOF8RL6c/H53jA/s/tkv0jXlRF
6XnPxuKVS4rOHjnnqKDRdIDgiZTAye/MG8yW0am6t5Wx7ZN7Mh/IEJVFslk28RAd
8UwDUzQUQ2juG0A3t+yiNIIXbLY/BFTaVI7CN21wAYlfwyEMGbbtgI2dZVAPzbZX
6iSE/P1CjO9feebsZMIQeBeP+6cfk+FHhTv+AK++4agXCl+gMHcMZcvtDrS67Owt
jRySjGaZGdLd/JuTAkslHC0OdzXLjTKPyWiR6eOiD13WU9FRLHU3iAuVN2KfaV8f
blZOVqxHSas1GNPPFKAUWsn7yHFSa8N+OEqzOj+b13mlKWLcFEvu3QfmuqBTggrp
3NHfSvr/6o/tRiHn94j2DTHWCmjDWQBuG1qwXYS8v2es26DM2utYjzRQO/crflQv
W9RURSk+DewjTfJ7vBV8WLzQD4ao372jJel+JDm82l3/YkJa9DGMYAuR42Mh1aGr
yb8LwhlcrT+Jmk8tPb9kk58AD69k3ebZMcrvZj04Mq0IEiat3i4SWAH92NOfoAc0
2ufSNaKk4NqBEahga1oz0IlX4nmtyZXKnRJ5/TOpqvkHsNdlEXwaZ99DJE5siluV
mvwYm/xR1zOX9AxuuCzF86Bl+Is8wHGt44+EFyLXVXgkOQwBIO8Ey0S+pOZaaWBx
qN2/B9tFYV7xsogG4FxH1tgigDDTu6uCWn2XPkftHDQDOca9t8fKlFpGqJXCS98G
4zd7zHG6xJgq0WO5hp2M1Cy0cJPjOyAK17T4YAMYaMdM9Dr/Sm7jBx4b8Sgm/Mbx
llxr5jNqrM9/5X4krvWdeQY9/D8al/x+O1DczJKi63KKfEo4GZplh7uSqDP3n55H
kpFWtvG97Sagu8pPby+RrotBwZfdCIdYKRuH/o5KgdNqOIFslo+XWjrdnGY872rK
fOs0nr5r7P4iX7AhlFf9Xj+vq6RPVg6CnYYBv3PspppUa15EGpEcb36UDACymwxF
0JlN5ptZyHPpjJABbpFg21kaI+5r5AARgI81Yo+kYrhGuJY7XHvN5KzK2hjRn5sW
JBqGmjtvYCcZGdzU3/YI3UBbtOWqlqfFnyEBTFCrzqmqhCNvugQHKHy3cWEN7U+Q
VfhpD5O0xTluKLT7kC2aAbu7pA9Sn+qyx6nQB5+GDiLj7Z5JaEw6ZdcUn8Iv/jsO
0+SF4NmGRgf4uFpfQPH68wII0XurRp+e2KQDPY83/uadLnJfIXtKMe00D7br7sJ8
fjjzg7a+PEsWObUAIfhbsrTfkOCEFfJsujQclJg/T4rSe97Anl/wXvwBqsNOW8S1
eX5YboVX/5qB2EXBFQf8rVrXnIhpe4gHiEELtgGll53aVNIFRJhllj+B0/JE/8g3
kRYLJFc79FssJDUn4O2WMkoavyQb2j06ftVCku47ImgTuxNNb2PsctNPlaJ2gtm3
SUOz5IqFwy1ShorYC5ILqkQaHgexcdbe+Om/rrY3ir4igSqCNbV9z+CZZEFKRiTf
mBfCfZFBS9s1bKgHBEvdXiovuGT3Dfa9hGdrn0RZ5GQ6sQoczbcHD+GsAAX5wiMK
N9QE07gH/ggJxEr0yuKyTREEX70or7c7hgMm7whJf73Bzozrc/2NGjZ6athghB1X
LzrFrOlVS5OWUcF7ebSM7wDdDHKVFU5Ym8ns56btPSMOf8hjoVoomB6SvQLvvd60
BZiODByxiqCK3NxMuFUa0g==
`protect END_PROTECTED

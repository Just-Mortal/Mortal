`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MS8aLTpePX1XXMngpsXYvf4DAIbVN/Ps2M6X8QhA+fE2WAm6QELEpX+y4oR6PYuV
E4xzEKSmf828q1/f6ib1J0+EyK2zxTiaQIZ9mSZogHoyENahoufLbCTS8n650Ksh
zS6C+JReCK774xBzauAzxFAAmKkaF+ZIUOok+C8Sfq+UC9HI1P9O7AEh+ibBqFlo
N7TO1C3lf2u21I51dT4Yx+cgcQNwDd7kspb+RiQAtae1KRDpUGkAOV/FDPx5jdLV
cQdKealUU4wPrilSp5hKe8Q0fKaxV6hBRdTpNy1Di/xfFl3Bg0pNuTlOdGWihJ6E
Gnxtx40TI3aX6D04r3yGoq73nuolHNKI+cURw3cWaXCreXmQPSq2RuQz4/wdwCeB
Y8S4ek2KUVjDiN+FzV65CvGK96XkAkcoUDUL68BgEYA=
`protect END_PROTECTED

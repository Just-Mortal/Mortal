`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
co4z1rxuWr4IjSJNuJe+paWrklO+slDDihxkTuyVGJJvOIE6K7YiEemjgO2VyE9Z
ECy+7VR4Y+0UC/y5DV/0u4pcgHglX0LhtmR5Z8DzArMMrMgplv2KeE0ErED/Hs1+
y5qBLx2haly/9AyR/ItQCB8DyGEXdd4RmbA8/WKCDidir2W/sOv81lHJ0sFnFo0b
agwriQ7tXaB7Vc5vTncJM9fZJPcSCM1UpRh4A77uNwJIayr2eN7t7RCaajZnwP30
COduZVjY4bT8F9NeiX/59v9AS2UeMNA8e6jcQyE5XluCe5yBLQabulHS1RE0r+/r
Gxg57zSQCeU9NKY4aw5z+ihn2q9BeE2+4izvJY8ZlqwX1g8F+jjcBaqJcTQsy0Nw
94p4hzDuqeyNBLH8cW0VuNIqlNQpHB+7lOV6iVtwvIBlErGdS9+qGUW6z1HMO2Xd
1WhLOQvzSPkokv6QRnxDDCnwePkdZIt/c/GNxqKHlTUxDPU3qKtZxDxPKS1edCKv
Is+FoPB0zrKwZNc+fOhX8THIz1tsRkyuB4TK89HYbLFhHfCI95bJLsPYQPoO2aON
MrXeM0xUUF1znv2oeKBOg7rYaJfLb1glRklbEu64rEW2tvvlHkOHDiCWZFx23Xoz
qTCwRRs9xD9Mk/ExEMxcDqseMcRz6mWlgINl2Huw6NoVSLPvy8WL0TFe+DNi+gre
o5E5Xm4eAenD2emq9ai6yvJWA1UP+2LNGm5UKRlp1iQNzFLllCB3jw5QqrqzbGlh
1Yf7tyJEzUq1SfOtWlYvp7bAKqgItxpNzCjp7QPWZ2u9Y924JyuAuhq65bxRFL9x
GCZd7xQ0K6hYBUDnQf2k9CYn6LJaVZ6NW/vlYSDJUUG8kpB9daOy0ItogPclfsPh
5OaOTFgr4x83WLT0SwNSewY4JCrcUsVJnkn5DMEhsgJpDR0W+3gQDxyhw5ovNlsX
5e1wfJ6PxYQaF57bSjSRKCKxuOwyjIjHb4CD4ith2ITRNtJ6d6WYSA+U0GFr9u/I
WQxkRDKrdm5Q0maRZBJL2jMNEjAsKXheIxI19q6KNdgPX59ZH1uqubW6PfE3RuuA
+Ar/6GgEFFGFyBq+wRqtZ7+kPT2VC3BKhMOLip9Es79tsQB0d8ej0RIqM/fGrO0y
SAMbFkNg39w1txOkBU3bipt5juqwVzmFkD4nBwAlkNbkdzMVIba6t6HOPj/ezf9R
iQhZam7O3n1+G8Y8aQO3SwVrd7DQoLyKrlSc+o1JcktMzDwP5X+QLqwnh/PtLPbx
knR/ARJ9SUfj2Ktyem3uoI4qHV+FasB0gSmg0rBP1Kr+6yZgI1dHYjqdwGaISyHs
ufoz2fc9ColEkZErw2maweJvslAQcG9H9OlIWUKWep+oRMv6koPHzgJVe+45IzGN
hA66NsQ/U+vlky0iLihpTPAGZRUcT1vCWTTHttgV3zaQQsqsIesYEzgyao2L++8j
jUk4+L2OWaHf7MXQiS1VNmjkNCDf7i33LXiXbF4dMpTqGXrTYufGPbFFC7cwoYxB
aig4EQZnO0iHozYx8SqE2VWJSTkxBiLP/vzxTBuZP4/JZ0leEBvS08EL29DMnPKh
Lup2brhlJGQxjNaKfUBFjezMVKtO3OwOQBjNJP2V0UbRfJ/H1E+CGuZrfYsUzqwl
qdoX8bhbMIy7IX3pb+e/YJRn0aZ5ElKfR8lbjAP+yGF2eJhaquGKK35DWuQw9z6M
08iWVgKjk/NOxAk3p/NqQ/3UoEmu+aAhh90fyBjAQH4asglkS5597SsE8LRtXWvt
LXdz9mrG1OJE/pxIYwwyl5whRQaEKSLJIR4J8PLBtj1MH+5qzm2HlFwY1rR5N4sC
Fmfl/iNRPcM+sXsK7p8KnwJ9NWHJcc6l5p7mWLeV6CzpSyAWlnNJmaBcXytCclLF
oR/roxLQm/e9EUHGJ6tBldX2POeV6/NRXIzeMMy+j5KkwSL/vH9mDZdxnrBmnDF1
cc+Z3wv8qaUwSzYdkUlttljq45uQbrVUcjNN9fsyvJufTi3uZnrtQLhHw0uHLyx+
2YICJmx1qj390PsWaFp5tvX2sMktAIfpDI59onyCY+v3yVbEcUd4+SVpeJoWWclg
DTt58z9gFeVOb99i09PUhk/vc1yLY6AuhHc0eZttFpbbIJnzuz667MY7A1VRREOP
pWOGc7nfG5CIDkgA9WD0DNKFP+HQ0AtbTJCfkwKtMvCfRDR7ktIPISRDToEKgDO9
Hg1jXMCuMVAhNqx2xwOyswQ5nFsd9mQkrVFfa74oEdMNEH3slCs3QK0IbmSIXizq
pJKcTphaZDY2LCHkIRbPK5hkTiTmLHeXJKk0KjpOIkUX642a/6Ei6eUYZ4uu8MTT
zDpO6lVIhJaQp9YGgeevpkfSDREDD42IQsT36AzxqNhJGvrrSLR0O3j8SVLP/3IJ
m0v9sEgDPG3Sza4edn3nk0YRf+S2tHfUEUjK+HpaD23QuJjL4c1NwyXFfs5Fk+Md
ux1kPOY7lylhUYaHtQGPNwwMMExoNzIQCEG0KeBBeQf3sGZBh6Oxk65+/piRqgMt
x8L3QrAfD0Bpn37bDJLn649cdwDf/wifjUCgndb3kNhxuo+DLC96tVHgzuSa7opD
ZGnVvXbdevjCjyGCD2vlzA+StV04KMoSOgmQdiQlbmKU+zpr4BYhHLzEUtZ4UeD7
txAbIrUqEXvUd9O+8H8czsJfRAkokkWn882vClU/CB/drXuWhuHq+x6AUiY3wUbU
pNHZuBjz0ziYUbn7406/ygC1AvYq+KdeSClhubw/bBhehlRvOLWcB1eDli3mVgeX
4ASG1iA5FPX9ciWACTYb2mBnjGJPQpKUjMuhQJ50E4dXyAtOZfeEioE/7aFi4Gnf
dyRAy3V1vLjAop3JgsJH7S57diE2K588MP9ulHDVYyEpSkxuhe2C92XEH3mC3PHG
2xZHLfNpPavaDabeVOOIZR7H8r27klPbpvN5mJrTUhyXptWfRecjl6m4n0XXu5G7
3IyDX6wZc6PIqvR8a1zjBJ9hCmDdkcIi3/X44PJb98r76npyzx1kTfrKzr0htAzx
ZMzIcvSvpVkFIdj8dRRsSQxEAjAGwg7XP1KlbAG5yC4qMsZf4RuElVk3fJGchEBu
hh8Xu2pZ/4kNW21Yz5j917/R8EjiN0Y43358W3nA+Yt9VQqCdZGBPeKs3vLidNMz
+qZHlQmiTXK0tuJfspNL3rK+HQi3eeTDedfl6h9ous3jx8QA0A9S96xSHFVLE+A9
Ca4+prJ78eRbQfGHyq9mtM+8mpCEeeRC/C5OJK81RNADqeGP2w/5Wsv8mPgyYW0p
FUmFBR48GueDunr5/TrH2k7A9jr31/PUkDuBebGk0yWrSnVxPXaZeQK5j7jZ5J+G
3DKkqNOL60S6TiQ7/70hnzyQRfJt3GosVZZQamOUMG9MxhnBel96A9z2I2kEgCCU
518+mMKIzEWjJhGFgCbsO30r+25M8/keHRehu6FWL5KL3YMdvMOsAr4dcvIuEBS0
XokQGBZ3aOWeO/XPm9WfHaAWTorYAcrcJyDVVV8hOzzcDVbuvs7JXLISS6zD1ka2
plt1UtyHQehjKhxn86U7KslZJf8ZxTzWTtSEI9I5atCoecjF0LNp9IWIAkQloNSr
9e+v3CqCkY0gcE1ugbnECOKWvG6I0SoOO5X300Cf9z601NS1mdQp5F7m0QcgjbcN
KUBiKhBXDPWNWV5EPxSSeaOXmUIboFx8DzK0go2RDT/m9mrb9CT9aqFYHi0tkiSe
Urz7D0D43rNhkVIjcSwUN1xENSyq/h4Zhx2/Tcz7mi74hW1BWd3/GPDS0xK2IcSU
R0UrXkzwKD3o8pjo7KF0HtnEzLvh2HlrRNxVHufvLj2hKWlKt2aAZryEx6o23N1b
3UymjSetTakxRffatCXmnYMYuoMX9Ys8vkZU5uZ+g10CrW8Xu5Edvkz75D0JXtid
Y+wchyUaRbajXXQMFdiQtpu2k+oALDleq/7KJHWc6jMVgG0kD07xYjdCq7y3NhMU
MtDKt55TtgdGuQfZtbezpqsjBj4ilpA6X64BjcerMB+UdWEq6hcVuQrVU9Oanz7z
BxbxklWC/ZTUprnyRdKUHgs68aU6FzRyqTNwyNRsy4w87iWjmDuREyomgBjZQ288
aijor7xLzukIE9SWkyHVNfdjqTT9F121FutIW+1YMWpXR5hY4HpBktG1NCCt+DRZ
8BaSVwX7rnrjfVvf1jPRLBLXYbD2T2gRigxpKD0PQ4nMCs+jhDyg+ypHFGuXCfem
DsM4fP2adVeA7nAdpLzBVohiqj7DRFIzgfCoGcMYHz4bm1NHeDo18Svdp50JrgIJ
DAzKheSza/UIhcJRsr2eoGkWgnnq/S0s/dC2ztAebvh1xrXQgOTKwuZTx0gQ1y91
ZBv/zK1bBVEDeLa8ADITYKMO9Re2ufiLAzV/He3en8erxib+vJWC/NrIQ770qGQT
o11HQoFnZYyc/mhEW6H/aD5fxdGKEcpsg4iANU4Dd4B+jgQQd6Wh4sSstk+30L6L
1VQpK5bkbXfOdkGOAa4yfcQxPmC4WhyVgBkAO2eM0zhu+SAVzVxCKTA1FChjkEv+
9+RpsWOknnH4aY8+m8gyzJJlzCJvKsC6e62u3VTcYDv0GoYBnR7hFJjHZ2jWgVXa
YSSTGu+nQG+xmfiRxtZPQUZE5z8SbK8bxow8jBWM78fNE6lhEAm9OQK6ksl/FYUY
mQizRbXnyJVrMlHRhG3uak3eoPhniTVAIVrA7TJGDDjTVQQiJMdYk8cgWzHOMuBY
5Gpv7A9/qQd5nPBoR4VOiwYPnAq6tqz2BIIOuYrGZ3ltvykr4IapX8CwKgGXywX3
0QTELgmbL85FkJWeNfGuVi/KVpe9qXr/bG84FmQS/fjN72jZ7pXQk2hr/AyCqclv
2MKj+faGcnoC2Cjp2AxUikzd+1G529YBcgfwI5ahKFSwdMwvnJIKzs5K10dEiGNt
Lg1o7aYxJjlb0Qger4jDMs7wAkoQ/+ygObHNYDaPD1+KWy+g+pg33FBwXzMALPkZ
IdFhGWjFOUPky46Yf6xiB+noTO/oypqO1Lbro5/61VgLb69TS7/9DszdBYdJtzv5
L3G29eA3H6HaG3VFnh5jLOwisFHPiDJBggZwctC17JqKMGmksOtAK6Scro1SMa2c
L3VzCc8BGIukc6mxcSV0VliGYy8s9wk2IYSya6t1KfoROTNnNmZJt5rUkdlze/7m
xFFvPD+Q3JWaE9MIbs0Vp0y+j6j9wg7zeBCpWSvZpQfrJ+mgoSs3xr0u/HNTu5wx
DZ3G9QmBdEi2YmmA2E6u2xO2Pr1E4cP9pJ03f7P0DcqgCG0EeqKojxshbH4xZ9+/
Jz6aGmLw6fsyCKMIN8H0K1uIeoMcecdOHxqa9lOtf+oJTRS7KEdaHtilxaAHLJHz
VR1lIP2uhXeReOMHxI+cp9wkW+oSqtUOD+arDhW6llEqDIkNsDlxWT1H84fA0Pmk
xV29KWhR5dCw5mO4swZ7CMoCcaQjSu5HB3pZt5seF9WXm7t1/Pg2IKk6V9IMHM3u
n6Q9c2JdT+9767R233zFeE2ev9TtbUfFECT3hfC7u9qftUV6aIsVJeJ/Y/iEmohN
HxpwSRaCMcKE0IbZssEvjXrCWwdTBqoO54mnt0XzyNkQ7kF4eGAKuOya6LUFlHRj
Wiw228uBvFz690ObdJYfHyONsPgKLwY1x/k+F26OX0RDCpoE7fiszqPaaZY0pCB8
CwzvUAPVqshvhSpU+cVTbiENc50Rn6tTnNCSM6gOm881Amd8nCdlJq+65cYnmMp9
MXgNr2FzpkXxVZUOJZRWgmOAD8HBhQtcrxgky+Tk/r+hYDy6mjlwyAQ45wsrvPgD
1TftCcUNm+adla6PfUrzFOCVgWs54urg3vKf6qzvqEB8qDL32u9tiuWbwQUkHeeK
cD6wxvv5I0PsMdeXOVpdYD8WDVoEIfjceB/a4Qumv4S/5XQ4xOg2gXGl7OBVs+4t
Yh7zbOOMFXoQ5/S33bzR5ZhHHtB0wQ0uzMufqayWc+h3os4DUW+PzWpouhxJxr4h
Zt+MJChPwyk/jjw4XjcWqy/y2E3kCXkkk4kRRynitjKKWAcPBsf0Pyrei1zsrtlF
oe3ut21yj97ItagJBuvsaaaVQMWFQs7fEeEKofTmsYmocB7uP9G+XaPvFwRqoEtx
XMdxO5b8zB+leXGIS3Y22FukEjQ8bGFi3miOL4ftt0TM92FbjGc/lYplP3fwpuWx
1qRoAmwlHmkk8fRW1xjBrT7m6EtB18JYhQxVTIGm57xKizhZpKA4OCbA0IGf9GaO
MZWrbg4Pei3xP7EStyC9y2tvxxxeFR/4gCdV2iDhyxmOiqwX9UGUTR2xnALvnaAP
zEom3WLvaYWJjC1RRr6i68YBTsUOBJyyhkQZitpWB2ZFLghpdabe0K97sNR4heSe
iiWnIfJLGEP6/6NFnea5bhVfOoJXLunMDEIFMLBBD7LFBaawZrxXRgXT5oA24GfS
HA2xDAp9dysFqsdkSAbUSgiKFnlOx510LI5nLcY5tjWhmAWniRGMdsTyCFL6w4pF
Xix3jX5YL8MbvOqeUA7dPnoOtCezjxQwkdNDuH7RB+vdG5bSFMwrjiagBvmNM05j
cSisx/+5S1JNgyNGyugqRbNcMcgN0amW8hX0FkYGyJeHeyTaewaEIBrvCSPHCOHi
vLGMSRrM5R7Pt4cY4KZknu8zZVrjNy9TCY5iaKSD13qGoO5u6raRDNt1r1/ZPDxb
JrukpHzWC2yxwritbJJxIMUvR4tq6XjELO8e4WAxDbUZu/jJYtasM0VKul9/fJpZ
0DMbGJkHtq6MVykkHY4nZ2qeWwwsn2S0eSwy+VOPw4c2CgkZT1n7sb2SLjxSOYHk
4eupccGJ1L3n4YiWp2/+rPdv4g9lqHRf07gzTgN/UOXtcPpzIu/AosZ8bguvdBRv
/a3zHtEE6iWpUfXU/vsO6NPgFqxaI7pmTdbpdRLLT6HsS0qLIMSWbSSDQmn/ukyj
Ru2rOW0kD//FyqjEfchdDovcizUxDjPkKLpMqnEzwqDFJkkPt3u57AgyNGC94tCT
sDF01F73FCfzU9SOOq9tk2pXwJ635pIMgmP47GHul4NXj2y2RDlMmygv61zUS7p9
yLK9QxXFYLFPIEvMpsaIywKY+iQle3fI+Wk9UdJs5zfDBJnHF3rxTIBxue9LFqEE
M1IEnI3D5c4aQbaTlVs06t1tPtOhMxfBih8ipaGKi66Qk/cssUO7MUn8Upx3zwWo
l5ynP6AVahZVEhKKY74Z5YXObklzFsSaRU9m9nSGJH/736Sl1wJDceM1XUgepp3E
eEuyJbUrx/fzGI+3tMv/ylyHinlqYsZuAPi5pPPvoywhSDvL6xWF/prGPeY9yPtl
s7oE0Buyt125lJuM5GvyZIOf0WSySN9xmUmF5F/cZvHUdAELVhQ0+nVYKGHRE0IV
Y/QL3xoSFiLs9Ar5JUVOAC/MwP6F5lOOdO1O8llXary35Om1g6a29jijCF/cnBSr
WPXjw42FHzXvV/9xbxbB6ZhEcO5rilFfgK1P6sUQiDXSetzRknbesefmMA7/lHiU
U/dNVEblBdIWvUMM/SYEkNU87MVjpTRnZDgaFV3JOG3t0kHZsZdceixKud/yA2Df
JD5hvqWtD9SBYewnQlWP2zXHy8vvdezUpJfQn3f92hl8Ghn3Z8TXmRJYNmkUuueh
KvzY5R1CIoLLpP2y7nWFNLOQsp7+GMQSzjDAKr2upFg2GXfAwUXi3wuut//3EyyL
5+Oc5S1vjaPte7rnY7ceoc2DM/O9ZyfrOmdwbIY8NZIr1sC6D/b17rL2VqsInPuO
D21fDYaLpFsasdFBD5sZV8sPGwYsk7+EfiktNtpwssSNjrVxC8jvGzO8icfIIiue
H9NfcbM1naCwo2GHgFXu7tkmeZSFuNLDU0fIiCiIxxH96vmJPgk52XzXzjRyVk/R
bnycNln5CVsoHU8JF3i6gyTUL3Y9Pduxejai88bd6kPLlkYxBAQVDu2boo+ocJBG
0ethNquZNJE9VylUqcF6KDEA8xJo2EkS/eNpkVqu4+3vtGqTs2dLR9tR830QMCs3
VX3cRKimTzWKHbMvg8vctO0Pds79zW95YPa7QYzFhLZxrXTB+W3NHBixrButf6Ly
eLh6E1dccmH5exNana6Ewh3BKyw6uVNFbGyNs9PCdA8dTaBs0RNs+tZLe3xLweBp
D5wNYWtxSFopGToT1yQGdL5GhHR0EfXfwO2SUWh/hazTuuqIYdf3/7SIOlOHczoT
nPZbFVLR2gPqu92prk9MBqUa7jAiGtQPvJRhzY4DqOu4Yva7JlLv7Q1bt3I/LJ/0
DYnCTfbbtyX3y1Jow6gVVTHVkOeIXJTL9ia4IbYhLDCHaopSSbXDHi6yVCekQY+3
AEi77qfFfx0QqkHuEEJN890upoEMoiIwh4FrPcuHYY4tOsRfzvGh/90fA2gfhoIZ
eDN/qiwnQQ5OncK/r0wf60y9QfSDgpUy/H0TrjMetVJD/Y+NYgmeHr5AKcOLKqEa
6ZJF4dKVVqkAEzL1j/RYEnFRk9PAA45jYzxt2D8w5w134UYQ0bp2q+qGrRyZsmRm
Fu352Ce+pRBMnSwvIx0LdKHVQd6mN8KbouHRcRAwk4Oy3AkhE/t/yERytn8U7XdZ
Nz+Rbi3w8u2FRrQG3SBg+ykANCnJmK9YhcmgW33ijyQ7ry0ZyFggqj7zRYlCsEgo
linPz8jP9dsU3EsQ21A57BbaA9+8n6Z8uCLvoYuOpfNgU6ou78zMYMAXyk0Sggrb
YgthZw8VGoi9EdeLVdAo8vn0DCIQWe3aSC1MGJeS+CvyVW3u+rpHz9/eYqA7aTi6
R/1iMnxY+GSnzcazks+BjHUgiDZVAiDrBuNVuwouepEfccFqEW1Dm5uZ8uM6a5Eh
SpeKjpqgzFMvJyU/qbkiTUIxXCkv8/30+Gbpw4oCmLm82uTjHEdzQYPwAqKLr7Mi
L+1ykeEbuvEM2gVarpgXGukt8lBBxy+cQKDrznJR5r+IFf+0AF+MuDLV7XzrTWMJ
61r7xCwlJZOahOFRCjylOqJdjqujT4MV+Ro4cVjjlZSg9XXQU4pfUz2pIch7Uagl
bGfMaYAKm5iIPlvwuf4hax+8u/8GpEKe4F01AqAFL8Z6TqcK+mLVfyOfEbbCWy9k
OeFDMcKZLO14rlTbaUqpQKKuBHXtPBWA/8nwI7Q1KuPT8eBqiwcnNFV794LwceAv
9uCP6j5mSdgbNaCk3ezlrSChMXmOicsAjJBu4Gd9GQgIyiZ9sBoHxk0zvcRw224V
cIwCH20PLmOSNP0sCR/hBfokejgDhAnjiGzyZCKZB0CEoUYv72xhVCH9gUmJV69f
xDHtO4udWPSsACaz/zyXF7tLFwpelS+x3oQCWOOYChnmPURxCxw2ZGChyDLLR7gj
+sf1v+i45qYAXBzqGGhoUbqvMQeNAfjyRok3GcFte3KtEUE5c71X/XN0Lz64wjvB
kmCYFvSCBpnWAGnWAXCZXz6uncFWSBx5n/EQlVsV4msjjLcfyEro0nTylCRDxRBJ
ufFXtLJPA6OtUI0Mzk1ax+qDKyUQrEkJslI/5vgFhrrhg4slwU2KIGX6hdUABOvY
8zPZAnUMADM1HV2L8re2td5WNgjtI288T9qkXNGlHbTfaAQVATIetczvJTVix2ZD
GBgjA4RrbFVxb7p5+02YSthITSD0F4KEQ3qm0Hxizci+bTdR0Z+GDxYfu/Q9X+sN
hf9vZATS9PStj8NpJR23GYCUP0MK6Z4wnPzju0tXY+F8x8Z5z6321l1Z2rjic/rF
rYBp7tD8cyvXLsvGQZLmhSSsStS8BQXU14+pX/QdG7x1Ld1H+f0azJ+kh3UkjQpj
ownBYn/we0ZDLbj4tug8w2qfAXAc3EKdeRVVt/wr1F354dle3NIELiYPJgUtedVj
ta3qdmXQ6XCTs1smY6FyE/7eCIob2S23g7sGIlaYeF4cULK+B6FZ3xdQat8Kg+0d
ihy896tdIUck7WQodoh+zmKamKFCqvd/SWDU05kt6MrBCVxKCWu5MmTjMu5cu95w
eodaP3niDU9y/qXDQVU0ZSBYiRjonJFMKRCeJHCgtgR1L/00+JjnTmh/ntkrJCbn
OvCakih0USNzmwBadhvcdQZjgFqrnAhDsSuLaFf6DpuyRBorRppjKGccohd4MQSI
xF8BjEklfbWeNiM6HzsUN5CwbtuBlKQJkUiIXg8Jy3xvN1yAAKeLQXQ4Cm6wKweD
7YndJNDjdbTbBrJfE9DC2QTMFpy0+Thg3VBp0iUObQHImh5JClEi2MX02vPssOAs
Z5MA4XyLXUpfPW0a2awE/rmFnUfdXbXPsr6ycVdw7B2LQAwwdwugEbevIzvhkNU9
NwFRF7ez3oYf6xmdZi5cHmYb5EHtys+5NQKR91yOjrEfsMMoV5t/wy5Bld+TuAw2
qaQ7E43fD6HJ35t48/oEGg==
`protect END_PROTECTED

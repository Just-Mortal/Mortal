`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oECjIGPl9d9bAMpxCa8vakpdhuhOuApA61PiIRzA0L2DXVNlri/UeEi3PofGIpYl
sbA4wsbbTvfd/aG1QDfSIxDdBn33qyynBC73WkWkM+nSwPZfkJ2CzOUJV0HQloFV
6Yx5yQtRi3ZNMUCHysv9uvActJXkFCS86dMujk9dA/V6XOFV/3NTtgpN0N2YSHoF
7z19uKvSi0m43kUiTq3Vn/5jUcxyRuciePkgqe0+vNYmqFnusvG1WE6ODma366Cz
OW66GGsQjbqjoTx806Jyfr9L5KXbFZs4ji12FZhriZCcpNh8zJW7ACBG3wsQr/dM
7FYOP1OT+IC4jrmP755dIg+CmLhgoqJoDEzi1OSZXkqImGEMP5XKFfL3YbT45j2I
in0sefgu0CnnwngMZuqnuDpgDqbJ2NjefUgZ/R22wZnQW9dfi89C/q98hR4Vd5d/
YxJcph/zEj03QtBOOsSLBQS2NsSO0OqaJpvY7Ut+SX0dF9bpMfD+y5B51kaT7DOV
RYTtepBLdN2wHMa3HLkw7XrnFXcILxqm3kCI80CFT6+munzNlhCaDXUe6iWU4/Sl
JB+EialCZtW8eHlnoXs/edZRsHRixKfNviRQTQMlLGOSHjbieTKE/N6YWenqZQZA
g3deo7s/sPhVEboncOVhqCHgwFplNSmfvMeQjWPcxuVGx37n8hL+HvUGPRjoJEYC
GiiqBGbM7OofAL0dwyrP7ps3YHpgK/z2CNH1NTwHquB01Hwx4jYLudWIaDvcA091
PXOrzRzRRsww924skjzQX31Pm6503aF5rW7ZDDOrk0Grgift25OIRSkJbNfW0ySK
fL2aMUYoNoZpy5pMzNqhbK2d8Gg7G3tutQhJQhlUG7LAsAuAcmsqs8ss6RPKrtuA
HbAr21K1sTAdH+juySbiz/50iLpbe5Ode4+l/8dfaOkBqZLBOc2/+dQZ4G3X17dO
sfBmF47oC3zOf08yAhe0mUXp2ZIoGX2XlQKBsWxbjL6qdDAJl/Uuv4I8kFJmhv2U
bziBqD4iVO6l/CYJGEfD++NPobBvZpWBx/LjxAOgWuhXN4SWsbHVTPESXGq/VvJQ
4AFO8hDV9Awz+kTerKHutIZKPUwbEk2bzAG3dOuYf2cy7nLpNceUvfeI7uu0ouod
g3L+XPTj1vK5fKttkt/vRWoL/cVvsc4qLbo+uOxweue4+VGjG4HomwxR6zd4F6lC
QVUBY7TnJ8mZ6BxogrhtGCIrDImuOrx9+k/hgJ7aBd5lkV93GignJl/wT3HLzNK1
hEvMGdtme2qQRyRqTmOhPWj1kF5wUy24ALfXK6081qaMhhWnCJjzpgzK+AHd4K9N
DQlhgF1mam5hmmzwKEk9oSwmIs4any/+LoXYBDKn0+kbblJ2oRD/hxbktFGCJtl6
WeCoYwnfYYRlSIeBilQVuiMoXtNLuPUxDyY4TDJV5V4oBasX5MgPE9rfLQTO6z8v
EFmEqVssxvJm8a2ht83y2NA7TXpSKWtWs6GXCKdYwt/0+r61EmsoAyFwJUWu48pP
MSd+2C5hjvzCCu6mKduquU5/DBP5nJrlRPsNwnG7amaeDrT3PLs/Gti9X8Y4NYwz
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0dXTEolfrxMmtPaM740DtNk2xPCmaNfPGJxZYD8wT7ybcKZ7OmPQqtP0LiNjw2dF
r9aRCCH3Qw+hcwKlqlzpZbYbuVU6peXO00YzXgSjMRJaxQwrOlxTbRbZqB6F05SC
7nDnyqlfnLHTXqHolBP4Ua1/F+UXWYmaKEDxDn47vDwpqLepvU4k9AZ7FhRPTp5j
DfJ73qXNZU8SKse0tj3NK0/oL/viYT7Ej8RSRnHv4TX7AxefpFkJw0fOQQ1iMo9n
dsBoWaMv064IJLRIuazsDylSRt4Rt0PvQ+6Jlm1iNwYJjRAWA2YDHCiTPyn6oZXm
NZlN2H+j6I1aBhcQg6ROwtVENmcoLI9KoCtD95Kd7OFFhpMZ0newt4bZMsYxlKAr
zLt5pv5ga+7TwHyekRrGghipvlTJnFYpQ0mv9aT7iVaj6GKEA04N5Y5eJYWKU5y6
gNQo7/DVwisgs8kODhs7lJLPB2pZGR0n6KEkkrnq65NnAqNK0ryomqBbkX/bGBwi
8Yr7bPpTvOnMJIo6XqUvk1nappoiN2dxBML2HiF5feJWRNZGjOmmQRmWnOIYn8Mc
eF7Tn1lgqZ5CeZLQwbZ+BsC1S2naHsOmxZTtbKlongyfdzjFnBg1i10qw3xi/yQC
X76P9qkwliJk2Ph5N6jibR4U0ZnYwkHavu0HjNG9O0DWD1pRdmQnS4IDnliofpwU
j5qJ3otF+MOeXVUmwXo6hiBMSdNQq+EvQy4q4dMTWYkCWnmnn8zOpVm7Yzq1y8ut
AtxQ12DbYnONC1BqeQ8wpor9KwKDWCusqCiPCAk5CWcgSFI9ZQ46nDyc6lh0NHei
uRtyfIb7cY9wNU1wHXEIk/6m5nnwpnWQ3j2ugHqUosuSuPVA4JdHguDx4CDJl/Mk
CNHEp0XFSSPDWyj4uo/JEjTGPVEWtLLvmxOyf+R6ZmS+K4FQ5VACoVdQ+tG6kMVQ
gkRG2zKCi71djWRknQCq1j7I7Cke8Lm/FmNaw2kBbUudyLnyc8+AeB5wyVBdZOxD
b3DF0QmjidNV4e6yPIgw1BxYg4tEHwGJsw3T74gtMWQkaNPhn271LhIu4wQh1oOX
keUIxUs71i18bp+35gImT4ssT3tZOQnN5W59EA0bpq/9LD02IwzGFHwwELtPUURC
8DX1+/LkFyS9yJ6L0P8xineDSZk5YamIomwt/EcZpLKe/FS1mjQcE9nxoROYdO2i
zr26KeHEg3m7mIWOjIGCyKi94WEAcUvuLQcwvgF40+x042Vmk69zDBQLfsa4RYPx
ext8ir6xjF6PsQ1McK06Cka7FjkQlwSIGmrEijjlV56OglV0b3eVOY27J+0DcaB6
+eO8r1yiVkG8dQcbGpUG7QnfOqJFvObZb4PBZen+ir34rBVTeOsgHzWsGYs9UUVP
P5T/HYND8ok+6qEA0c6rID7WpO6TQe2oMLVvsEa92RPpEMWxV7qW4Bbnnn1wwXCd
e4AyMeKvA0iObG+t0azJHNVFTIOSYJ0FUrVmBl/OvJepcEdJo8Rbv2qEQN9GC36g
xlO22N6aT4QZOH0/TRczAAWX2SSeaRC1b1P8lTNh0RmUL67KYnyRDIC1xJiPWZQt
vUwVvcvdlPnDiTl9wDKErVsJZKpD7zmYiAammNTui2oxoCKY3Kv2XA3h6hzc7Ljh
voFPIsX6Q/jIGfI3XLPNcWs7Puo88R1tIOIshgw3aor+rz3x9w4AnYIiTJ93r1MS
FTXDRK3whXoN0sPepKJqv3Y+1Gxi1ONHLyCuRaIrzJtUmSqXBrRtIIkTfy9RyucT
fAKCY55jE3p95Q3+wXbgSAheIgPla3ZEsEskT4HRLNcGvl2zT3jUtg0CERsrP6l0
9fXRZlet5xkmPLcb4RG8PGW45pZZZEX52NuHPYU1zv7d7cMjulEHc/8/VM6s5VZS
52zf90SIXwdMIR7Vn2md8jfV1rkbI2M5vPLAJuztE+XEaWhEU9GcqTZIRbGDEHst
mxVGXhNcfy8/KmqWPuwfvDSJjM73tGj6MKDNNQ4FzX1TmHD+qrZ0P7jH32Z1P4d9
v2QuUzKXstYTseH+3v4QL/ABzAHHh6WiMA8zESw2jkPZV2ztodqUweLLyXHQUPx6
CVmeN3En0X9Pa1tAL+95AA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bLpU/dnUzuauapvsaDLtro26van5h+taXG0z58maLUJ1Kc8CJMwDJ9TaSoywM/Bb
2t1ronVNg4ht9/ChjKSkqaCAQzr9SGVaWHGqT/6apsi0QkT6ZzLaAVmTcFr5Tkw0
7nlQwuZOSw6EoBnX/Av6EezuD7GmfI9CmoZKwGeM1Ewj9DG4uYwQxnqDVNirHAS/
u5srGnzUhOP/2GZz2GAOkZphbJDeWCKZnCJzwyUNw3CWNm7vzQPvxA8kB2YanMkd
gbpnP31GYRzDBvuimXy2IGHDni50QkVUKM+Hh8ZUp5x8HjNatQd1DQDPlAGeWa5y
370Qg0614V6NRiM/74u2CJuFOjlJ+bJM6i3FO+9vBUEkVexS1FprPcohuRtfLQe1
gkG8xOo9g3DVefYLJiUTG8BuFSMadZQa1r+9BgGUgNjvLs9jNmIi90BtiPlK79qn
4vKtLQKIG5mnAN9QakQv682/8UrQAQp76gicH1laARCVRDcYbnAavJeKMoh5RuxU
6AGqDPLddXLeLZbivnWDuugOi9QoTUoVEprIP02ZYByYFUXdGsorYh5uc2zKlRcf
VIFNDFDJYpzwERqoKzW8sNnLArl/7X+6ekPp27Ks1pBk8mYXFcE6YFFqAi74y0Mn
ZkKlvOXwizGHz4TKkJLEUyXk/cw3p+uD6IXQpznFc80yJa+GmUxt4didIfE4y90D
CuM1XRlf2lDBHfvMRW30Iw73hN7ShOC3icMXt/K4Mz1ffwIOB5W4ia2UmqHvKNP9
idaxRld1wRsxzOoJQXctdD+HLvwkl0LMWHCShQSHUFcmLMOmRB/BWuUoPI6QE909
e0yBO6Gy0FfZRJVhukrP7xFMxRVs4/u7KJFfHFNriZjpVglBVaWaxeVglm7aOZbz
jzLb0Naj4eOX+p2F2GJ72t6AuiM7uFaJqhiJ0o73aMs8ug0Cyoj8EjdyZEp4SAAQ
JeJHTfz4/60fBGTJI0qvZTaEA7kTxif16YpRsocGPWOJGsv4gOm4bpJKnjgUrLC8
+EpBupAsFdQBrM6rf4euHfskkHlS/vbUgmjm0zZo4nPEkf+NS7PbM/TyMNYILo++
o5tln3cYi6u87b+R6ogRtNJUh2v+U7P5NncfOLELK5ZlNPKCt2A8JrqII5y5Zbrt
ehSA3WZUq1TtYP24ABoaZM9a8h0HdIF/RE3GisoY2UprFjF877g/SdkGRd1nPAtp
S4vhy3tgSLdJWudIUEeyLeoi5t1s5MVDWQELPDGDPI+M/yZme9QF9goA1+SD5thn
oQp3QsmM0JA5fRFFfqFhIaud4KOYPjZG1OvaLiyrpEgnrXycyoTQkzdlS9rwmvLs
FQeL0uTdOA706pXsBrI9ngKd+YQRyOckkDq9OZg3EzXJKM9UuPhjdwSr3jo2ZkOI
VfH4NKLOzKEPtOFr/P79Nzf3QcRlPbDlpMJTdCzloNtkPE8oASAlrw9cTFyjlMlx
U7UVy2Nc7v+uvvpvB6+3hAJQq8KXceJKpy87jpIe2ye8MIS9BzwF/E5dEIHThePn
nm4HjcOqKfCc86dIxQ9q8nPepYlGP6MHjE24oXAg0gS1oyysbP7kt+3TiE7mrejR
hgZx4a55Y3mkSPFwvcrn1USdKEZ+sJLr2Okh3Fy1cOfq8eQN3ap/yXySPN7A7CD6
UUEirqh8S5IPVRE3HJtfwNQbXCGcgo06gT9tuXRxkn8455wo20FA1gu9VHorRTPb
yFgiHQNvBO2U5r87e9KiwmhHE74gYzsSymuM7W6mappK8leP+O2Hi9ZGabK0l8Vu
f51tSHYp9DocfGE030cJjZ9Cg+33IJXscxchdXgz+rpDw82fRglXOn7en+OWhwJD
n1n/TXVcaOpK0G1r0wdQ+MA2JLwSHDLkLhEZcOnFzN+d+/TcFD5IgS7CgKZC6cpG
C20TkHGeLbXtKC9a134m11GNTmhd8paP/kct17/U4l2+OjUCdxpGHk9wHFXJwrl3
V8f6rZqYCoP/3fqutRWJ9PueaK78q0KzkrVZYC9/gtsMKoHljoZQjbF9mTWE3C1K
tMIHOzBc5PuFJzCc2tCcKYhhZaEPSx7fJjFZhS62EFM1tgHonMUV63syKY50mHbv
TyyByRGvAThP9ejBBaoQqWN3iZu2j798cquG1fk5IRn3gc0GLbmRA4mYdpkVja7N
8VU5pt4EUjaLmYulrXYtDt5eWy8niMX/9UyZkVvkUqZrgDhLnkb9TNG1YwMofB94
CKR910shYLBGWINFQKgU7l6kpwhq2QXrfR9Kw0IK4j+waoOc1zSGEcsCBWzhjnJC
IedtgRuTcFy8A3OxI7HjJb35oslVi2Wuvp+dJ1E4qPiXPyw+ZwYSJmTwaGJDfUhi
aLwykz9PKM4g9T0PXD2sgPwfwpZzbFhkPecPxQw9OT4FtFpveiHR1tSUV8d32lBs
fNaeuBxJOT/grwRFzC29J/LJjrnQVneGgQO7VUHeBHzQn06Nmm5s3JCO2fWL6Sbx
iLOwRo315/h2SPJ5tS7GQibX6feq7pJRy4Fepc6pk2xq2jsXINvjjYhDZ28BjYsE
5ydrhIvdKwsySaP0wuXSuQLzdLt+Xd5GZ4yqaAkQ0QOW7KWZBBVWGR0r4PYPoUNP
nRM+5ZjmTWlTgs213slOcttoYhaeiq0eNYHp8Hm/00rn0Umv9lrD5hkoEJfE+rMm
FVRWsJBjvR8MCHXVVLKdipMOD/HCugfbXVRIu9BmiiDecM0U/iIQq60DXwhlgcB/
mA3/uExu0/KEGtvB31Ok+TW2wkv7Fhr4YK9rpdY+dD892s63E4PaomkOszDGFthg
bOCChTUCDqRwyel040C1KGQz3BynJW2gqzxOdMs5pqzZUpzuLx8ATdQJsW3YLp/e
dcynn+3/I6Ou8rDuxedPLFkutmE05IiyY5n+pjsauDiIvBfv4jdhDrENFTpOan4Y
Ro0iVcYp9sKzPUJKbTTMas3sftVy1cT5NTNn6X6GBWrlW7CA7pFgSr4jXMY7o1+v
xa+CeewpkCkRpfxw1JVd/R5EoNVij3VuAOWY3pTF094ct30Dg1Lj99Q99PtMSgtH
jq1WuBw3sDGtGyLqioWmJ7tJmmiab9+z4x1BU428XszzB1pMR/6sE6YDRaTwpUr7
EJY0oLk/H4solvLpcwZpDlY+6FSIGBNayRLLR4L6MzGmnVCVXeTkpyb7cJ2w0xci
OBxy6CGFhcWCwwHkcQnulpuRqjE2okvxnUm630Kq8f33EK5li0JbulgIXlGwmsYa
wD1sFLkDGh1ZN68k2SGiW/vf2LFq9lO4vwRT4ijWPTPDoPVUZ7rKfDbWC6Vo1SVt
bQNMI3uLq6imazzNdAFf8uFDMFIBqE7huUUpeARiupKWtmM4BnqxSE5nSyXv+uqh
W1mf9vdeYmhcjS7RVnejHy7u90McHBSzXYvleojywYM0L+oSwF8s0MUlDjH2efuf
lIdIml9Yl+bb2pHh44EbNybIxvIQjiSFLHNHc1IeoH8Y+UfEGEPce1oGsJiqtnGU
w/tb8VCBKy6x3kd/GJtI8X+DWY5Q8gtrviJk5bKZtz/tYTStIMRlaxwYvoVzpKje
x/JShJYXlkfaYUN+hUZCgTyd78vNAdOsIRmrJ+Gg0vQxQmC01ZVWSA6XsZyES0PQ
`protect END_PROTECTED

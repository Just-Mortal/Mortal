`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rg7NchsbzReHMoZIj/wsnZ0dejeY7IA2ielSvc93I9DYGxy1sGQZw4pRokT3wn13
2c70Dc03Snu+Gr69vTIxWDHy1E6v162utE9C3ugDiiATAR1vVSTmnOAzfsHN+zeZ
3uAwdd4Iporr+ne2qz3tsXCbt9aa5M+YbDDJO+I78/xjOKdaM7L4IMM+cukhXDOo
adPVwhGp0ga/oXx0kvLMBNK4OWmKiR4J7Vh+ETnTI9zNOWBEoXUsCc/ecAq66Ftr
Hf+JLAaq04Lb6qZdhdMS1vISlMX1nW9U3kMMBaBorlXM5lU+AWaMl5/K2UY44QJP
JL/nR3G4vMrcFSzAHYBccQTLbQbNYHfHjLNk4rui61lBWxU1hhdtrccMV7gPIGWB
n1OrStibTn3D9QZPFUmYecz6L/hDlQIr73FY+pdYwCf/2gW1MxdkXMrhXjEfSe2m
xJf+4TDCM4L1CwmUi9KzLkAGlqXPPDKZHVOMHqE4CH9y3E4AgE69owIKR0WypQ3s
EKy/EdKn43kZzgJiTQDzsqQmTzY7kbHvK+DzA+qr5ou6A6rFxAAbfCJ5tEm8maHM
hxL5PNKl2DQpeAY7kpJyWMjDKDa/3zKLmEFFgJM9KPuF4W6P+uOGj3PP0Yogefa+
W20X2ctIXFyhAPWLSxu9AzTumY4+9yDWEy9uHOgwjrZBlcnXoCyBjLdFsPfbLypN
eRay+vNSiuhqiJW0AG+XF4EUzO5uq1MLeNQAIYsuFa32AHnBtK/3bnlHlJddugWI
2ErJBUgvapeKhIggO9foODHDV2mFMDYIWc7InBkKyHBM1OCDqpfvxNb1oPyis7yh
MWd0dHT5ulfOlQTv/9rNWD66jSji0OvzycSsK8sycebLAKnGVGDNCvE51a3jG15r
DZhywkJymjMoFN+APqRP0S4QRppId+B4eYRc2Axutv7dmnlivbiVUHPvQqZpfyJW
9A0fP9zsLB/VyOgREy6MUs/mAH8/mj+JGKEohiFzrWGjFnHnekvrX+uhsee2RxsQ
Z2C+x/31ZyfIIyy9z8lJPMlz31jPwqYLf9OMTv0cUKLAQql2kl1gucZWOWzTINRI
XflnV/21sl3Q/8MOlBvi13oCLPAEspLaD1LjyMI35YRtgNbjFtGQNclCDqCEG8mh
2FJREW7jX+gBNengFG56QtMAjGyHcqbt/bF+2N7cYff4/MFHexkkUVfOiF609ru8
Ufic7T9jWohKmmwYk5v/0kR4KLAOO+oI82gXSQ4a8JVGodmExJQhFDFntieMx+Ia
Ru2JHCVPtgYz+Nrx7M2bVDVguZlm/xaSQwGvsLnaLww1G7YAzKf0ll7CWUELftYK
oltoBHjtJiUVSwSRhrhXwTBguE119MGV/Vn+z9QmGYG7xS2txNxoLpM6O7hjqrZ4
Q0tudx0uq1/rXjkeGwoIDmhCb7uwyKKsOydsSSIRr1jT8Z4v+MbOSNlj1yYqY/SN
`protect END_PROTECTED

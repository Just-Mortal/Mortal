`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
56fq+YMnW4mVsimkMNDPDLah4l1MbSCKavMEa9qh1MDZzF/txWRYovc8jz8X7X/H
mmEqeIC+7j5wSr8iJfKIy/B1oz+UPgYrSaVglwtDkc68zKcgmLJ/N97l9XjQ15tn
Ul1vf22+26CRpTOML69Ed+JNi0U1k73Ebi9WD/cSukwjorv3IcV5UJrpfz+ZC0Ev
NK18iNx4yOZm3Zm/+hr5Y/8s4H5Tl5rGUH3Hk0zCOamKob3xcJ+AzB9K41GsMrlL
9TwElGIA5eVBYOvpf+MMh/HQ68R0otxzKlRbb2N7RkK6UBS9o8AGt3CS5FJEOch3
aXfVHy4psWwWrnlo6i7Nsq7Uu2mTCWifZZDWN9QcVAey153arfpOWqCVButvWLDe
k2D8Yb36J+FVuRpumzCL/nvr/skScGX5/nK4ffJwTDWxR6MszvC03CENQtYkVkhK
VS+88WGxCIjHcAWhayJDQIGjrHND3vjsNcCAi5d+7C68DNm1YEbkNmYTyWnFMndz
VFpC2syq+k9aLxqaS4Qb0wKuwKoJT4u7EZv2rQlnPz8=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmN+uvfbrsiNTYjnCdifJqQZbjqXpDDNtXyN1IvxIFwFVGtTwT31LzgVmkMuK8Oi
J0/aBLBOGUagLEgX3onYQgQ//r4axWPV7WMVRDGMLls4jLmfjksv2pKA/SZ3rXFu
yVnD6i3dlY2uhIMOB7xHIe5F5Jc3b6FUaMPGe8qjEj5nVNbPe1IuDtqMCBpEPnZy
xWZM6lUB571FDQYOZyNJZgyeTX7TmjG6sxPgI6+0XWhToVk5dA+LByuKXfDb/p76
oRTvasxfIcDW76dA9wNNlWJYDOUkZEvZQ2b9XpraGiKmKbl2nARCw/JK45tv7KLd
ED5SvjJJCIiNX4TpO+915bybQlpbfz5CATFWdiSJ1BfVy/JXL4BGca+hV5DSTkm9
Mn0DA4FTL2lVUoiSCamMSoDzUKDWti0xbCBJ51XfiZ8zMDsrpJuR2FusIsDb57Gd
bRi364LU0ZS25eBZs2CEAEDbFpuz/EtF5gjktXyWxT4=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I73CCc1XsK6cGyLu6D2TPkDpOIGIT8r7LD4gED3/271Ihl9Q2Qzi5aJBI+xwWDqm
Q2eXCPsVACqmCK0AQgzBWEsjatBTBYScruNvLrmLRKriG4KpAvBp5yUIRHpp+2tI
56vkDint8lOQ5OOiHmd8t31D+4nT4RrsYJ/T80UoID+mvWR8P7kw8ebYu1+Y14Ns
ejh0QNZHXNQK5b67Gp1KulPyCW1x5A35/E445g8aZS9wbpO8ZN3sUr+fmDIreLQ8
mM7ndpFAwzwvFqsFVMjOxffaNFgdgwXABaGXjEVdbba2UokbKS7DHNF1YBZd0WpV
Lkfd9m04ZuCK+f/z6QW8+zaLB8OX2kmvP9VoOdF40geKRGTLmBuJrm+Gm36SyEWc
rpYTs0/BsupurD8somJiwWL3HpjGgtEjrPSdyjoArlGpX/wtMz1wGBctwLPT0NXi
UDa/cEoWoWgyb8mvTHde7CrIdcJWEkSxfAX+vW1k9qZjqzGB6QGr25ZGLFb6ux5O
t1xqjWdTqD5i917PSc3oQ8AfFxtqXWjaPHsz6ONc480U892of8XRx2/4rlvjJmHp
VCPwS3nauWQkWUB93e9+BogD+mlFKonrUTHZYSUiJFVLRI24IFDqznPyM/aKXk6b
BP1H8F8iFGFDaZJKJvnAVkamlI1+j9uW9TWVo77xmOW7OwqEjJkQ55A5MKc9/jLx
JqwjFd75YUIDYNzM7cKVtmEtl9O8AmiayG0uNKizq5E=
`protect END_PROTECTED

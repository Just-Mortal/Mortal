`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19e2nps6bVKl7ETHR8RAiAcaZ8RE6sz6r5wgjps+uKKQ+H8WcU6r4qP0mvcMv3Ja
n2Ld1k0q9brXeAmV6dUeetXte8fD/0yzGdrqOrkd7BK07IkifonzT1PP3fOblWtN
+MnGoItLD7XnGZ5P+dqQ+E6hN+SouxBFY3cm/g2jlMt8EP7ybXss0zkbN7i/Y+nw
EvqiX7SxiypkV6Nz1wmq7yqIHbK+26gg7SO3hoh76YxR1PqVQqKhZ52TUBhL4P5J
jzX8FIhpOihV7EUsBIIt0ZQnY3gTSz5zGEl6uPqD53YG6LN0SThZHeggwbFNHYmd
c1Z57ePyBsu03qbBzFAv52Gf30zRowauatXzoAyfHcNl0cWiW0xVJTEWdmnZD4lZ
6+XMD/NwTPG6C37aqqk1RXgAb2/Eo17E83ff35d6/FWIaufReHJFEhsKk+weK6hU
D5SXQt6RLOKVTl28I1LAIojXLkIH3XtJ/3RWsSfS4Mo/cVuwOlUxUQRjyO6Cdx4f
qKNA2qPWB15KKKIG4XQO7hwcE7Q0KWgkvY57CwJlpOp1z7z0UT2BwGA2OHjgVPrX
dzVYHQ2F+IdearSNtorZ11SE3SviuGgMpwQPeW/TdK9e0oiC5TPsI6dMVUxDZMOJ
aIIadrZovebwdpTxKKXjdph29qZp7W/dhC7OpudrFntpom+nfnp5/p6EDPLK/UVF
BgKGxscVER4/gw1e1N2JRTbiZsgNfNOweq6ldqSJ4RW0VcoSf/9mbpBURvKBM8Tj
k1yI4T4TfASULwIpduViYKEpnxnI2cgDmYMoOqeU2chMghWlaryLJusM9tSsimNl
zY13HrereNXwFCtrg1jYxYXZGK9QSXkjE3tO+B+FkIOSG5oAuxs3fN1nr47JV6wN
j/61OIgrBbz/bcSSUDTK97R+N7jZ4KFT++arD5Laz45AFqTeUDDZ6yOEzCMVSjMt
CFgUSmmPvTvFqGwQ7PYfT8iBC/iQmMQf9JxsEn42cFWanWuf4CXCEVqwdzuhxsOM
gIsLhNCTJOlxu8wynykPAWSbLB5WwkUmMCwXv6s2ahO7PfkFtrQ4aVTckPbsK7UO
RTZ7JYzf0ukUa3Ct0n5tQxVj1bWiN1Q28ItE0nLQsp+hW1CdXlTv4d30Uixu+Ppm
Btc4gVx0MiQ0NykIifB1FUmZxq5KXJzHbODx7TGruq0/oi3Q2gMI/A7Q9j/Hq/ix
svvWwqVjFQlCH1JgFawPAPln0EZejKVX4sL3OZ8zUKSNtrb/FacDNmKdj6TgEf3+
8XJB4pyjIFl+y/jgWdLM0e00RJLM97xn98toNDYV15q0IX5ZXoCLD4z5ACLwd6uD
aec42AnURkZT4FTfl/8G9WbDJBNjR1RYnQbQl6e1R8z0m+d/Z53bQLZ3a5zFRM+E
fDLh5D7RFdjBhU2pj5DaaO7Y+bDsEqcOzEcKhXYy55CuNf9ClCivooCVg+kQXEGo
+uUM8W4JOa/26TZogr2G4hk6HHUMJncMrZRyG7Y7B6/6VCjKJrTAf3KPRTA5C9aa
RWbPtpJIzp3dbOOZe/iNU9CWa+jpcqlJlULTzGUIJsllmZNpeO1zXE040nQiFKaU
SKpKfAVEGqw5JZd7lsOm6lAkgTuxt+2LCHfdImG/DtlQ4lIqMD/uXkcDrrBcDWM6
r/La82Sgs48mLmpq7ZvwQxK0et3teXJ8z/MDhXKk1mpE7dRVLiTeOQP7aXQb6Miy
5ByAn3XyNgTvYFfZ1LraVMsLtxTn3zfeAxvJoFxdpJ9cOp/VHsAmartHsI1wHmuU
yYqi8NIelCw/9Hae9gjYzz0guCwe8QbolRzuvM6gXAH8S5t7ukbPGTrQcU7en4EP
x+KImuY7EbJ/sKZRZdXBpEEJjfGI8RUnn1tj3XshYGpS/TwrsUJ+HMJXRRYnn9gk
7EuGkO/VOHWVYVxfubcPA7IOFz+yTs5usk59bCqf9ePVi4m7e3iNgJznI70JCZ5v
tk5I2SuiMbtNX8tYEPS9ry8vvT8tXUGe+AvubTBK5FzoDJhdM8txKv7kImAhKKAl
oLKUcQRpVd5uWvAuiw9crXZDqYaEkG3FtQUqjhiTO/pdry2ZXuWSgZVzuAIxLK0W
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEMni7eY8Lmkrnfuc0eb1c/EQ3lZaXcOtSLw3HCqT6u/mYdvOri/uYzO0IiCPdjp
HOBXFA+IyjXMI5gKmyWSSy8eGdUl1D6789laT3N6ZueSpYBFXLKdhnoApR/C9AMU
/LpKgW1CDQyV+m0ixATtU/FaDLKt7GeQo9iYm07XPNVWSjXpu73WGPPQqprZ0nWi
z2QM4mUvP6FoTUqBufvEkuyjYXapr20Cr+XEmu05gUhdLv5TH3DSPpcFBoBSX2Yp
kJFKU8RzTaCFKTZflj75350q40NsBnOFdBFHXHyhGARG/JbGsIgsF0j47W6vEe6n
3WYWSQGbMslhK8PNc7uRU5iDnrHHO3kgxD3zDrMts/CekAo8LT4K9vRgLXO38U6f
en3i7MRjYBhbwwGRvceqjrSst+Ro3pXQwH5qlKREZDvT27C/pXVAAgBFFD8dL/5n
DJXcOcUOKCNE8P9NR+wi4PpFdhfps9JQDPK6SaDWsu21GoxhHFQ0E4r+oi+b5HM/
LDfsljSuCbKjVAvbw9Zao/cLzm9NJTsNSiiBPTqxZqpVKZCTH9qwQibOZqK//ked
3oDt8RtaxOMwuq/xAgaccURGT0WDVMA6NIkI5JsWCg8xz2mUgzfUZIcXk/DzG1o1
kRvzOsPGwzPP9P6svhc0XF9nGnO8eaCnUoW2eCOlxZkEfyb/wRlJa7U9tNIB4GCh
jTkpJM5aT/MUdUMgOJS+HNjKb3613lFRR5U2o9/gs4+ry7QGCzVIAWaZC/1jGUoc
YkfNaim7VlFG7wuLAaSy1a1K/61kt7YRPO6Lh1JwNsQ=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNg7yEQkTe58IrDAJwCShdaY25/z5nIXf3ZbAVRYVJi8mtY6g8LUO2eVTXH4fNcn
aGHeOg89xF8bf1bywx0ud+FRwR/w4Fo2CZ64g94jq7UF2Nm2ZdAS76JDpvK2PoVt
aV9IxuJNemEZJlm5aDRsI+f0k4HKnaoteGaBGmRjqc39X2LYmluBuXixUNbmRyFX
tZ7/gKdr1OZGTH/GZWKnlckNtM5Vo4QpS8wKx4qigddkKrqiB/25f2BmUyYn1scg
h18w5z5quzpYF9yrBpvWEQkvAe5Y/Ilmkf9nIGataYRQ+npJhfXLdhSstfZgU0qH
EQ612garSJnnl76j+Ii2/rWRYfEjagySQ1oPkYZRGGnmBHF3HDFzvTxcR5BIVsWS
5mZaei1U986bOvGMT39KtToeRmDvlf/X4JalK9sZi8w3wW1TCktqwMqkWQQ/VhcS
h8++2sBh3d0r9y9V7PaKoYbvedlFGrJVa2LEdoS0vMTI74gKql574/g8+X66w5k9
yyqiMXyLLrHAGvVY2OzjG/MG98vtyIADBwAIZJ3mPFqBG0WWqJ6pn00UT+++PoEZ
J0MjuoNNpnxSTAQJAB9mvCBh2ntAMPSm3grLO9nIBRV2cIrW2+zgtSNZhJ4mdp0Q
CXGdMehjjj4I/zqn26dstsHtR30/sqFMCDcNO1O16lRqx0iRoruDQNsMdXr8s5Q2
U/l6zQo19IIGAQDkXBdmbXJAKCAyybYQue/w7Sx5qeN7Nh58rqosIRO25O0OdG+3
nG5YJO1vznGKae6W9OgNiftPLY5o/7ijEB4Ys5RT9wzUVnvq1Emgb4wzba8GrMA8
oykmA7GunP8kNOeE6NZUjoulDqaoojr77to6h65WEU7x/la4TbL67BImrDLoBn3W
gYJFbd2hqVKfkfV8O8zA2dAjT9exQMqFsLrPZO6xVe28MctQw/dLF1B5FxtPafxA
EQv9jF+lV3g38iFGKztuHofCkm+/kvvnPFNgeAzuXe4=
`protect END_PROTECTED

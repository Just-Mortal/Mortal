`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fPQI4aAz4v3yxj/x7ysaiAilfmZkdGkJRAx1WCYuRaQHMHFVizDbs4/bI5oxVOP
ocaH9U76EKmDYeIn7NoBCfNM40uSj/OuAmZJu6O1FRAzhq1lPh6EcGLXQp6+yH24
hAhLJubbd0UCVITUJV0WIVIywrbp9AJQjSHh7J3jXdALQV6SrohgAO88E4WrCo0W
VHONa7/g2gUVCQZzHFwzOGdSbnmtbnyt1HySIerI+nVIxHN+KsGsO51q3+Iq2qTC
Oz4TpjawkNAQX0Bl4sxfnE2FPJ6kG6dg2b9EDei7pUTb4ONlS64QfOUAfge8yol+
yk6ZqI7/TUvQ1NsI4dNbV2SZmK+Y5XXKxY7BTd7dV4hG62OBcqvLGBKw3JC9far5
NMQG8UcXylHxv1wN/ihy/9Pji3LnnKEpdk8rtQk9lyGz6fhXWFxayCgSiuMQyEla
TjSRvMBgjSJJezqixeMleIrCm+5KfkKrQWJR3aWrQNUSRp6ebbAl0rL3ZNXDMYJu
tY1OjYyNGDx0kVxfunWOLTdWE/EcGdJi29F9Gh5OKqECuo8NIVCsnFkHYzPHglpd
3VBnviPj6s92h4tZbY+vWJca5Ljv8+WwoDDE8/dhPyaygE1gvsm1TqaMvWgAm/Jn
uMuSq7gYMCnMDUQ6xzR6MJ2iQuh7GGeJDdt1KuzzoewMNH+Qjn18hlss8APAIgp8
KTPa1mvyfhxrY74rbpWQ+6MEC9pvJxYj73P7sfgnPGBSjeHjs8NoEsnCNJWtswuv
2fQBzGU/EzITiJ/8iQtgA72tAOF8IqhGwMn1KlHcBEtqvCMcrMXo7b+L8XMyFsR2
FJGEIkm5+6iSEfMi5FItPkmNoGUmlTmvphz8mth26uQII8mBIstcEO2w9WsbiRY7
HmXCFX+eYMelnfg31iuR81CsBu4da9v4UBaF+TVHmXjoQ2ALzkGL6K0XTjp0wXVf
weF8yOnU1RZhubT/FmxOvQlF1TgdPiSJzufz+dFWNlT+pSfUO4O+2d30SCw2sYh5
so+17GOMBoNthycZPBgYw1eNtUPBthBkKlV+S25RTJQmPaZ02lPTT9PiQdQ+nLP9
mJAB6WpH0gXL5GY01d/IKQZGpx8kB0KRBUfpnZRWyCOEKeven6Ve7vx/1k9/mSj1
cXP5kv+BYbe+p3ZKtsoe0hCmfvA0hZ8VKfdwE5hS8COYPoDFX1fYBmCTFpBw29kM
x5X2RJNmaJ++wtcw+4aiyG0yJvwISm1RqgN5uZDpBbFpIDyO2pFvlEmt55NOXg4p
2cihmEmqbWk3r31YprTgpU2/nkTC7YvuvlI2WMdc44J0SsNnCRmZBxly2aYN7c3y
OC7SFwNhopt8XS/aOzcPYZlwKNq4GIpBB4jonlopM3h+PGaxaxcT6DM4MJZW9vdF
yLLMG4YNLNkxYefBj7lVJ1GzuV96sPgZFXFTEmwiDDPLGE+CJL78PogTr7hksFGk
Z5sCPkpAMbEXQhch2TiUOjYr0nJbHTlgLhqzedVdEsD8+X+RY2tXbqQXwLfm6QYJ
+aVjJFotbC3KKWAemo4zii6uLI7jDbT1IfJHdw5fVciDkdqdfRF5JqVkraOL0vqC
feJA7A0qEG/H2/JTFq2GITL8UmyU3sT9SEdz0v3TfphCI6MNz5JlnsPOBVyi8TqN
ar4mFp1x/GiWWQbMFL/wB2PNoVQUu/VyBUfqF+i56YpuqB+b569JczC7fzK79SZu
N8td2tFAx5uh/BA/T766d3MGJN175TztLdoMw9nobtqFB9FP9GRx+vxIhhWpcysG
Ziw/1x13VSs2aLe3vuh+AsB3Ba79awSR0aMrFFzvI0AlQhWsAyN3m4dyD2ym702n
XUnOt6S2KZ1Y95vl3wj0Yq0gnX3L2yPzFHuAsazIJbXMD0z4aBkDKhsghbIv13Y5
QO43rlmFWGZX6QD6dYb3zX0Ndp9Q2wDZIuYaRQmfSMIVj5zBRcz4NDKHJoEkBRNl
bih/mZcoP7k2QRVz5hnydVnlwloLZ8q0radzGpBhgDAPX2c5Kp6PNllxz32mnpxN
ShGeKf20qOOosW54KisUsfkPDhxs+D7oXz89tsgDwsLtOIFlN1oV22WPVNL51nf1
kMl9P5V7uW0l8qSJJjP+sjmEsrFvegQqaYlzBL0V7+3mMk994jlH0GkK1k/USLk1
7zpp+yKWJbwuVy2ID1RZsI+8P2loYVn+PUi/dy7dAN3q9STacLlI3E/NDcOpYdJr
g/E8AyuyGTVjUGuxy8IWMDicfx2yf5C8ysAn2UdaDrca5EnMObZWuOa5FfFec/Ae
IwvTRAfs2W0JZKFfF/hlYjAmUrOFfXQQejWuWrDlYdZToMXCG2a8xAcETabk4uK3
wXFQuJDQdkEpBJznLgMo5XyI98zgyjOTBzvmrXFV7p8WHeAasXPFCzudv3snT6yA
WHYKtWQ1qkSyHM9RYedaPfUjbjRMz58Ex0GtgBmtU/qjtkNTFYIE34+0SXvSTN3E
LnrGeJ5WiRGvhDhQjvMlVs2rDm4MuQfCG5YqplULFd9sFCXlueDsYLVz4X0xjrB8
w1siLoNOef983+0sxZrydDVRXcP0QshUchaV0u40AlTQBkiE20VVz00SQtFzn5MH
yw9A9D6+EDmJoYEhz/mWxu/EEHDGISC5SvXH2MO3geGz3V40UkPjJObv2aUBIqJm
JccG5GSJy/yroQ38vL41yhCk0NZctyaCmTXxEJ5AZLiz4bcWLX8o+vFaj7jV0DoJ
SClcmpDP6FsKvpzslSja2N+IjU7gTRpoBUcoNW0aAtRCmS+qvcOifpusK5bnfE2E
pIBxSTeNiSiPJRD8xVyRF1MAuGa0BDqGj0L7XtMdRYnCK9f4dMdgog2xRZgeFmZP
iOg3fyIjgzDtRGPGjt6Cq50R0mJ5B3KiIeS0Nv07lITC4xE9t9wHQmm9GRiS6ycH
GBbz8VE8aRVT+y/FEYHXMUAfsICJvtoptSL8fKGUTHIbTwrAFfbFtql9VVNDfb9+
xNntbBnREgZfxBEFc0qMCB+Wh+oJbCKtFUj2kYFEA0ABAD8ncUV3Jrzjg6Po3dkg
UgyCEmorAJsjtRwC7ZQuohBeLoTdVojJCRcp2ZJ4DtrBytHuU/0yH9Td2I/eWtEY
fCmYFOh0GTRDcHYaBT8jETuQxkbYl/UrrLGJZDUuwG4hV2XDwX6bBHcrlI5x2/4c
6MbOP1RkYuuLkNiPTNgbfD+d1nb4rSbZCGBaEi9N1k5jVls+GsHzvR/KKrlNYEhD
7bsmjXQmP+C3EVL3MJ4uzTqZQl0SNoZJPpwKHUGIO31uat/IWOd0OVXw65FBK87E
UWz7FMguQOhvy6YVsUXPALwBjuk2OnJjknYIdcRYnsCAYd+FIkm2pwDOScZpK1xm
3p5VvJ1aAzs6oHvaBoliae3XMnkj7g04Zp6yU47I025IwhILwH+0Y1MkfLmDUKjE
HUbSN6cB7XcSZ71NYRu94A5UHioEzxEjmEvFqs4jbVxSiUGcuX1kDMpDid2XsxWX
hre+uthunc50wl3iywrBOgeLjlKBO+xKGGtTC+u1CbNArYomr7qwiRQc/Hqpu1N8
3qPfJegowzU9z8rHgJc0AW78RRdeblSfgjnAMDwGZ0BzUTVcymz+xPATqh0DIDHh
tIHX/gOZhpPNPVjI+lAr8Nn7wIICEbTEcJihLI2z8kpEnhZq3vnAN9Ybqo0ARjwJ
pg+aE1YtF3Q0Edi8qrm1JWV7WH/aiOMCpsF2vaTEgEco1rlXP8JycBXtNf3y0S5A
8NXLJutgP1qO6kSSxYGLFg9Gnfe6VJYIZ9VtO5CigxZPl2FQJ3kiNzJCfHA0qgEF
dXqTxqFLUSKoX2ILqeSC3zNVcSlCQL8sHh54L0HGD+yCE9nSHVCR3h/D59hdIaL0
vVJmO1q/QYqH9pXiwAY0WgLZFtmp6Vkf/CJgjsKbKRLGqZZ8MugY+vlHnkVbnt/X
PhtRHw9iVPmZFKpfcmYNlX6QxNa01wS7IdIDvLGKLaxbyk6Wtm40l/fmxt+Jso17
3Qn7CPWJlfxcJ7qoGbo+zgPxWWNQYWkCEqVtpu2AZRIGzgFEbTmYiL2j2hRwmvBu
NrIjnNODGi1U+4hxfhe2CixeCSzXTpQjnQNg/+UZVFIlcbS4Na39y4MhZjAo8cdi
WS2JarCnxO/oRMRbgWbSE40PH9q4mIofHw5r1itrk2PtNxfGl8M8iGpSJ5uYEOpp
2oNgpJEgThL8C7vNdh3J+u042cKQVD2SkJEpZQSbAeq60T2FQ6YJeAPXqRN9GZAT
pDR8vCyn5KG3/SEVS33ETVL2V6Osm3XsJsCaqmaDkurUTyJ2TKQzpzCTIz2tiAYU
T8dn7MJ+O6lze7mJPvyynYCVZUQAAwrTz3gUNIcSvxIxcjrkktMTSB8iLx7wfnL0
aR3LY8TrZOkV2OH1K06rs6FnB4+s5qlY5mck5/lxUhxL/JYcxxZ5qMma0GA2iXc3
OM086Z6h34gAsE5O5kDDhsTsPrKqNpLM7+FeWQdMNi0B3lCUrAmx47CqzcLM9jwL
1iPszX/A+Scl2RKnZ+i3a4qgQnD2TL7blIWg7kw0AOL7ErnF9UUU7SQ5Z9o5Hqhx
r9oaVCUgJlFVgLK32YydMl+rgYNIX5nvqQ+AIPDBAxQXHy7kQ3UnB5Yk4wPbeAFc
Rjw0BOUTMllS0izvq0ghjiv/Ktzxnsos1/VsuwF6Fq+SmWVu+d3DTKoHB9tjojcB
eWVwjoWGzqiGsn970ohOqpJv3MNmITA1wjBVqh/d8Jh8NQ1R+CEA4FqTZsV8YvlO
3hhGrlML0onKSd+XQwxDdy+GrQ+JEEbg42HVSNIg5mdKxOQfr+Qle+modphzTOtk
YnSKv8I9JIVTWuKR1CVj8Hf2YHZqdG+UgVz5a4oXI1O44XrOXGnzXIqAZgjLz26V
QzH2JC2p4xkoUZ+H6GY4IVApZyuNsU91mQSAdss+4VKikdkfon4DHvP9M39dO4dY
zK3UXVnLe2qA3db870k9vWIL2LdDyb1hLnVEChUjiilzblESNd2zsJ4S0DMMLfkY
EyCQcslFubAqdm4fpqQMpZe7SKPvVLS6aSqwfmD7Vw9glcpMYTrkuFgHzjZVOQiN
haGc/GuCuzYdL/E0mIZm3AuDJ//FTFf9foPMlwUXxEHAP8y0lt9jWDXWze/nM3YO
jswYx4gP11SIBuuw2E2AUMTngWiugIr5anPBq/WvcM7rqGpVRLXErikGLdkx9Rgy
6jSXkk/CEEFadFYKwJXH4g1Zf0zWL9hDS6mrtyTXX+Om1f19QBoZ+HCegpVlPJ+T
taxOTvFEmh7a+FmjMc5zjfV0QqEeEFBFPZ4Xy+N1MEzBmmuWUGXqSYjvParzTtdu
EoziggPg6TiKD4JHTTdJBtsixyvV9f7Blr8Lcmx77Gg9cprEuhiRvBorVhMn3C6g
ZBYRPPI2vQsEecKUORgMHVcIxJzGeM0IuyRsybUtXfVZuf1S1K317SwYpF7XCbnA
YCFR4V6B8KwyCxLp/viwStLFT7glF8TBbmbp/zK1TVrok9e9lLXjtrrGVGMJWAO6
JdALAiyih7rgw/kXOEU1x9x5S81VXvol6GgYWqyXKC/vYsbzS/g3XwJqOQlOWohl
rgIKA48LMe4dlslRaMbmouAhV7S0egbwiq8fTRRc1szX7JtM3fmOcOjInHBxT9fv
M6FUxqbpdihiPtK4TDHDl6yy+QZbgcPOYXNHZtsmr6KPWeMhlB/DmnNHotUPZdJX
V0VXsmYN+Z6HuR2qH3j+V2vN1EBwFtvDlVkQxHdqWDgYOQklPFQDOhpSu6SCjffe
LEhE5ay7J1Ag/13Nt9hvUVXrGI3u8xst/SyO/mxD0shKl7WtADkG67t0m/9tkVJN
RvlUca4tI/lqq0L0zsmJgdqmKaDXa/OVIFRDQozBVdEVBwfqCDwpmE+TyoSZaX1P
noR95kVQFLts3PZ4CxYmm93DQwnd1zR8R007PLkJvLnbbJjERXV9It8aatxJX/dO
88mJ7wMsGEyXlI6+Tq3owMP24h6XZ71rm5XeqkYX9rTpoAEdp0NTql9Cyty+styl
/nqC8wv/qDIlThJzbRqLfBkw+pAikMI+xCvfd7sCD2rJSOSsUHVrGz+LhDVxM5tE
z6NKpx8wLHmPyyJKkRyGgI1tl7mLY57Cm8ViivSG6RV4SR2+T4WEzIzNWzK6QUzH
N1P9n/KBaMOjCGcOqHhnzu/erCdQuKAkSLZOZTHAU3BNU1cBd8OTsbBn5d7XD8DV
5X8lJqh/WQG2uAzsvIuBPDVdyNFxzQ0uIP5sq0bOMGEiybN/u1EFIrsdNb0gHlmM
jDesL5vcUOzKWTqh6hYnElR2Y3cS9HrVRxQN2YjqG4dvIEyd00sdeRvxSh97F9RL
2fMTxnit/2fBCoHHSgub+Z+t11SqtS295gc/ezpDECLQJTohpteT1RJOXllP1y9K
fHFWV9bsZBBlabOozRxGlY6Pm7zaB1f7f9swXJM+ACiWvQD5JkArFKwwec9pwDkD
m8Ah2NnGq9finSw0YCx/24Ua1E9W8x4m7UNI9sMwqrqUlaiL62fxhYAkjMk5eAUO
mvWVu99c/8gPcdhZ+BZl4EbLlbAUniY4OGxesXvgaOwSyDU4l3jypNWpvV/YqB23
LvP87LbemcijFLMIp0nNVwTnPbId1hXu7V2sPWieXTTf9fO9UuONj5swRARdv8J9
ux1y/qYPqgg9L7SYzNJx1fDAD3YTtJoe+RC+gRSrp29qnrvVY1TzmzzfZpCsU5Wz
dzoiOlDcA/L1uoaPQ3Dw07V3UUPsZ0NvHQS8zPtoRTnhbNlhWWLoPbgOdBBsAsPe
9NApqca6N3Cs+7TwooIHPVLIe33mLkQYu1RpWACc1RATbEU31KLZDg9D4JxPLx9n
Z15jQFOKZEO2td+VJTfecxDN1Loco+OW7yUtLEzy6XeLvAdxwdyaZmHbQaFT0kh8
q2LALlM7h2BICJIYeEC7kRAjiNYBpsBGKNYjrMIUDui519ExNgFrlFHW3b/kRFb5
BfMw1iqDuWig05Zo2jkfF93exKsUHIX/gzsSVL+R4S9p4fataw8kwJ9xvHOygHyF
vcoIOH5IM6ArjGjeXvgYu+n84Qd4TO6uZ+5limcn7ev60jRk6bLblMuN7iw+FDVj
XT55F30Mo2rOPx27+XU/4PNuW8rKGP8jcblgaX9WqFv/eRlTRLURwoqt+qgnbQdA
OiHFGXpmXNFqDz6CWa7WyEuOcw/IQpu0Yeae3neFJ2FeS6jUGBKPbPwBjf2/Ko5d
HFGIiB5qmDE3kLpKJQkBXL+xt2yRgkl1hOP7usmUTLYMvwriIjO6GrVC7RDINbjf
jspDY2gmSriKPacURj7t5S9mz1x1lFb9P+zLYcTQLcrg+OCbqVciL7CAncvp7hlj
WA+P/oHTEtQ+inxRSvzEg4rQwAupzPovWKOh73W2A8khugctQrFbY1p8CCkIzf7/
EfdwLNDZpkIfd7xi108KtM3oVi/Ku+0d0WFTeAi8acWWmEKhGi24QmXqC7Q+n1Am
D/8kh1WI8TxwaFE1ICyxDhvIlKiLVcHJgBjoqH3mYSRAnJqN8WnLM61y/2uLxCqA
3Jv7oL3yIpwKTLNm6ZmhFC00pUpMwBz+JiAv0gTsz001GvUsrTt5Q2u7vGfvZItm
oL5hxa/kUcGSLQpGomWDoNIR9OgqxQyR5UMOWUiklvhySgVFGXiDwDxqcUfg+kI5
qHBNjoodV6grmIbzqOOD1R73n7BXd8+mbZjjbf+m//N/ln6jdLV2inKyMW0bXYA3
sQozOkL3itQLEM5XHs5XslC7gxXnKCQ/FCRiha5ZfBCmEEPrxBgNwQyayJu76wi1
qv3+rTpdXP3tI+H3D5HWeCjtUe0Giifxi28ZuzjyuBFnHJ61FyXRiDxFreJlLS5h
lI7Mm41MxYUvg939wg9Xd++dtl/agMXJCoA9zxY5SRxpl0ME7BYSTK1u3/K1ycOc
SS6k3lJWV1d/v7QtJCyF5CoEanQbJ/LKbEAQbOBr7BX0rRygSUM8qWsV8KO0bMdP
wG+3+6vaLXQsXUvoez+Z6+77XlsGFHrGLl7cYDOzhuSYjpJlrRdOi+MszFqp/UTc
5Xt10v8g3wPw8qdBTcs5ckPORWF8Xh38FHNFC4Fxuviv87mgkKrhH4bPs9VnoJgW
bCZ9AalSq5jM5W/SiHrH6Nfai5BmOY+w11wbpuU55ycXtbrZwycqi73WHSCqt7E9
/0yw2rYjXQcl2Z2S2B/SbXWZiA/bwwygpG3EUizY4tTCqFlcmPprb2JhDund70c4
yXSm0G7KDI4Ug4ipug/www/NlSrBcc5d4IGSbRtB0w2AEYKClnEJ4vbYJrDUO3YD
fJEAXktu62obVwqcq3j2ksPQOjy3W3pXOLEj9U2WtXeb7ysyG+DZxurfoBi4W9XM
KUF1676xT2WBbuoiKbetqtSYiv2EfjvzAmisNekqSy7gxqfcdiA+JlWNziwkRPKK
9yw4FGpjii3gKdnyYqPLLVZdVsS15Vrf3+6Q4KwY9XOrKpErpFGtkf9z26JASQ41
EgE3Wca/vt2eEgR3uSqFUqVEcqMnPdvrOkLyjmA9SQ/s7PTV8gIuLZnpNq86+1Ip
MX/6wP0JvMwfOT7CgpBf1qQNFx51AzNO8TOCtkiZPGQKQPqsVuVgoZYW/1m6kYJx
GJvUHIrvrGRe1e+VJTu2+Ff3XhhX9Lb8NSMXsdXj2DeQlHwpE7q2y01eJl4HRc8m
dU4IHGFAK84tUXkfDKlSdMIX/TNz9vEKuVnu4aIixcWfSeNpg2gefCNYiMiJ8OeQ
+GvLmRFRkAbmvAvILmzX9ZK7SHxynLJcumeY8DSuC8aoxmzR8bPhyeP9aDhB9C1N
i/djNW2x9K5rRC/dautpWTyvtjUlyfoY1PID7uLdl6ePrpC0rCroLLMrRZil7WhW
kxDHku0sYhelzhOj0LTeRZYILLZOVKAa5VHVsfIeU/47fO4QJbL0B52BRTlRHuMU
Vdzl85dwbbtH0IrpxoZhd97s7juVE2P379uNfghgInPIzLRJHsgQxtvdcWBi+1fS
geRxHtjO5li/n7JLJ0+INCypz8u44iNOOlNEwywmKJA6/H0aEpvhyolX7DupWwol
GIi6P24D22XiqY5XsjpWTpc9fsujjzV8GdlotD+B5te7XWi6FtQjljcLnSiyDBD4
iTR3ue3UAM+qbZ3OG6NfTnZzzANKf7dDC4j98r5PrkpN571OzR27Kmg30Gkft7nJ
ZxWfSJfPSd1fm/bvgrHpmA77daPJHlHVtLNaySqN4wNz9yHypZcejsnYFAD3Kmsn
jih5dVX76qc4fo0TIOPev5ycacIp6f6bBKM3DHTr55pOZSZv7gQJXFncmlUYpJaO
3qkOqAlM3ob8isWyHldFxu23qRlEyZk1qSjHI3hAi+r9KncVTQvMrSGn+eqetMoa
8a7GME5V/J3P6mKKig+V2hWOzI/w7c8ZAUv4v229gTKvphKgQZAhcbPX6vpJjoVY
Y/TbhZ1DvWJazIsZCHglfkYpQwUPWSVbmU7Cns6pJm5A5deR/BycvcI4enNHY2KM
uXVQWn2Ve2PaNP13RcZ9pTJlaHxGXpEnpiFpNM8vpuiQbKuXWD8tivRBhA7WxMTD
jvU5vtXTTvCiFMvfc1R9YCKrdCrWY2pL8163HPB5hh/VAQybYkYyOXg5tyF+qPhy
4scp7PuxY1zr6XWg9s60ZGNFlKDbOCP9QpJc60Q1I5j0RXG6BCu19k24XYEFKFhW
XqcUER7n4k4oRI/z/FlZTdWKCQrWwou0LnfvNDdIqsZ0WUAs18sv1qkwrfUTomk4
m4BtClVRVGkhWscSq55Yxycwo5ATMbnp7fFOfAj/nLbY1x3m0gqz+6JyziHQ00Q7
/3LNIOE+ZkPz3OWFJPGPPOSWtTeAbZuZm6Almor+/Cr5Ifg8tCckK9vhyVFLUiN0
P+naQ5zgg0DPiexyuSIvPz0Xsw6cQKmb8Y6FoBe+sWBO5FxkVPWFqJ9ILjalkbWk
SJD9+FniCC2rkWFNKe1dj2H0pdOiNxoN72+V7OPrX2wjGJcgbgZQFcDmrtoK7fEg
BoSmCcQLHmmhYi7o8ZN7J2OFPdBx2aSdLb0PYztzqLC+KP8QAHa6UbMDZ2DqWooy
DTIh0CoggDGYHQyAQvpw5b1ub3jiJXhiSG5ebR4sVdF2vy9H3hTgpc4FoGf819Kt
oW2MXje1W0vRbGDkVuC+6FRgrrWcV71hkvgVSbZa5KPHtQgfGWXWHOlok/ubND6u
lwj/x5qtTibqAJVJyRY/A1V8fGebQG9kUfl53cXqBjXWgYJPzj4EHanciXHPV2Wi
Cy7lA6Wqu1CcCRu4RkfDJRm17Pn6YK2Uscj266Y+ws9ZKqBG82YeFs5J/4Rw1rIC
oSz8XJeX06HHTcSqjzmnRqVmgG2cl2qfkXCHGfBQSB9Z1X6/Feb6M1kCJEry45wY
1RgDaVdEhXBH0kHBHhozpWdLS8NmO2lHkT8dsFfbSHyh+ves+EfityjnP5pRD0zG
QURLWxDF6KuX5Kr6+cNeRQuaLOn0OD4x0BQbdbTf7sY6vTCVW+tIhevG85DlQ9rN
+x52/2FvpHmddlgusVNZhBDAfXixJmz7xyojfI+7kYXHPTFawNRLEXDuf3nHiI7r
TiYAo64KVwFUYAYX4as8h8aCEywwWJSwahkQulSSEkvPS/irmVwKZ0+lpPAwzgvr
k+PAzEnC6q5wtPviglc/koPwcY44/hDz339rhW6MebqYQeCVfExGk4GHXuhEtmjK
++VuDWWiFbSXCLELB0PmU6eyDZMZ0kCgrDCkDEnnjA88r2zPgpaBOf+s3NB0+RvB
cKISY4yqFDVGjAdxJ0296198HchAAdmPaPrv3EgjGJ0XarVMy1rtTiOqEIxcJDNF
IufgrXpOEw8+8J2qO9pVGzq/jmcsWheyyCT3YZUAorwRz9NeAhzk64OHOPwboFa7
lWakuNebjFX1v8i6lVyACqDXMIpst9XVS/tsdkD5H+48xWBZnNojBQgGP9ULMflJ
23Pie8dq7SmlXKL9UspDsDNJ2GEPd1+YnznO8WpBF41X0yOmnLZNFCYR9S1xpDwW
nJsmFE7NLM7JxaCfyq2mwmy+QmHSqmvTcIhGe2/JFTDm7+ORSgWqMVAzH0ly5tDv
5WPtqafq1uc4k8Gev9+hA1l68jnoCmc83dV0+i7sC9jMowwoXQGXQqMapYbk6NYT
mZY62PY2OlJbD//k1zZn8c4zRwhSwPtKmks40MYvJJe1xWOwDrtuSanQSt/nSwXf
ppkm6pbCp2pcw25BxA2rtr7D8rUH1LGCbMtLjxVq9aEK7WjnmvoahlLnOEL99KZF
4HgA08tY3lpy8vQ8bzjj2q4kcwm/MfQfckniNi3Xny4jjDHS8TTQLqE1r7NaJrRD
RhhQ7X5iOEIvmInbLhQFU0+i+9ktuZv2oAMArvVDzfj7A/K1AvzcehbAYtuGaWJK
giwguBUf4GNLWpH385MLVTEWsJACqYEY9kMZjRAb7Z8ylfuVevupZ3MZgpEBgQ0B
yjMRIp2WKQ2IfVstz2OYvC4qhZhj8NONSrd4ZDcenruA6f/xLXEQdDNVsBR9JrPe
ShiONJ/1w9FnNlYL2z00RIXOyogdVF56zgq68/ofPfGQy6RD7tcrI0JyuFSv4+y9
14ddqpvr5Wi177Sivba+vO+jfnf5B2ptnm4MMm0jpAcdMrgYKLK9b8t4WuJ7RKDv
3rNk2+2guqJ3tnDUQVGYZ9NFK2fVg37CGIfdmv/UnelAjFg3qXflQ0KkwAHIWmaK
G//h/WkXsHiw2SvGM9ZV7MabzDi4mVoPQ1W7uDdd+Cca5UdFMhBjBlLgIRlR1NDE
xnSHz+Vatvpv9Tj+S78SOYZ/qJMUEmyjhYR9QF8/loBHucp/jZvRJvp+IYxpNZff
nse3SnaCbRZv8fMMZHa38CfAzBzqHVV0S2DUrpgL9tGuUPH18ureZj3AaHSQSeMT
JaSpDerZKgMax82DyyEDyFaTKkzMx+0gRjdYU8zPEs8bcccwuDbNhIH1mrOeH95A
zXocXK+wAsMUsFyhmeBw1pO2HMfh7hGqroeuuMhbSqn8apsDp0iagtsFjsbDtPjw
HqKVV2Mv41eHrSvkK97RromzVxUwXHJaiH4CnZ8FYOJ0oDB37HE1CZjGiT+y2U/x
jSMRDGYb7JHfRXWeNlk94zW11QN1uusKAIkm6wMd/zcN3Fcr0QCesIGIa7bf5t/7
giyUaCnPbiki1yhGm8x8h5Gar6vqAA04ESv0ivXpwYvOcHClTzv9BlS/m2xiZVKD
clcwQ1g5BpQbILqyYyItaU0W2DPqpI7ugowfDEPXKTvTbwL0kg5CZ1YqIhGdttv3
C2LQExnxuFRouM7oHUnVGGTwqlyLhYX89a700HaqRAaOz1AIGEV+UF/NwDutskvu
anJcj4/oSrPxYVUvbGA8A0/RGVAriwXnx46zXftUNTEr3wjrL9be2g+w/6E5HH1H
bjOgFs6v6d8wHiqLnLplshW/YN6obK2bn7jGf2OJSYpDpRMfyu4XYQXyf3VvGCCQ
hAS95mHBgdero8P+G2ViLMI2GqRWjIolQf5L4KLbl9ZzkTB6kItyHRFWI/1VgNGU
wHxIp6MYWRl5c03HRnQGop3bJ5z8ixrcoMJFg4/Y36LMEq8JpybhbTzOenk8Yz2P
b5L6ynuvd1Aw9HRjUnnuvm3sekybKDOeGJG1LFvHvLxAmAI037nivpP9fGVIC7yn
JJkTKq473sy0shYI0xBC1WGzgoChZ1DKnC1HxmgcifMpx5kN1dIf5z90u2k3BW+d
9ki0sefcV7+q8L3A4vEnswaeRMO0GQZbAuOSRmJ3IiWQLHg/uzwtZsLailMG72kl
ZjKAYEmkGBkU6rLZwfNrMNMj9nyg4G+lmJanuihIp2At5Du/AmKsA3ABu8OElLSD
JAnqrO13rTlJQorW3qghvwOrs+42nl/Z+5z3n98cjn05GeoFWZY8E/gcc30Pdwoa
AF4HzTGWRSBkSjGbsuRPCQnvFRT3tNWXRNfpIsroV9L74GnFTnZJSBPKMwC75R7S
GS0NB1RqM7TrPHJd59PC4v38w33hVoc0gU+5RDWY5ikbVdW0zeiTRRaAqZeE10fM
oWi2Bkod6S/nK0cV0Y8NE/xsxr3+MOtLkrs9uk94ww7jzKHqmFs6wuXRL1aRyR/z
meqsHF8DPzwChkOKhzBeknBBfdXcTqB/XaaleJ2y9yVs6dNYAF47WYLRpWqGHqyn
EwaGVJVhZRCFuEf5RXquiGACdv3sWGGotVfZtpvXr29HpoBhdpGCFbRgEufCLQwu
PMa2yNHufZe6U6hYVxY7k2/9OltIGnt5JpyDIn3E7PRjcl9jE+XAw5gCv+kceZtI
6LYA1GBgZwLxBB7gUWot2NoGNCUYI9ED1SVGciFTIHHuYc6L8E6YqIzVTWYmyO67
lEvqP0mQ4I/ESm1hhtOttEJEe2qHvx54bnnwcVPDere702wddyxKL6v6LpgPn22i
S5G7IZkc/QGNzUTwjZsP5ZGTR0vYl+mRTstQBOy5CT21JEr0vzkOBeEfxiaxTRuE
nEcwfGixT2lHgixKe9wHD6Zty1hkXhY3o8ctdIb1y0bt9p+KSQZdiOvBC+SLGm2s
cINua00oFa1ox0opk1lEmpPffJAm9e4XzWdhuoII/gNwmTgLq/rpfELT/t3Yf9Re
Pfjrb0XuToYArW8EBaFHgjxbD4MGr9igl0jnbW+OafkQkpVzrH95NW/5fs/oCmMX
JY2YlhbB7g1iO13iaANUoW/EiW+LbHD2ILFoYQQJXGwuqnML5GMTb5oeFl1/6PCm
75KqJKuKpxvppwhuBSbRtnwbL1b51uaQ3Vp1L531aE7KtJ/uZVKsNaLnals2a6gS
arcHYpc0Jd1wg28ONJZPpRhe7XwS+dFybNgssJBJ4GNVs7S6HbtFRysKXLdJbfXY
gLgUHKLkAmyGJfgJHOa7nSoAMxQK2pFAKLHMHu7oM/2djzDmTWL3xrrlg+ADKJ+9
HoOahxGREYFWttl3swSpt7o5ySz9KS3n/VOx3GTsIF6vgwBSXa4TSIs6jsLQcTbT
b4VUi8RU6OFyTaezsR6MhBiv1JwWGnJccH8UsLI19+DmsBNN4g05oDBoNZef4kDx
xUHvx8bM3IT84MbBSCFSYSAB2Ptca22le1LqXrpGvieXvTwx0Zeh2lndcK+xWni6
nIgITyfeRzKcHvXjPB2+oPuQgbgS5rVC7QFG2h/AEG2YFfFoKAoa3DdxukrLTwsJ
Ccfaoz9g3qWpEGrtXUwTFe5Vp4XVpQ63oUK1Ei4FHbqimeakpcz7a3hyOWpqWBU3
e9Yo1uJEk1YtGvduQwn4zSWK7kEng/ouuWEa8d80pkIoReQDWiZJQ6REXP2ykzDf
nok0rhwflqOvtiNXvj2JZs0ucq2JmGBeYYD5NHcq12BpGWiMU/mZ3vPuAaWbBoCB
KGN19Q9uvz76s3xGEG9OP44BSRSg2wflJRy4ufdlx5PtiPmoNesglhezads1pRmp
ah7Zvs/BpOhdoTxJ/IA3+M+zL/ATKroA9pGDlGw7JNb477ljKExKucwnEwV+Ct80
mMZpvp9NRhtg4W/D031VHhMk8Bs9aTlxKvaJRkeQSgRUXQcUqOjU1ZoDNDGLuhCA
G6oVCKFjxw7AhcGV1kkI4CAsEUcpsOeSt1issGzu1ObvLHvwtb7bVy6zt2/1vYVg
e20W1TBKoWmVDV8m3yI1Ci0O5qaRainzzFjxNtVPNcGtONhQJM8nSsMNpn3s/jnH
0JqdxF1gATRG6KiVPKkt5voIeMr8EUI9GtcKYEQvI+kQK+GcWLre5q4ac75uaVoU
8YVxyWXGTAVfthU7QA4GM2GHJla74RgyaLwjDJOCw8AbQr6lUEpPsKfShgO58N5r
mDxXWRqXPo9SlX+zUHm9U82lrvgG28cxIasMOKK6NeL2a6fxTcJDgdeQP0mNOxhk
lgKs+2ElwA0n3Mxd9R42miVnNIycpTveO1t5tZEC988LVAhZ0NIOIh7K1EQ5nI7/
/zjC9304W380IbEpojgYkq8Lcs2Lwp0ItctT7eYXji8hEp9TOcHdg8OloTJH7IaL
3mud7j5CqPgINcv4N+CtABV7e0Y+kD57fnHdF8bAiO18WbVe1Ab2PST5F0Z/TqTC
YxxmY9VERfwY1IjaIhGC7e6+fcyVPT3gT/7SYiQnCKgQuF0zRCUe2hwSzEzQNz5l
Ag79NmvlyEHu3WzKaS+fLNd4MDNLCCmsRHUYNYysEkJAUtrxlSiHnRFTlsIKdq2b
MJgPuDBkrntP/UuljhbbswSsoQsCe5f/N451uibVMQyp2Jt0TMTdq6mpj+duRDKd
ZRpYaJoJ/9QztLyJtXIdYuaMt3iOR1vF+mPcxo1nb+0=
`protect END_PROTECTED

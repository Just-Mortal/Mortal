`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqIbilnHbu53sQB6LFUqOBG80Khp4zTx6AmVogoSImpjHdmq4id/lWzbewHm9w1M
TV1angj5nMitV5JideCVovpCyCo204tW1leT2WomivBK4dA35VO1v0Ez8wXB+e3k
uSTJQ3DfRbWu7HGHUBpV/jF7ii4/Xtnxccflf9ZBTACTAkQcOI9u9vCWjJTAF/6v
8DnIkKJ4Rco12vrvvpkCG3X9REOtqlen4LumMBgILBfIImRTtFQ/ehH1fIyBzCCX
pMlKO+pwM/cAqwGnlole0iAZeLQWaj3E0maqEE90jfYiidHOcqJ6t4FU6/cEUsHS
loBeUM21sp0iIEt0T6QM+xm86sfVXNwnoY7dD2CMmcluDzDR6UI2AQuGYMThhUYk
Gf1cRR0Dll+tFh3dSX7xop5Dpg9yxG5YTN5JNAUGSnh5iid9OkY6+M+WntNrjQjP
SM9joQ0aic/cYBqX4GDxwra55FzDdPX/9WVqrc8RniMMLLI3zFogHcF3mOKk0vOo
fV2y8ZxRnvqpL2kmzgUAFeumo6fpxEqk/XTYRouM66i8ztbd+vLOOEcf+z5XZBrD
LRrDWcO2BzlOhChON8FIC09UruY10B5ofP3sRW8iJzYhgqiRwhelN4tzC0jBhddX
fi2F/z6rSVwmeaqeptVTObVBLqf86aJnVkmXtK0TryB63XZxtKGS3M2GHu3cAwIt
Xf5sQJZP3jPuZe6SxW1x7zE9yxUmx2YujKcLaeeeY4T1ZZ4iQwL2+06mm/kv9mnE
jAzC7gjY7zLPHsyvNE5njA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WT6+0SAVuaCoK3pFiU8DX8sr7wpN0BMqwBYaYnm/4ARI0kSmpqdPUmQeVgDLBgZp
u2lzJsNI1fCkW/VFm7xEh1NS2IVi634fWlEWXMJsoFlj4P/nSMjdBst/lewPSj9c
twpEJ83x+aBR7Q6+7299DtVN/mvWbIEYOSkkWdBYZX8PARbcasjL+6IrVxdtpp/C
L6hUA3kErdWOMBKrCqH7E7c1gCQq54121xAc4b7BldLJ3EWpZqPeEHhQrp3kSPQJ
aNKqmbYFZKKgFJDVHclho+gZXC3CX8jE0TwUDpXEXSA6LykYCYKTawLIbkfKqhsh
Kr0hLA4o/uO6fij/6Wt87YIgxEuFjRqEwXUFPY+rIBMHu4Hq7ZTd+uamxkYzaZjm
CLDiAstzNw3qVqk5QiVjRBg6NYbE3wISzZFnm8xAInJ7ol9W4Hf5w/knmMaJIPLQ
y3JmSESDVN0mhn6NDFPHLfQAuB42RYmmTBGCTtGR1D+nnNrNWW9sMK3wb0z+WhhN
fZaBhHjC/tsNMpAZGcTW+RJZwgNzwNznTmLFnYH2nK4nUQGELD6BkH+zWoFmFxXd
RH6XQ3TyB7674ngRQTHtciC2+Fy6R9YcDkutFhCKcPnWpfcvjF0FY7k5ujJLN4Hj
/NhI43b1/mGqtkw4WeE4kY3anPsfdMrf/On18GoZcARGKybgF1h/3STUPSz2yVWs
hID2vfmm/JJKLEuBRihVwBJtRbrAPImlZfynR2Qmm6kz2ksfG1A6r6llSdYmm2ZG
lf941kzLox+MrgG0HhIQlq3I//+WD3OZhz5s0C1b1NKL18NFD9qBGLZZbN4L8U6D
S+QXIU+Jf9xxPQFUHzecx2bzi12JVzfiqjFFdbQ0o2tNIrBl68vu+5iSm3V4UrPB
pDyEY+yx4RJ8lwsEVikk8Rx/VLQ/1lvSSdC0Y0Wm+6Q=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uey2Wyb4RAEE3DW/DSxAydTqr/Uxh+fVnn5Z2mAY68eEfjiOgpx+6h+GX7UtWD5v
etg3Exp6c5DWNJUFsFWeLw2BkUjVGrnTwdd1EEU344gqdRfkA+xcs7YzIVQFPl88
8Bi/CjR0uUdqh5Ag37Sc29Uq8QNCG7zU+UCYfr5BLOsTUf068MQO2f/3W8dQhOGD
aCXGxzMczpOTl8mghyr/Te4Yvt5ajiMm+QeBTmAKrOG76T3BPKSFTJDpLTVDKzcJ
8vrMsJE5OsmHkF2HunZgb7gONGynGRg9YCwUNsSF4hauZmffhLaOFmFinbaaN1hB
188uIesSAaNFHmYZaeWSrxDv55cWThPQMPp94/HsaCYsAsrozCAWFQq7EtMnUdTU
yE7tTgPp/qPXPDhzyVvibVI/fCsdHvLh45N67r9SXiL/oSy5s7knz079HSdm2y4k
lmWiWGGrU83jJ4IxuD0Er2iFG7wcOTcawQDS0MI019yZW/cK7BLHcFXpNcjeW9CT
IClg7EUB+clXmLTQ0aquRxlW1KjjzARnq4TE0ST+4NQpXNdxO3A9l0RyLdA5kxmB
84246kL9qeM6jF8l1CQweOBx0YVqepPv6smJTh4U6BxTL+SSNbElG/cCny6BaODB
+4mPU4lpopzqi5XhNahjsQ==
`protect END_PROTECTED

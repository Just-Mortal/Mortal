`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tYKbqx4DsvC6FLW8ubebwixUfgDCZdvPH+DgyEtM+M9PPLetiZWDGle2M/2FYXmn
z/t+M1FoLdpXbBXM7TUUno2kLtvh7MnUKJkFzcECRtzwpt623DbR09dPwuL8d50a
AjwNvietZdnDAujbOXNap9V6Dv45Gp/0sow8LJ/a5o/+yMaL5UkUaozduc0h3TZQ
/vcHH/TLMPfoXtPJ+65eymdBT/jF85mmmaCZ5lYDSHoo9HmAPlAZ/H/dMz7UuBeg
VgcyaVvBIC/lyW/HglH4SAlwoK3ZigpgmOsWN6HkqroJTfp2LHXCsqK2tNEcN/eC
5Is1L31jkY1rpxeojxx70ZGFhjxnTFrpCEkWwNVwVvrdd+p8ZYicycC9rlIibgqV
x2SLgmWpa90AKbvRa68ufCumVTx/5KHqw40fqm0Gp/SkLww7D9G3FXN08BWcCOcb
S46dJJUMv2I1Tfw0SErcWNxuIOlImm/ZWT4r/Hrv4j+/qV9miEmqa7ZQyVKiQ0Gq
0pWBzF8zGk5/jl9qj/pwA/UpYIgvDddhQMZP4Pi8bNJd2M0iVcrrHw5TVHwJOno+
zDUU0MA0pBi64KwAH8vlsZdqbveoEbWbWrUJA8V2JFT8XaZLewTkAyL/DvoaQWJ2
mIFl3e0A4HxePDdmhVTc3Klj6XAi883ojL+oJoYpCU4DIh/GjUq6Cp8ceuno8Zfp
MhgPqx1Y1O6Bamh3SIusp0sJBrrH8rd9G9x6+15F2wLwlkabWcAM/xC8PCqL0EOd
LC5twCaYhr1DOpYOczdi4prOGnEx4qdH0eaxsAs3wT84twE1zcK4pC8UtHBOnWUm
dL5EguW4S5N7VFac8ZIl08IcPCz6tfwCqQTKtO8x8cRHoPsVxOVhMZ2kOdEa04Hv
8oyYD756R1MyDEiRvMT9EvRtcrel+BL7Ki+Aouwtgz1rTxyC/6ou1i5PICJiFe29
hoDLCi2wDnvWrxIRqwtAGipS8ueAqgNu/6oguob5gKIoriwjvrg8KTgRmAp0N+EA
lbf2n7zoK5MJm90gVtL10lq5HUsh+gtjvrE9sWUEsM5QcYREt7LafH14iTl87AEQ
geoXT+RTfIeV6HzhCgCJXD/2NsFJ+FFLPfNsveaoVQGizHxPo3dfp+HxuLFNd1YO
ZdeD8nT9mAo/DwwPZ8T3gU9UDx1NhyI99pngNv/kpMng1ZmaNku0L3SmIDeNxupv
YvFMB34isslLi4muSa/6NSS3KLV+YlAUwpQF5zxa0StOOcQZnx1WrCje4416442F
mrLHmm/EqUCbSfGEheYAEcNn+yl2pehcMlHkqDcvS+UEwggrmMzcCqRxtr10Mrk/
571CEugsNmQIuvYgIuztGcbR51AJdMdY/M1aAtRl1c8Dfe8eVNnbFH1P/SekBXO2
l7pIvThXJBuo3PhQLwZgb9ZKDUJ2eQAiY5yG0EEz5MxBYEFhfaI6kOCciYyaf3yC
+GvsMoHzUNYHCJj6rhtW/pIHIIduJJYJAmgyvetWfKMoIwgrbTIegDnMxuAK38gU
Hb/QIHCMDQp934tKAukIPpSX/iyqLBCubV2vP7MvM5HKbebM8K8Uy4g6bVbvFBu2
HTq7tGeOgVcKNud3hiprzO2Q1tWnvyWsjh1mCUTFtvpIC/J8syg0oS1IsW6KBdlp
UEmGW0mu/fYCPuAE+ehtRPL9RGasE8BN31W5hCObQEY0MHBdHkJsfNuiLfWiit+j
H7whQH3/To/9eFVQjxPitxu+ganvk+Wli/ZDNgFjHejrtzbISi2cqlGFDBMlKH7I
zQ0Wj0Vp03qa6Fb65kSSPxYatHWiqKx1+CzbuRTJxU4WuCUh/WcIatWnbmx+xpbu
FOT1V4Eq5vHqG26UaskuzhpYj/MBsJoQrJXjmZ7N9AlR+Pd9P7QbX/3WE5b0yA5+
PndPOd+qNVqinKps9ncYvfuC1X1wuHrfjuTUKHJBl+QT5ku0CK+3XP9DwHHWzTPt
LqSdr/+YYa7K1d+VPuyXj1QcDJz+Ict6eMKl4OK2XWyWSKJZ9naCRPl7xkepGn5Z
YUwwpyUlIWkv2ZiVmzws5Ze+ijY3jwzUOLEysIn+JqftF5XDDbHuczgsA0qBYiBJ
ODWIsyu+3omd7yf0mO1V+H8ZN5BuY2u2aGBWpWxZ/sG87iqBbB7FWJZSBadxzXsl
ZS1hNALACbG5mvkfTlHZlqKXgAxfitCzrYgPWJFiR2TB040P6xXBxJ/3stEszDMf
23/8cFxxupNpjovSuRWDpER5HNJUh8OdPA1SbZ1Kywib4AUdlQB3lNRe8ae5n8R4
k8AZ6DLyEXwWP7aWqX0uvBuvEK2BHdEUnF4aZEwq9SZ4trfeCM4nm0DWWllncyxS
uPzs5nG6iQ0ZG6wtJDzMMuIYugNQHUPIe65X4YjBwelW+Maxo9nvWtcz7mIwvuE2
IqECRfswuhNpZSr8gkid1o/ROBS1jukkoLd0H0S/3ZwXnaThBosgB0s+QSxQhtZx
6TUOi5O+lo5A1yEDhnhb+aOzVNUTJxJ1CByxzRlfbvvSmEqTLZ5Htxf/xv9OpcOk
8eoA8Ag+93c8JvfztIiDE8JKgM0OE9ass33cD+KyG0OXCN10GaXKawZt0EWqBMM+
TSEXXtMQ1RJh5VQIEL25aTY7QUULgDBFzr39LRqwajo=
`protect END_PROTECTED

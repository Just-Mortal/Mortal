`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xxiupaQC5CkEDeDnypCG+fx5AIojd0w6/3zHDSt/vC6xyaCXhGRzY4CAderqHtdq
nODAMhhP/qA03n5J35JlZiFkeeSmSiK7/YFBdKOlUnVei4yQSIrNUoUALvbCdL71
Oj9sJe6OhyAqy53FxqVMjh9pEWl5k4HjAkFfDvfDj9Q9kmT06bX02TFacRTJqW9F
7aMqq37uhO7hAqN6Z9JyTvI20QC6TMd1u5Q9qRBC7wmK0ZrjeJOT5cjwb4KjF4eE
Pvxxm1+2TCPZGOTqG0Ez7rGU4BGeGiEqwDPScLF+mNR1Ep5i4zyAcePoaPAoNXju
ToBgBKiH9FmgbUSxWSvvxgPcl8T4Ma+/9j2mdV9nTtvyiUKSGtq6HAaMFaZs+uIj
aSBOwhdfYQJQh0a+mnQxrK7M0KG8aAv42Ue1jTa3fqHyGlX3e4d+BPiOqieVvhpd
cjSj80Vn0QtUhnAOQsHc0zepO5rbJBDdcO7bfcQrKNIreLUb4coJSmyDvICmhZoy
4y2JB/Sm8/mGZu/S/nWvQ94ta7uji33VU7k4dunkqw4k/vR7yrNyZXVc4NRVb6nT
DrrPo1XXXftT8gb5OMfhS5uRXBs4OiCony7maTcZWBi+6dGJ2vVR3Wk1wK/Tvcoy
5Sup8xav1/WBDZRZ+mYYw3p+MM5+CmSoU+PsqLfJEub6maGPONd0/g+7hCGTgG+m
QCHB8+BrMw3bCghYCwLDpRkHK+uCfqms97AMvVzz5DMDTcDqb/lVGPCwxZ0PA6lL
QUMBDH0dvOCHg4UqDRMKNvVXc2u20aTbk5gHyaFLgWft1rtMRS8GDzbF/2/nH+G+
dMrf9bpNu3xtfA7YDaocx5TOqLPOS+m4XLjqJYcA0/9JY7hR4eFGx36KRMhnsUD1
jsEfSbPtRjPxljg8HyXRw++tlxbciiD481oXnQTkDRp4oSqOsXmIpC0Q2onEgSoM
umaCfBnnWe7ew6SNiKcmbtqVX8W8mVxLX9+MecJaQ8NFAw3OkBbx740/wI6s5gBE
8XEzn3S2eEmXLNpHjff7YdQYGLcJ5pfCI3rBU4+9cH++mQsMvuB+ppa1ExZPidlp
Gitx+cjA2IQz/GhzkYWf9noQbipEIdDfHVJojCpE5xdAzJLH9oo9U+v/6dzcWIUj
waUI21XhwQXp9jFgEmcbFkLHz/XsyAfcLHzExEo5d7/SgJcDgl7tRsqxjymq4W72
KSebI/lZKMK1SSHxfqviRwRXcVcAnJoykLBWNSdqryHt7Dd4OHh59JI72pGmQFbQ
9Y7DgS2GxW5MXvJ6KuvN892lnkQLv/Iw0akI6kkOk/7d7J+V/De1V/Tj9rcKakxQ
DWI8abhKESJiTVT/Jq1ZLhiRVYVSMvD0JJ+Pki6OXtRfiJDK4dUonFhTb/zV1Oe1
3jXDksVGaoK51X3Zm9IFDNLFf3ec+zRSSvmui7uUyPZC5ETuJjVGHtUa7MpbEO1X
DVJMsOllkCfjqtk8IPFrjpbDTV+6gPj4qZIMTdvMgBFd6+NpRILfLz5SvbcnIjJ/
Zp6pN2xYiKHgNXlbyNgdZkg6WgVxDfFzDgZVFkJFvAFuxkMVVi8NpCOag1L+LHuJ
YnWKSKHs+Q5DYeoP7avnXJOgcXu5w4lGKvDyVMb209PivNmvjANl45Bvw4AXF3SG
S4AFV3AItvdiekSJbAmso7SJctNbZNGA0w+QJ2s+IgrSCOMjK5MF9gt6fLcRNTWp
lAKhtcvE4wyas5SylfJAz5ppS/Iug8Lntj8M9XjiDFrVDOF4rP2Q2bCLM91LDTL9
MR6NkEXeqx6kBBg+4kFN3YnhGguEbikYcOOdGpVRnP7dUqPmD/d5F0GIxQpynoYT
NXRK51XdCYsLIlwm/R43Z/RWjze0Nr2mBGHhQo4cxn25QW9zxW4lpXdpAht1OIPX
M4fC++/PemersBJUlPnf91Bba5/CVHgsWu+FLurII+MQe80ANgK0ptL+q8o4KEH7
eRRpc7+UstsUwnTrgK8sCCO7FOhJ2nXijbXD6pJy/Gany7pt67Mbn+a0bk223K8v
wNDo8+A9TPIXy/IPrt6MslLv+4VzgzCosDfbMb0AQypC87k1NDhPDMn+oiD2KdrH
QbUksuOEQEEw39twfOwX94i6WK2INauFm8TzFDEForb0tkqt2k6B1Hk6d9EC7/aF
qEj/zXUXS3NbuoNdQojn11g8zjPTqPw1YqJPqtAsUdmQxvxtClopJzRkhjGNXHyz
RGcUv765aMLtEZYJdruJSpMgJolzL9oDszoa63ThFJR+vD2uj/wEgmqAVV/aybxU
2wlLWxjjyahfm5Wq4EnZgZQMjb/zVTi93rGDKWnB8EghLwWc7xmRJy8nA0s1hCxy
hYLeXTb/1vqal7ev6kUeXhkkWkLG7gw5y8/Uq1XY0zOEW6yXMBd/X0Z/KdW1IIx+
B++EAqWqLzpv9frzINYmjIkt+O2idT88AQF+AApsgVHnxM6rdK4sVQ/XLFfROrnn
3IlSTFSFcTbifJJ6AowTLxyqADtLQibTKPoY+f/7S+4VorBOuFm4USSQpqiw4uxD
wMesSIS5Rg6kjQEh9kdm+IDanMe9uhlM/ZfI7FxPVrz/tZoK0N7yINAfbZ6Z29aG
pgdcGOtnEwQ1TAtx0uHv7YkZWJIMbNni9tYgDtIChDnYuyeZhOtqunTBrKYS0pjU
KLGz01RYcJcKfLNJ4XoaNGFeiOHZNvViCLk5+7ZhzsHGTnAjiqbiGe4x4EnLjGId
YbFgrfZiwdn8Nn1NGp/VSkg7xYOvUqfKgGrOvGSv6UI0biG19rXmMsa+2+ou9zk4
zLFR5P0u/NJpJYpw58iw2hiDXZS3y0nW4qSf2dl5Rc9O7bbBNHSWhaox3kdTwcJ6
6RymlL7gfC76rlf1f+z7YYALxffQ++gpACRI6bat8EuR+eCm/W7ESHLs6P1Iec0e
j2fJxM4+4EeUydnYIM2GYwh9iXjZP5hL8KNyFYE9nEOoFpF9cer7397JifWnPfdq
i7JkfhCohxpvAg9AuNeWv+KUT9hqIMwApdHpLvjOEPtQuvxdj/6SI8JbBAT3eWQH
uIS/rHB85uBwBWdYDpszu8CwzeMNAaMMgMzPjBv/CXAG1znMIfQ2To+6HuEcSdzR
IqnzEp57jeDHo5XckP6mf61Pj80cgGoLvcLxtU6jqxCMDekA/PFmndSpy0xsRdg2
k1Sg5og2ybNIF0EPfJqZYQlW+eGuO4NJ3t45MPzELBCgvZcBtD5GV2pk4rQES2Y7
ypJ7yFxRy7dpqDcAngBeZtY1OiQ9LnDFh5dQJ7/INHP74e6lfduQ4u+4kCvlGi7B
+a2GRUMMjftNTqJCbG5PaXvmLH6ZcIUSx4SIhTbf9rNhSq8cJ8OkqncRmrpQ0j6O
3hcT6r/cnVMyR3Qg6LGOT22aU9pdBZ38QgollQJ9nf0cf8wZ0+CM+B7Ipy+NGFj1
6heYk99idyllhpD9S4HvSN7n+0ZHmo9HzPlAv2tzbQmmFLaY9ezNpUa2IRnryI3W
2/JB8Hz9zFXlOqOUo/Q2jmHs7FiSducrnO2EVIUq6QSxQs6QpAYVeLYhEwnR/B/1
hKegocUQDp2q1xbzODJd2N2yTshyRtF8CvFPhquOsukxLUfo6JdrKN4BdhdvbL0b
KiWXlK2RFMkyfIvdQmY1qKV5OQ9qw4CwWBPP27MVmNJQ+bK2E0Dyw/syHgoKtpkO
pPADYQF6bq2672SqRKKFQfLS7qaBF6J4fYCEbsnpS4rZSMqvcwn5d0e7z0Qzdmz8
d/ZWUjoq9DakO1BqVIGpuh45Mp+BnPzhLRKafcSd1VZcAc1tNPKNgrr2lyj84T5r
Steypab+1rPtrg7QWFsn9hbrsuiCHn/9E/A4YVCwSc+JxHCDwfZntQo6Z7peO4J1
Qyw++9nX+oK5+uCjrSyiVaUde7LYlX+wFTac2qiShgPcHpYE/labbv2JXSJUVK9P
f15u0P/07GlZljMhN4hLblSmZwtDBNRiTzWFeO0ZOr1DteOmcLAjX7GfMywhIxMx
8wZgZZNm+nF6Uv6IKRWgWWDOgM2pdu3kL8RQ6eYJ6CgC5OHnvvottj4I28Je2wel
fpGDMvtfvl7YkkzcW0jP9FPUix1VrxmXW3bRXP89MJgrayGgPvVG+F81o3IpWFrP
lxd3v8PfCLZCyeW6YuC7da8M/1QFrDqLowx1nE1Q3rWVw+oS9KNhvKMYYJs5oirZ
Nd4ZwzNgz7yQgZozOmiOUoJFfmaG9M3BBWxeJ1OkJiMsdm0vB1A3CXHO1GxDwrRi
se+6zmnp5lrkHoZP75+vx023CDUi5JxTjLjYTmOSTm0+OADK0nnbHtXGH85/DTbY
ZRtAsZX+ym18xTba75mJe6JTY+8vMs0rlCJ9XD5PbBsadwm1zezi5Q7oeWnPZW2U
z9Y4aSddJBIBP6iGh/loV4EfkC3oyo5ezJeivm32Gw9NbY4lSrCWeVAEVEfeYCkr
nwLhS0v2MAd0tIGizk/moBUvzq5Rjzh4zsHGmQ8m2drvZ48VYzph0shWWogaBPqM
TyJpZ1yIhjgQOr6irxlV0E1yvDg6I90WNHOvjwxLUyCGNsB3YnzMWmc5fu083Ovl
MP80ohLeaE2tWRJbZO7g3LkBz+LTp3PqyAeZP3kjp1+L5UvEMFYUCHxuT2gOSWXd
82250c8X6lmhbnHn+GYIXrXR0h+//wZgVjxqrdXNOWH3Ys+MzJR40k+O8MHNR9e4
5xDBHOEyQV/+d4qFR9IzA8tgyFTmJyiCDHmDp7DMOj/JheuUV0encQ15sNWhdS93
Xakv8yynpSI0tIKpoBYofcRap0L8S9gMWnUFVD5HeWHhB2FkKS3E+xftg/pJv+Md
Ez4pM8kFYTxHOnVHeIAXZvMRoau69aCmr1lVJ+SsSRq6jBtl3hYHJT7+3mIfWkDL
JETEiJdsABsp3LZmY0I1vKGpjlaVx51ZscmHC7xcIoaD6CNUsTtk6xWOmVB/V1sp
YH7kiaJH5Y7Hizhj4hLVaqzCiwzq31w8w/vMagkBeIJzWK+uKpXwZ69yveAp6a9u
l1hqmjK8W6X0N7T1hxEHIfO5u2mosYd15C20IvanCt7/ADW8TcdmxOtnjQa3Uk+O
7wgVhDDLkMJbwUIZ6zHlLzSTapotVCmjp8fILyj/9QPsteuzqy89NEkYiQ/1k0ir
XdvT9bNS5ijW+QqHGX6LxZ4PMVFQk7HWqQcxUERxMgPheDhZQye39bJgPHcaZ9E6
6RU181JPKKKcF9dE4ErwNJSsbKUDlwQPN/BOvmvWOMU7s/QgVVlrodZ6w7GGy5ll
jzEcyFpTr0mnj2+jEhwuUjym6v/RDaQQInt/jxjDA4EIfNmkejS5sH/E3mWeuUvH
G5IlZCeePzJ2jb1roXzvhRwfMRRTgB/C+eiOoDRuk7JCysQNWcMIXZmeG2z+rQ10
AJHc84N4Ueyj5ZJjL56n6weEQSAQd2S22kUeLbt6BwpiYOh3gyVCNUYU8tIpHHKe
Mnf1DTGTEmYW9MueJxrmHJR3ebH+gUalwhBgQOczW4/XTnT6JB17vjI0UWjGZc1l
Zgj96UWydLoYww0k0WhBBiR0kA6d7bY2h6NbUum1b4wq4AKJR8nB93Hr7JDfV3eQ
76o36tEIXZqdabvUhBwy0s1gro9iVfOdG1RmJI2frV1/JhcGuL+81T0niTITrOGo
H/bp3dndduWBx7xcbk1v5DF4Qdtv7WKUXdBYhbOoFQV+j1Fk2wr+oq+qPjJKTuZx
ImmO/WPvtVa8Yxxw5rEqg1SQSx/iGNH/F2Acr8Cif8yHFO07JwtKxv8KPn9f+B7J
sRuX8kdWEi0tzAe+G2UUOJE1/M0BPhju13wzBeGLP0Nt29ed8Za957Ckcy5oUDtq
J3jeVK8N7VdxyF0A7LlWOdPwEiYfUqOkW1Poo2pzmGjw8v1uDyHoWAsDv/dWo6SZ
DvBqGQ3JKkmZ6WBfBiekTWa+ug29/ruYbWBhFkiUyLPRBfFwO7Cj2r67rkLCooCN
IE2QzK5jkLLDLWreApkH4Uga/8yJsDMyqu3bgL14+hrKB3sTp3LkNKJe6BH/ISVw
1UDZrjkRoDD5G6L9ob2QmLhPPWuqV0vt2U8TdntUvqTdF3ecOZfiR90x4e5oPfWa
W+alAZZ9qNo0Esdvw9hXJdzEL0kmcbQK9CujesTG/SRaM+jJbVC43hCAZzTwZ+zN
KKKdYJidpedqgFncPxyACKAeTQg+b5ppCMiCUifaxBydD7SACmBlqyK2TNmHfTyc
Wf52mY1Fky52F3V9l+cJ+2oU5SOWXa09/m7aMOQcuK+7ohctY8kPirzjoagePuKd
BStWn2INAZFi8gfjzERJ/czwm6k9CEl3cbOKrEPFBzp6O+CcGVZecazcssBArjIK
4aHmdQq7TNjpc0OoWGpWzdmbEDLkKEMpToGJUnhhcIpv6FyJ2M86CMd8QMEii9UM
CfBZpHtXrbOJVWHJspkNCYMJP97n5KYYcvK01ZOlXTodHIzFQzA665jxwBJWoeul
PXmDV7zF+MIO3qfLEwZZewxLG4dyoLeG1X/e49OP697h73ArEQffR5JJAnBOddWh
byiDEQPoR6CxjmjZx5soGBvd/UXpHgy8W5Ftk1vyLoRXE3tNv5xTS/5AQcPXhAia
tJZxNHl0WOkaKhIhBN4MekzxWAopI3alVQDcPPmSVWX/Md8DRinrHFCSG9VZ3UXC
fNLyTXp5Aa0Z1k0Q5I2X5O9oXSiiPZ4UMawYfU2Vy6jvnS8v90+F60rZ/bzl1Swy
t0bsXYj1+KFIaIYpT63PgRJ+qqPZQ2GtXQuTaz5USvHt87MznaDJ0uI1d2oUyDIs
gCFDA45aFUZsi0HGh3J1blqW51ttCDOsw/Fvs6wTFTuNTWDzWI79tRcgq1cQDiJr
Fdremi2PiDVncSbEEEvvvSdkfH3j27TR9IB7xDx7aXOAnYv68qNnFbR1hf4XSfZx
y+CD0An1YmuphiZou5hs/vg0U0WHNqLjS+0KTb4JZ6Eps5X4DumeZSZzXhjeve5C
x5ABebIqPxa3n7R+iubFxCPXnhKlr9GA8WqkkmpgqE0wRT1FnTtpeJn39W1AkO6G
FXTuRL0MmiYvHXeQYW+E2m7SNj4egWc+NOV5fvuwbFNcPqcmjZVBHedeloxiIfZu
vzSS5VL0BJUqo+5u+YX5bux64V1dzv6tZK7ApBa6hD1fGXSV3jjJj4BW+FyE4gLU
sTi8lKVNyG6zhQDdYlMw7qsEd9HgOWxU3QtnADaoUvxerhTKtSqxDJQU2BoeYH6S
Xcp6GY/A55LW3FoT8DEulLBMNOIde+SiATi0kTcnUmRhyLIHt0jQ1I2JzD75V6L1
eEdeVbQsVcJSQFhgzgyg5FqYsMv6sVOE4UjWuOTgLbciyVlC2KcAH2IyuTqXU0FN
856hxcBJEStD0H9MWMFV1ka8trdSUvhscjKzNyxAIZPD/H5CLQ79oTC3Z4VFmSRT
lyAEZQ932XLOYFN6BF50LSUnxwp+yxLE03UDoyvMmDiQj7OML8V9AcI5x+EEx7bW
2v7KwFCJ9ZZ0+T9bLtDC60D//g+LO01fM1jpdcohPJudCXOSVMxiMCDA8n1coe6P
5oMstg2IPX5dgZqwaMUrCYM/19oeuBebk0f7l2OWVrIzlCuRyhk+6hBLOXkpFZu0
mRniph9U4Lo2YxUQgMh/4RMmTXqLGyhn4UxFqY4k267VDAStchOvQweeQf3/WWFu
QjlEpkc3utrcWVYSZQEa3UAj0Jnk/QHJJFpVG5MYnU0IvV7fBgd3+VY8qBueumbI
MX1qP1n51XPk5XHftYB8RV76cOoqYuzV2+LXFI784vZX1ELq31zN0yGyU1OqW/VA
2eBLgDNMRs0wXemChyaDl8pXUuvAN+zsG/gBrSQpsSQHShSojJGQZceVVL2Ta/qG
vC9TlRwRoBIoWvH89cw5LfVFEjvEMclnyCihQ4DCfSsI5Jd9I7BLc9L8mTGi2A4o
vLjSPGNQM2Z8NZVlASJchIn7yhutR1eibNjh8/qoPtlvjV1BKNhuMyrB2MK6pL7u
P0lM7fe2tdIDVrgov2wLlk9sgiUYRHIZtEfPUsa/4jB4BE8ha1qpThCZsZPhgMgm
5hW18rgdzCYins16Q3xuPDQwj8GfVjW4O2+Bw0DJctX/0ZvLdFC3GJOzvk7SP2Le
KRycXiIknZEeFat/EEUeJdmZLuBUJKHrpP/hftcnJmrHwhEcW1dILfdNnXrfun9w
iae9wv2h0cUqOgikA9SoC2ZK5rUnz7Cr3vFIqpzeBvXjugstVi3W24VZB1+8090o
VxQvTXu72XLGuHog/HpteTxDBaKpMtoSBR/Vma5xnuVgQfnvwr4dD98cch7dltbE
wDhXR0Tsbuq93ApQoNcBKHWOiJcTJtn6jAYJjOdC4BWOrzS31YdnPDGpijlj2oFi
xG0ankSR3+yfblYyxjJcxUqeOZoGRx6GSV+6EwnBvbg6eQ7pE5dX0IGW7xWKWQl8
IMGiRMBDVRSndORxd0qLsNip41IalCtJzSkmRNbJJS2IQFbH+lzYLazbOWCXbn48
KFyj9KcLv77x6/Yqkb7f4l/mYDUyGssed3JCBaegtAEDLZmCRebGQKm+FGndFylC
ZdHY45wXtMTpcoMpiK5XtdfCznqWNdOJMoXHdfEd+XCEP6jZ6sVXmE5GC9da7glr
yfG1Y4y6HIScn0v9NzYsdykLM9v4KpmLkqRP76qPktBSIiRNgJMD2AJOnIlvSl4u
3PhSK5sqNXiloT5BVCD9sM7SGgkzYHgBnJiTCkgmP7XsQ9IbjD4QW60dhmWedRoK
a5CZUebVjdL34e13Fco52z7oosoBI/zyM2m1pq1kqkmYcHDQHJF2p6OlfgJyB2XK
b+opZVLoi6BcXW/4PiiuzhxJcLcyM7wzG5vsrC4hm/QyAace5pU6QiiBjzVniWoz
jc5FSdnFbsVA4pWRiCrVArux7plTYo2VPQ0+9mgxYHZGXBhwa9oZcC5pJHLfYiA8
xX+sq8g7spkvXWjlF4KevxnTHY9E3DPjRdNy16Uims+xfN2EsEFw6+Iq7aw5x2HT
Q8tzAsIYGyUSTrRYvvfbY1I6YAdoHY3YkHMqYmzsTkxF5sY8eX0I+43/kM4kGnQ+
iuwXcDUUakm4V/ZlJQrf2kMp2s2ApKGXrnYo0uBjLYQvT/mfu5BSt+xZTWsLwTvl
LaKBHlIkc8btFCTEsmLc0piZ3zKsG9d3zPX+g5b/BSasJLB7nvZ2M3Ar8dXnXadn
QyLXHsM1PBQFzXH+MHKQaLgTvFjVsG81GU+iLl3pjHd3nnEdBdqR7Mb3gVSrhJbT
nZeasMQphXe2fnN0dBD/AfAwr1VKDo0NDNmxcgRFkInu1y4oDsAhXku08p6RYjx4
L6Bh1fGRwgcRSd7/C0whCcDnOd/Z0Kbevyu36L6HudtoqIzH06DPXzRBdOPZIZ22
xVvM2PTOwFuRFwnJk0VBJujolrm0AoW1fS9dgRzAmGeUw+cySHRnaCJjDs6q0vhh
CzViXJm+Z9FY43CK/a4vknEgJ2SOSdNwaog26teTCwS9B7oLpWJVLeYfZMEjil9O
COc6MzT4hjyQQMaDGll3QUKmDFLtsjbbb7kyv1ZaDT1fvS96WN5AaaUlIG0O0ynb
EYbA4CD+7vaf89H27XCwhjFHTBiqWxDsDDqwgda6QE58s2lDb35T5M8sZBPLZNHX
esCZOjgYp2YaX/V+WkHA3y1eyMvkmrwyUP0cl1Hm9vZtqjFqtRGJzOHmVAGZVuwt
xuBTrwZ+uBweRge6q28MrY9rkN9DotvSkvd3vi6tDhI=
`protect END_PROTECTED

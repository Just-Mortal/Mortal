`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
grUsQjxJDvLTpNHMRfimdXrQt1n4FIRVTmtVxjJfgwV4rwBurMSi4+dFnaDBPcpU
lMcIm5P4UNZ/gWtIXihRscnuCYJvQGwruVCHKor7uS8KfgbpeocS+BVu2gW7SkjW
7IblQfZjBEkf6tWNTFu4sUJ2Rq4VCuNdqUus4S5f/E+gWn21QzvxZNFpo0csbTmV
uIPLARJ2zt26pP/warnRxCaTpX6r/5xlUOyFHwsxCNjF2+nwfNYVVPVxlEpIRowE
i/zIPpYw8TlcBsxUbM3XynAGCw0agOcfXE7uacShcOaQBc5/m+1iKkMNYdng2hYt
ePPGjBKGYLWdsyejGfDheSkoJvk1ctftfsbX3odp7Huu67RY0y5JKvqJoC7cK4da
XrXD7XKSIlBqG8szRlt0Ghv93g4rFjjV/tEo5PyPAQyG2vpqLQbvN6EGuuv7un9a
DW6/XlASR2aOiB7yuFRr9suQYpu1amddNE4elIUjm8LIMYIpYoT1E8WG9piGEw++
w/BAfuVuQU9BpQzCI8Z4j5LAndWirALGVFRkDNXQe5fe7+y4U2DvHlLcC9NEs504
AK2YnFdR2N88RyKvYj5b7shAQdnuy/vGKc8DgiMiBz1265Fa0ZqUT835wwi6Gxk7
lL5+Ak9pASur7MVhFy1XYCmMNAdAFtnZuaGlZc5dfJQJu51Feolz6EPJzzqKQbQK
nS+74NUXT/V2l2wBaRXtQ4CAYtOxQgAXBVZZriuWFFetZ6kRrYOEr+ArycHM6yQC
YcQTnXfkJky06c7L+OrfHbNPFTmu/0Fom8oTd1ot7KTuwaPyQTQr+wJKIv9CayLB
nQXi2ulNvalfL1uyNuL8qy7JAME9logx3ueQ6ZiftVeh6dl3jxLq88HgbS+1d/Li
n+TmMRU/E3tbNW2+eRN8OUa3/Eot0EwOZZMznyhlM9Uli68na0I2EKvt6bH4JCSy
d5sv5UPhRtK42veQQIBL3KGyrCWe+Vc5ZH9wC3LeDyplsp3DOaWdFRyiX23WDkuU
EQVRBHEM4x5At6T/G2NB/qFXhUosHC7QKHJaxySaKHEaOiUaXbtIiVjHUcsMo8bW
yqBUQLuPfchKOfYGdt1Las1h7vnTZnGT22wCrws0AXDHlG0rPDWNTXSztUp0OnI/
GioNolYDM3QGFsSiAD/UbZYLvkusoiSrOM4ineT9ckKVUZ6FwxrhOzJnd9PcL+ff
53biziBt02qTBSNWL1J2yn54Nt4rx4yapr/ESpx2w6URtAlNyaid4VJ+nx4DLJw+
OWgzcsPb9OoZnq8C2Er+ZgkP7HeO2IiWsstx812852QAoLE6GSeM5H4fu8LTUezM
Q+xcU1rDP5Ra6S+9SUWhwLOkUehR/tGKRZ1W3GTg3Dhs58TN1aPGFaVem+exvVFj
Aefdl5KPMl046UNVTd4GkMrCvWKB6zm/1V0usAnUTdRj1t//gK2A5AwJbiIZSyvD
Nz9Q/2UKVKV71cOIB5+K9vej0grH10julOu8HYvnBW6w/OskO0xGxJcLD6QjjqKg
/2jNZqXkOeyPz9mti07dxnVlpBGANy2LFNEsq/FIrmpSzrXIaaZlD1W6RR1EdjCT
QC+4MoYWl9ImHrIjuxs8ungEou7zNAMnqx8tjYGe5TuEG7/TVtWovJJeEG/+sK1L
8W3RU4nQ/DL4JK1Vw/ozl3KcCpR/MU5ngDNHZYZ3LNDb77HANC8FrBp5WrNCWr4X
ecDGgbU5p51ovqlMERFkJwUf4qUF8vkDt/4LxUeRkTDUWNjaV8RsfVpHdA45n5sI
NDHlevfRxGXlca0DTm6SSB7nCCvhvra+kKd/udPak0TG//BKNFgHwVD3JYNVanqH
nwKli7si6a4IocETcvh2KpEPTSa71O01ZWGRlphalPRoIKcrGP5PqrWECuVroFDQ
tGHo+I42alxwA4GBnYcGYKmB/rYbaTMqKvz/NzzjawCV/PCC7lqYn0fzaQLViPRB
l7UiaDpUC09BKyKsPrw5EwhPwusZtWzQsPiq+t1pPV+ezGMmNMrQdkO5lDNJjGOZ
qThGWW1VvWFPG2WfCeNiomNHF5fq+cjEOr4kCO9LZTJ3wqKRAkeiRF+6aNLeZf7n
4jNanXDQcovUZCHkXl63ogY/4SRevK+2GY+fvL97qRwekgg+gikxf1o7BNH8FB8U
YsBBdgTY5q5gSzAxGPj+q/O9AYC4pRAOhsvLJIdZ3ndHWF2cBH2YsdB16NfK8RvT
rg7/b6xOdO8C/8eRo+5Dhqqk5K5+Ja+KFKUCsXCst8zazVQMezZ6DhgApYS0AzwC
x0yFJngSTvNNoBecKCglvlm0uMq1D63Mnl6Eo/mpQlbYVtUmKTswkT/u1G2s3mN5
59rEWqlg++aD4h5Rmx6dtTFcTb+tcPehbwFaOLdtbgwSjk2Ko8BXuu9X8D7mfo/f
wyVOmY+b6P6+qTOeqw5frjJYPzBCOR2K00DlxD5cYLTzVYDsJ+vcWW46xdWNUleh
gUA52DMTeM1FDky18tAUdg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmGtpdNONnGnIQEbSCZZMHJb35EliV4qXKRUSNLtQ+pKboc/rgUd2FgjhPh+w9Hy
5KXIDxTB+qalzesHmw3cPTAAPy5PRAG/+O/B/Ez12TUMLXd2PHUUkIBka9vUbAvs
ox4z/s9+FSwMrcVSrsJoU7wEXNXSmqWff/J3PSeAPPNFM6eqKSdY0UhX8hG45kfX
Fb22FCh8/ntExdGKIvH2WkQps7bOZ0C2pvckqpTQn3bHlyvGUlpXtMAzZsbYIIVC
k61Fj6DuEdw488hfg2SHogXLKbrjRDLUarEDzN4s9mIVEif23+GdJc3o8Fd0xzmw
HjCVClZSRsdlyaasceVvA7ZEfQ7IyxJtoSl3BI/h7TFgdTqWp/r90t7uCo3G8elb
sdjg2P3SBI6CVwp80cyxwtmCS77Dl7r1hfk23WDpYj967iewsW8VdiAxalWyhgYr
GaBpqlEWIuokUS3gy+Yps8vWq1DpYqa4Se+Nbg2K1nowzCFvd76RahCmACtCLu4P
B0kY7YDS+xBr0pv9FfCayvnZwoieZDuI7ycXMAoH/GPLiLMzvYUMF0GnrXLmkO2Q
6U5YKZIl/I3D4gQbhSzCVO3lhouJFa7qZvMM4LGl4V4w5mbpdoAQ7d+4Bj3epQzr
z8SC7IqMmgeDNjEsfRUjtCZ4m6gL8cW2lYer3NRxiQqIsgJpiSw2HlwKPXp8iIG6
FwqDFLfQ/UIXVoE2PXugpb6TSD8ag04CzmcjOZOeis9+xW6IMl7cpdnz/DukMEu7
fFA5V0COQNh2c8ChNOy0rgPB8XDFae+YQjWvJcYdV4mDgcB8vwxtSuhc/SF1k4Kt
wFz4LIvA5/vg6HYhq+Z+6f08BOPfMc3cZyKyCe8K17s0MfRwPLeFsi/hrJrBiyvf
oCiri2JhgJrE3AewWKmm+BqkVXZOlLNTYHHDFkpLlwtYnGq6o2et7Gfsj14JodT2
CqCSNf4Ma3FDEkO2NMPON5evgH6LRPrK9QaNEWlUaNnH16RFW4TAJpEXITj5Vjh9
qjDimscNw12U2ss2mDulMoq6w+qtYCCuo5J7KsI6Ic49G2WwZHsuZ3B4oL5Ukwbu
0oIILURwm3DNkquxoiODfNKTASj8dIIdC+75euCPjqNW2Xq51RB1Sf3ORYQmFMg3
hbUl9a3fHflrIpJnk2hz/d35uMQSbazNlx1BUcK4gVMTopExKUgr1sjYffHojZKI
iKyUcFv2VHfyZRIpCfBFieP7Psuz67qdmZ6wyustgFB9D0dCUgdx7fAZpWKFV4bI
thJ77Q1AUxP9145edjJ2hN/KWI/MAhMa8VcgGsdo0F0iOhVdBiyukfiQXgDrAZUP
ChCdL6OzRwwZkZmAwd+xWB0sx3D22VM0hC++OsRPMmrQ7CtddeobV2JkgUFN95/o
rG93O8xB/VWvU3tb3s9NjtTV/Cp9+MffbfbN5TgPtA9OkMh1VPvNTZlPi+5MTHnq
JCQfwcMmt0WwDZH02ETR4t4AU46KFMMPEZwAIftKqp252C8ZFiWt3QVJ4TyTWA/Z
pC7i8mjuWOPk1G4NykFwD+PUf5HdlB+zUkGa1R2+l725MHUozqXXhbPhxVCH47JT
N6XypR3XH/oar9tsP7RUP58Z21fNs+/Xt6QCB46TYV6jM4QQxbzsrLfsboCuB16A
jCGFJdqs85wen86hzGny+wjFnqvYKUFUB8hlbjvunKxVv/hsgvAKlMeRslaFfJ2P
i7wc4Lb/sCPVsjEtUIO/pfjIG3tHBoXGIn2wtoL2TVjTddsM4Z3VkOy+Zj0gnXNo
DjPK7FIh5/PSSS8kRzdUujOxYEx3z9avYFC288rnKf8hL4JwLjLIPoQqdHQMtNCY
Gm9p7mPTLtI4DRKdMDmJOSHwNfuvyQPoVYOzMktCx9FP8c/mFUVjUzfCbrQ92BHI
+Ei7YbIoz+uMqo8ao8ndOyGC1/L1qQGqMUX4dxWqPH69bK77t4NthNpgg95HHCbL
bMl5x7y8PUyTbz7JWbVQNMYVWpNRQU0aqC+SR6LXg/vmraxFMItlxd2tzBn/hPjE
4vfBiYYLwI8U3jDJagQwpxD5+982t2ky/ymXjVxMs6sI4aLYX92EMJe8PDNdL53O
BNf748QALNHrBGZOEIsa9gJgu7ikPEpBqqUru1QvFL4IEqRXWTioq9MOIDNglHDz
riHgLeYbqUJdLWh4okM1qFbmMrTHFGvNOga8c3JTdmQlqA16h6bstLGfeVF1v3xb
AOF6gnlPZNja+rNwA5c1O0WAjPoUP3bv2ZWZr51bEXlQAK8pQEt4S8rmBZegccZZ
My4mgFjNMb+J6iczwSyyrk8O4Fa/BSJeXmJ6B36kB+pFz5bRXMIhjlRrBVI5xoGO
SYxPe22caHhcKw1A98FL1TahU9S5xIS+aG6Sn5A6wuO1PXZzXpaiZ+dBSjvopX64
mQtysKkYhaevWnbL4oU8XXBTUIqlUosrT479KnHOIg24g8GrF2zv3GYtlNvJ8B3U
iZI+i97fxWLLVK0iKgdqkqU2WoVEYVN1PmQHszym63Mz7HCe9hymfLRJ9Y0gKLH7
yYmufATJb28z/2HGuSk1GKq1KwiQpYWQ3Ek4HOSqTZoesadPXJeTWcCjMedK7MHM
UMQ98xSRz2C/nNLbMFa6kl4Doqva/xbdcFoPikKpUEVuG84M1LM/ccMg7cXW97lI
IhgsC57pzn3TzBGuXWEQSoVdaAcz+OnuldoIc85YHpZ2yhTn+M1VqHxb8D+QHF74
gi663leWi9XYUBPwQXXSrOnOlYDnwo3CvdaXXOz9UPfQkQoGlYSV7YA4y8PLGCnb
q9Ck42dLbqUTM3qqMRrzwpHfsNVhdTj/nE7wiLTe1geURgJa8so8NLegVT0YgEgC
FStyjCH+nwfd5xS+QFHBCl89b9X/xORvRzw7L+MkJQvhRRqUP9dsvkPyTZxi0g0k
J9wiLZqVLsQ1rT+VaLmo3Zmg834NKxLtgF9O8cVn67gVQ0VH19nFWXmbwvbSENXz
cjnrenJayar5Oo/p1fLptBzzg6+cdKNSpQkW9RG+BudNcbEihu/H9rFIjkxVBR2D
GISoD0HLd77dFemk8hztZ/8o6GKZJfSGvv3jGm0p1UemuQ5Mwzrt5wmHPFF7d5It
1O61Ncf10uJn1hm0Rh3DjBPvcpb70otK3w+tRhRnZzhW9zdsy6KOETj7DVBm97zU
Z/2XBhWthhjliYeOFCVtqJP8dO3hDanDcXuR/Ja8sH7O8fzHxVrxQu3eGAotULS9
CJNK3e2PPYLB5qZ24BjkG5iBzEIt48509T4H9dtq0JKmpMY7L8zQhB+uyeF+1d4Y
uTEmZDxxzNTZfQuAt2VX5ZKr4oGTQdsCPDexoMPU9iCspq3wBQiCoKB5Zc6RQvvn
XauXMPic5MGInL5Nf8enj+0txUZavN7/kBWV0Ajtc4+Mehv9ECboZCm0h1drbKT2
T+nIXi/F7wXibxQwYxPOduJaOqm/rLuHulG0JQl9tpfuO1wCzPU/pJYS4t/n/ys6
vgX1goMR9m3F909gzkZwd0T0kxbHhi+HfyGeRZCj/0ybf0ESAJdh1kkTAwVBty2Y
nZYvTXjYGm3cvsAjNUekuJFsywIyzy+mC3JadWTH/j8Bl+61vvqoDWSmO4byXA6T
qcL9DJ8tHvjdJTC4B234nZRyLQ1HpNwTPUaJVeSR2YWZpKvPh+cZueeSppjDEmaw
COJ2lXONQgsKJAXFlvyZ63nkDjM7SlYhHZhxFua15nOiU+GBP69QINYrtls+u7Kh
vYbFW8XvwtpThkuKiH7F9gLPn/aagY/LQT6rJGCXcCmV/f17NE6g25ZtXjVmFQZy
aPO+XP1gDltoxk0nn4bxcGA9n1sVziUp8HdS/wW1sUZo9X+2xY5LOqK4/rQsG8bn
V6leuUiuI97zu58lhVC78VZNy5YfFY2jWgn7OGE6cHLqUS8HJIJKiEfEC6ifViud
c4Ebyk9T7OOww8rbhyx5FCUbq6kmmcbMKMSiqhd1h+I95vXscE6zfh/QiD8pFF5b
r2RugM6Vixo92P4FG9B8oNvAwmQvRklzKGgPoYzExEVOGWWkSnhBxOB26tosja3j
6AK0np+ovQlPbZ0frN0Twd8G/OeqT/CWlAzmkCHbzMdu9cG4lLnelrt+/s0cgPjo
Ob9Pcc1qIbef9YzhDsnsgBgebwU/i+fmZFwNd1ibtYrC0j4PMsWpO6TXo881rIkr
dxf25L9/IgyDQHIW2+X2aKIZokWSQwZG5q4f+/JLNZMTxyrrxjt7asUF3DEmINfA
dFIacBNgu4yCCw+C2Yn7CVO/RVnKgO2DPdIEih1eWmmUf8YPnlwy0PXDFqOoHGLX
O5fDfgFGoWHCRfzjKyxyCQSHbEs5CrH8vKy8MjrY/buUG5Mc46XCmpAg0U/DK8y+
d5ymdPm1s9Hg+6R0XoxYBRJC0gYGwuhSpIVZkd1DQBPbqFgUrq54Jxl851xYz27E
pSDxy9Zo9SfYgjDAQpEPyS4KrbdH+te+1kB9xPgbCUwXm/x0Xt1M63kBDh9aDAzu
kJLFnDdQtGdDjXrKS+Od7HilnZoqbe4s2wCr9zIQO9OxKTdx09AZff7VFQsU6h2b
+oiwK6OfBaO03zNCwU9M/lXTVRyRANQs50hFBVZXFWiIsZ926SvZQpDlkYAEcJfZ
a/gy5pcTy5etc5if+NLhjEV41lTWhBVHzyw+B8PZkejqQzu2+POSh9xlG7HXmAYH
qZYZ7X3p48Db3TXtUchVk9iPSDFu4IJZy6GlYfgpg5wE53Eab/+NqifO6izXIbdn
DqalHXLvumovgMUNuAKnfPJfqi2kGfEPQfCG0GNcEpxOhwUvCH0g/VAE4gh5fCEf
OCgOdcDntcsSWgqQlrgBUVc0sasUKleDVILYZ51CW7dOcTzoLYUmE4PyxhtFdHkY
Yu7Sfvxvf6htVmRD0EhLJp1vpj4W1h88GajDvucro36XQJmpuoq2I6IxjkSQmMkK
0Pw0AbvT+s5ykLZlvIWN0LU40ikBj4wNuIcyHReyocAhzqslqUf59EGcucoQ+J+I
Ca/FE9CMkzLuXP3LM8439jyh/VOrjRuE8X7s9KY/S9QbwmGLe/sw5IefeKKKKlBc
LtzW7f3KZk5tHTVw4SQ8AaywVD9fy69Cmekn3E/vjI/FyjNA8jSGjA3/iLF9C5Ay
ka0ZYkkF28KWTgQAj79etj8TVWzzFyZDPMgCXV3KchEpf7QkcBM7+PTLwutqYqww
OkvaWEbVIHscKsnmyFMU/ylH4nrLdC5x2jSg3nQfTQdhIDscu/+PuXS+nmjlxQj0
V1U5+km/mENUKypXBz8MOGyh4mwn7gXc9GT4twuks/nBANb+cfHqKKPL8xOu/lQd
uZtmNop6aa6STa5plHCaPCa5parEzxOlvj7p4eM9jUAD4VCd7KlNEnbKwi+Odcmu
OvrhCQDFjrIugqdOZ4ag8RmA7OLl0v+ppw/URS+wkmrk3pUXADnWwvTwfehHDZgJ
RWcoUkPE89gevomc1LZ9krZ5E04FkgaFKU7TeDcZpjRivyj5Ty2FRMIm9iyK84ew
DXErwQD8I8BEKyUYR78aobXeALggkeX4l902WgfiDC41DA/OfMC7KxdR+TrFRYJG
qbPlCiijeDKSJiTy4h52eUGN5e7KLtKlAgdL1R04IR8TaCmBNC2PvxopVHeGNkGA
G38dqgnRvzVcV/SS9uzocPkpVnyqWsgz519RenYrGrSi5fPoHMFNkRLgO87YhU5W
Uas0ru5Z5YBYkANaR7PzGysOYaGv9TYMOduykJkt9CVDPocbH9JwBbwgtdO0ntsu
5hcMvcqxRH50IXbVnwikaXWKs4NlAHExDjviUhSz1tsJ8ywQAkDKDauqbxmJvJsM
WbRAyWc+q96JeoWivqbzTaSYR4NwxEPpXMkDzDjIQ5f347QYe7d914JVKLRCXlAi
CNzamiEnFO7lQqgtUxPxgO9Q4cB+Tz5z0tA90AN7gOEeEPxDC5RcbksfW2/zWzUw
eH+JwTGCv7rhmAurT52x5BhdRl6V4YEwTzhOD6FNOA2jMg7JFc3YwynsgwVf2uBO
c/w2dY1h9QPgtcwdDF+ir2Zqbv+DZalbPirgBHEgKDxLfcdaH0mE80P6dhg3H2lu
ArqZVb/VBOKNRJGBnz6rNVEh2+/lVWyDQSPjDjcQbPAcP+fnNz9vnmD84hPP2LxW
pPhfLfoPROvksyzdJE8NXeAD++kewTv2pxHmG5wQ00/iOpDGdOx5UFYIMiaDtEMX
KTq+gl/J9xCfwxI0mtxzhjgKbXqzHxxzn9lF3NBucOgTAqPB0N93FIZ/1aCyOV6K
gWCvwMVG7mzuzLqOVJMs+R5rBRgTLXB+8XmWKX2vAfQdtoqjrFBS75n9Nms+zCTB
SCWd0rexPlYgA+Yq+hsryp1nI9A9gBea9H2Vf/xLHZiofcQqWInaYaRRKw51s/Gq
Sk8/VoCQyBGmd8Wc7cb2V58kDaG4cc4GXwL2q0nXJjZZhiD4JMvaX/t+GhSY6Gp6
iXZx7g658pe5RpYTRS8rANE2q4eEQga3eHWQ+0FwWrdrZXoM+8A0CuZp0L5MjUSu
3Z0lzebBAjpKMQTqfHszFliPBjjS2uU8f5K42UGt3a9i9vtB0vWQPTknFZWdVuzT
7f0e+pQougXrj10BmFTnjltFzUroewBBRUMoKgRBwn/o/eIQO4y9Y2095FdkHsaR
pz5uIufsIb976+jDgtjxnF9OZL879OYJj9dqipJO6mzJ2WdzcnSucNouPCI/C+vH
1H1Z/WKrr+JQm66LGOkP/Uly6NKeOyA4uSMzAdkkL554JJzftRp5mOXrf9ImQQfD
7KDdIowf8F//8tLhvTRHTHugaQ1vpw/zYWhOxGtNHOoiEXiSsuQ/HzIXmj9FodJH
n+LfGubOrlKDi94G9TR4VN2I9uaNtiBSzCZQse/YKoq4a9EoHzHteZnL2o8uwyYr
FIZ58ZwvBI9HomE2mkaRq6AjkwpMU3+hve/d1GykEDFJeqQZnWhNrS7Vwq/EdHx4
od7YwhcP+bVmdzsCSZf8Ka7Jknq33PNABdyRRGeoQ9YOryIIxScN9+AlVjciT0Pw
0H+PtJvriUNk7oiluzWOjxOVEU8a2HA3mgqlFwP6mbQoYjMEdWKfPcceaBKeQya5
32OziZZVlguAK1qYDdyiQY8v7f9u3Ii7MulWlSF/MUMZtRNsGc1WY3mKz8JUMD22
50668nkv+vLebPvylu922Jn/KIq/8IOygUVbxBbUqNa3tBh55gOT9J9g6A1hVnZy
D7ifwOB8h2rckaIezILm7NAT9yOETn/ciDbO9/SVGu7+85FKlACVWqDVMHjJSZqG
o9570I3XW8DYuufZu6RYaCCdpThERZwboL8UVuQBVADsIEtSt7oeSwOkSR3b87LN
z5YdIAuKaYBQjGuA7NqxkB9KUP5gQLXFIlA+FqYQd+zMQelMc54LD2C2epZQThpd
ak1Mrcmf5BqjlhIl/L4p1mr6PlPZLccwSlNd6DhISAr9MNfEUili5M2GYD868i0S
HrPdhZvMSgT5ebk7bjdhhFLzhgsJBPL8jR5smythdXsvz62zODpaXPt809r8pJAp
8gEHgWLx66xxciHw8jgwVNk06gBg6EyfYGUc4CVnpa9YJ1jbElEby/NHSJwnf8/z
68qO5Ro0MPvw1deA6fGyzaLcraIGQeNsLjSCuNIfaAGqrRAyvJxHKj0RhMufzh1W
mlLEEnNrFnYNJpydsvFCNiw2baBip/ps4U3vDYdvQTmMwBYgsvnHJ7ZbcSmnhva1
S5zPilLpiFtsRT4Wbi0kgaHIwCWVEaw5Umdqnql7rI8IW68CH7eI/DVTfqUqz1Fu
xwtUm5KdEPaJCxa5E4KxcLiiWT25Pa7pqqKUlEjO4VcbC1Eh5hvUeTNZaus26G9/
17vjMPl1q1mO1LBY263Ll7l6c/xMH5xfdvPuQBEtCP/2Y5WB76qw19z3DFhOUqsB
K83eC7FYFxEjrbyR0p1aEbB79IGznAxPJSwDHlvpUEeX8JNXaGm05hidxyRAokci
jZAve0QFqbVKjpiV6JyLltXDuKy9kHggXMpWVaASxOu1Eio9x88IWv1Iyxizbbbk
GLrscYlosr5F3bO3RHMfgtSN+TUjtU7+U/gb4hHuaZGYaTMzRgo+Qc4teoBHqejY
JEWKbPxJAIdAM8582hMIqBwZiv2h+HScrKr6+NCEdyiq0ensCiE5t/gHvUj8LCF2
cBabpnCc8vrPW2DoNw8b1YnygZDg2yxbqJtpaYcQYnpNkk6DSkTwbBFlFrIYz9mh
TR6V13qcJvy7S+kiPj6S5kRz0P77I0CPS3ElOHW40XHlrjFiHuHU0QELuD3bkY+4
gQZDDOoXN7mCfjme6h2u8yzZ+dHgRCDZMFTSG+y1xtnx34pAEyMQ+kiRxT8e6l9v
YjLqVGctESFzyx3gnP2OcCR7pM9I7Je0tNGGcNyYF+jtk9dqhCpqU8sfOjlIg7b1
lfyOd3kiQCu4n1eRUeSjzwJFr2+zT63GjSydEeir0AaJV4gDGssS0B82l5LHi73H
vNrTOj2Wo1ahtahXVLcpls/epHMyXP6gEQVc9wXuYkQCay4otjEEr3CUlFs8I2PB
Lyv7yeU1S3dENeoOaE2wnLOCDecv+JrBixRwIyiWw+yHY8Sj39c7HXu7tM//2Zot
OtJ//jYeksO0H/fKzmfPeoeLZ5tka2KMoABYb9VKfHEkvGAR301CQk3C9Tej4B8g
pa7gqPJ8/66mhIRQnGIrMmeDypv8YUlI54zfJxKBZfrrZCqeIat6Lw+ZfOkFydiM
fFe15OQWPB9hYMUcRWTVURR5iSdZ0D8dCBGjMg5MV18whtGRbx1Fm5DNtL2T2TqG
3rFCi8No/4x9wqWwrtPJWJFf8nAXSmLna1AUe5N2AaUXz4GdTgfqzuOX5RVZyDJG
KVlkcJ+Cvi5zCT1n7Y1c3MUyLLDNKFmyQnR1KwdiberqXwlayYUC7fvalsrs/l56
ERk0vg3xGvjI9A8NH4BVutm+ZlZiwtfOjMi8l9N2YdtOp8VR10Ht6stKuqQlyC3V
kuBxgLyAenx8jC3On61rhuBWBqC2WmFRDW4v2Gd9nHronsfGp1jrSwGUyoQvI3CJ
9O6GPaY/ZkdCU9uU50yYNLVephQXFW1NeHvD277Xstlzmruk26HjD3iJ6EutqfKa
Pkt/M5cVSXLBjC1PpwuTwW42r51/sBqgYm115shxPfq4kyb8nI0OVJhGAkp5TGmS
LtZ5quwOU0l0R02psBFzHy6U84Hm+jvaCfB3x/J3EgGW2mRtT62UqTNOpoutNZFk
cguxrztsD77HuUmXpcJZzg9/HsOohD0FGYjLv6Ru04IUC5j8cLEQt+X0K5Ncw8js
s2mobihVNeDkZUccjyG3wKz8FLR8rQog6HlAhN329OXU8zg90uLpuIjD9+34dk9f
Cb4fv3NsmyJlZuqfGaM917n8jJpTWY2HP/U9kPd4hI0r90ruNWvvsSJbrJJpvhuU
UgWn3hN0qw+gmkP2DtVByGXQ5udGurzRkZC1xvmIBSdvB5qBofaJU36AEspPdGns
LoDetI4/VdcEawHzrVBWBbBFMvU41kaoWcjVlbXxSuir+cat7zWFC5pa3XvdGdxk
QzGoE4jA8rlMwlPH/8bVUCyKfLc0+I+YfA8MHUJs33/0NM0p+KnyaQ0BkBVm/kxY
vOLoc49HsS0S7e50nRD6aoAzz+BTw+Md/D9HPM0QLPh+/kX6hmjV8ovhlKm6J/Mb
V17gboylJVOV2abSfMG+YnQoOqEFyBB2mydQAuy8guxUs91vLbikgUyQk+O1mga6
CTzzJMNuZVBM05dyzvQMSrxfVdv0FkA1hfhSd2NFtKD8HK/AlGMzYP4dNEV/iLmr
EhJUYuZciALuX5vW8df8gwu4LT7SiROwml4KbcPCupG0/Vvjd/S4leg98RveDOK6
gleNe+t9ZVYzD04l/lug0KQBimyx/iHpwIqGOi3yqisQjRVgB/BZ7OibWOz8FNnC
vcT2hYxtCpW9ItPL/FWngNvNLj1L0/F8Ochfd8m2DSsSmqxFPKAZztAZkuCRT5tU
rMEH+9LA8/u/qrc5rHNGQ3y+Btt+XldthQdl5SRW/Fclz+55jlnXpp0f+NL+WI3I
lQ7SCfybP9xvkMFsnHFVI/F9BfTb7xSAeaITZU8XIAMO9zLxYw/kCnC/R2KSHG/4
dMIdgsi8HBKoJ9agWtXNWrh2ZruTWsgjlT0yaC45kEVBVa5uB5aGI3IScc91VnUn
FtK3s5QR4SWG3K/moxm+qKfBCC9K9gjWgxQPacZVmWJKg6Rob+NfNqJYJzszumXS
IuKTE60TJPjBt86Br5WXbzrA5FTbP1XBtUcmzCYms68cVJuRyZl6Q6jzW2IbtQgx
IwYNoQwkXpwZNq2hc3JE5pZcyuOnDfVBkfofgoYSMQw/r0VNuk5ACgiBuMvwUG1h
jvMPYkYP3P+0JWHkWNH0Zw4O9hRCxpEQP2ZUcmkS5AK6ZrnJugH+2Pl3WdnYFCvQ
kGqouDT5I0hW56A8RRH/XvHmOkiRWn9cOp33C0xAiHEkEjGORWRE4ffPouQ1YLU3
vmFGr1J2NCN79TTLVrCE5Fz+mEWG1jkoL25hoAL18H7agFAwvq1THxU2xHpWvC6L
3UYkWUBZBsrMqA7SPWMCAX3Fcl0OF4YS81yKxfcR167ZY6VY7cEnAS6o3KgM4CI4
U2KXkNsF+5GHWF6j7XNp16/97LPjRLTv6wVnx/6eQ9yIUWtpkOoRDdWTbKO2vRN5
psjtgYfgbBo+glTsFkYc1E7aNfWl/jFlGu1K03i41YpCo4+st0us2okoyY9P8rQn
GDGLc5WoCo+ucjgOOwnVBblr20nypzIsN6weoBrkGKfXy6qfrl1pWY0eFn8YL9XL
0UYEQ7Pz09SvDX1+nmPLWIltcCqPkQQYdqC2rnK7pZC3HihCgnxwdNWxuJAuMhqL
4Y46h3G24W3suF3CYorp3a8uU6Vd8NxtmMiG94WqcO0dnuXqwYQ20W8jK1Vzxv5P
KC49vsTC/5x3AGzljHhENLX4Vo/bTsHVUMZPKgiKig1iiyQtxyGIL9qChklLPdSG
cMM4KkfXcdhk+dA/1DRdmK2fbK65VYrTrEjkFVbIutnetpO5TEdWyL60P6GTLFaX
T8QTLNZ295Kwj/l3r0NQ5DqHVwasjfkZOw3zPsaDglkV/5Efk44WMPkY/1BMyMcM
oTIvMRU5BFlMn4fzGkCEM0tki4cb5PlGNUn1lrg5xwMbch97FaOFBcDC86yRX3nV
2UEtDaM1UozZ6wTS1FVwIG8JImJBcOByMwCS7zwJoLPx4CmBdvGKfH+UzEKiR6xx
hA+6ZH+il8wswXDF7WCOg4/cdAp1t6LrGJcVRuViUMz1qeCM/bM4BRDoLqiesuQ6
ZFCmIa04+z7TSVfSAL+qXqFH4IIUWer1JeNHg7JoAvc+075cUl2NTCag7k5sJZaS
ofBgRK0WG7lQDyJRwGPJHMq89WRZlHVVvla8npAH+BurrYLvRTX24TOhk2lxeZi6
4O6Uob4XXFNKA5AyjXtuRWYxjQUFwToK8HaQfKKVSMpk2247GZ2jC7JZpINDIBct
I8tg2py381JnCuI/FkxG7qk2roJtOdJoqKpe+4jDraTnYXdl7uv/1Rz4qJPyWPyX
jivJP4dsyvrjLbr2Eaoa2Vm5QiDV2f0d/rtBxnqDIxN9r62+349m5fezONtb72Cu
Jap4nM3EC86dU2mpvqFiBClF8htdoXKYfRHyVUzFQWIYZDH+RZ2LOrABpmcCKBLK
q9wi8T8719Wv14o7km2RU+sz+1YTJ4Zh4DACv0gSIbsbZ0NRbKbDS3m8sxPDbZMD
MHNbFHqR1gysEP+ERkzg7VsBZw6TZSCgEFR8wSpr/MJJ0ZvAMpW+KpRSyxoCdc7g
bDka+lX7wGtzdhVrc1TGS6Imj4S0jw+RcaFSWiZD700mLrIoKfwKaU3Rbom/C8sG
9uGlaFRM923MElV2q3hELFC/xHocl4KaAVyn4hgkOXrJMHRlW1z+lLxcMtvbG9Lf
wsOr1iIDOBPs5/xQEuXGcs0A8EAf/NXUjrKxWQWWa4BNr5+WX7YYsBxv4k6hIAbR
FA7CpXmNcfCE7tkL8ph3m4LfXYaPe1SBjvaMFi9oWi3VBVUt8y5GC+GuyUgYu4gl
QZcxDfa69Q/rri5g0W4aTc4CklwVFtilNfWmV9CwXxBJc2NEOYaVmH8oKCmYiNxX
KomptncMxQtjsM9dT2NKi7rivPPvnblKtUjntPteSLJQBokFH2K0QxhMFSUvwxMo
dn7qGlti3eurM5DyAigmjcHTBdx5Fr+YhqRrKCgDpbINv0OFVLl3ES4/WHmz2vj/
16alvMWI7IyR6N0G2wprVm1p1v1iimeN83dHxtJGD045RsbEtxmmteTYlRLPhUiJ
9kIDrsu2qaIpE+q14/PApR501ZPtzwUnXFMZkizquPxIxb7KFEYzwU5QtLb6OlVT
kNzM+auWSDA25nd0AQyA2wGFHTRvvC9D2BoYt2dPVNXG/1qMNu6bxYoBQg/ZA2yK
2yox7qnqFhF47WjPeQGXYmutas3H8fWASZ+c8bYeUugeaxykiSYjE5QuON4Ko77E
1yfW/b3p4bOeAE3AzyJfD4z+PEqRekeNZ1Lve6ZRElMCwDkHgLp4dneHa45ATQ8m
XOxphZ1n07FYeSItpwfHQECSdn/scnY8iF5o/10BkjdEjBjSI3DjnYfYCFPxI8gA
JupUcdiR/N60x8oPp57a0vCzVSenFb6qRgkPRsXFhknDm7mFEY+MHZru0E8AhxUT
UfdYBYVizY+aplTH8d2My/8RghfdVnbhpAqtCh7sHeeSnQFlsAAz2gRd3OtYyuU4
l2V8RO44F0rsNvqrxFHaunUnov9PllDnfsPZLfQ3jaq6r9fETneOxRYyCbKbNmqI
DmygYVwNuh/aAKURCZitX6llYL/UAqwizn6sM+tEetk8hv2KgEpUn8HA+n65HHlg
rYlxQJ7EQCWXsCsUbUQK+F0ds7djF8bzUlX54fclk/+HLsdt0xAt+i/8JbWOFUew
BicvpDMEH6QaZQjBVkvBQ8vvdZTZiF399qd8x17GQ1JBhaYCNCpAYtFsuXPNhFFl
R6LTWpTW+51BZ2wgvjTDUL9A/4rLKMuJjD6WIBBViDOKZxJs6fBSNx7vOhRtZMRU
9I427XpVWwv/HQo2uhl8HLq0CTKKVySXEVmme5LPbPfZYi7BaWqpBCSZ55pR5DYB
zMGOgmiSb3eZKrVsohs8NgF1DPKCXyDFi0gIZwOq2lP80VESGTQ5j2F+5Q26wb7i
8JJlSnfgvBLBL7Cb1CQEJDbrh1c24WwdM1VGpM/hvqzYrP8tHUGDoM4KnjtZK+27
QsDZLx71MOyKGfa8y9m25j9xpSVpjxWdx5JraNRWy5eBK/UIuNO17BEircyhdQKg
xWECJJaLbAJXiydCAc9xkhUj8+v/Gklo/3vuRvJZzXNO+U2JB1PU8Kt35KUbU3wN
xyP4KMBsiY79dVEQYvyqytZJwyE6/4OUwJ/Vc34OpCTC5/CxI23hQcWpei2dnqmW
7ed3ENRva8pa9LII/vk2p8UV1p4AzW+MuemQZLoqI00MMRIgunyVWnYH1fAJWD2C
LQ+sp3yV1ttOdFvhSNumB00ofHVOMQosy1iVuOZ5y9M7VrKsW6PV1VCIVKTBA4+d
omXxQIu3Qa9yDv+C8uf4MxoKT6YoTFMjN1arSlc4RQCuGFZ3lBpu+40V4/KZo8Ll
T8SQlC8Q1orc3jiaokFphAy/KSEEFFW/H0VUAEpp75GG34dW/vSjk6lPpJA/tk4W
hqec3HaaUtNM+tZL02dobWdufYHdDM1PsFJPcDV1JlSNACNTIEkDt+5wqCbdMhtm
HVbgcuRwAJWRNtiEnvjOFdo8FtsKzl3/z0ezxYrKlwyulGF6GOf8b4G7IpKDqECJ
JFXLRc4iWlWUUL2M4FZZpHE2wkjAYetD5dnUuOCBH4fdUp+324Ya5ut2xl/ePpyS
rq98tzFPDlSFHr7r8TwfUxmQMuV2tguXyXgOxEx1TiYqUwVnk16zPN8F8PX+/t0B
SgYmlF9p4DhOH7fKLPfkYAMAtCkplJN6tNKr1jcKrkZddchFQLrlhY7zE0aD8Cqb
E/o4ro28xJOS5coLNKN5fNvAriLks612ujafVIV8HciZzfE4xsHImwstogUUp8ey
1Or/KvyFqgChWx67BUg7TW0G2i57ZE9YvpOtRAnNvoc4KqDM92aPVqnVfqAfFDJI
BpzQABjw4jFGTPq3aE8u6eJvBZYMrfbiinhvHqMR+dsWyG+ekLlcz86wo1fxD0+z
XTJ8YyGnl7k0Z180FQt1nhaRNATTuYjtLKgNUx3LPyfO5BoUMBfsTgCAYylWKjNQ
5KuyIH/6SSww7cgdwgCpkN3Cs3tDpwS0iHkHtH+JFXggDCVqWDfDdx+4UkQM/06w
gFSpB4rIgiPTAMPhem/CvU4QuAzYnD4vQoXOjuiSyLP5vsMcaRWIoEYcQeX771Zv
SQj7cpbGPs0MPS6lOLQ7G+YQha8hCE0kKnFckgGnJvEMx8rCHUWEZjTeTsQPQpkz
x/PLHL6GnY89PPeVjrrqoZINEsBBVRbXhWgTyUa+DQBCVz7zIi7whv2JXLIpIeJE
8vRBDW9fshQrtqEvAviEirfREnkqDyazQpr7r5zDzjCSTu1uinW/QRz35bJt1j/C
CDDpshrlSh8LMrNvhNhpfw0QNhMzhQNu8Z+/mLJRjMPllmYeGOb+8ezmMjaiElEN
wkfo4wK2qmawDcuaqgiQsGZPljqNp/wk9Othci6p7Qj2D1XpeEElK3pJ4Qz10FNJ
VKHs5WTUEvoUYbsucVkhgHcV1XJfQda6MxKNsGDY+LZCDPbmh+FngdrbKCiSldzi
`protect END_PROTECTED

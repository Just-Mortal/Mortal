`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FqX7tX8Onew3pUuLtlJSUp6qwzqWMxxiE6Hi98kO0gXwtkviBUyPNvOzxxSCon6V
LEBY00SlNukYCBNdBMj3LRgBeohFwModOIeG5gVk2gVfb5l/IMIF1sKyhOyulmVj
D7RJJuImDwXV/NRCg1SijbTt1UiR9jYH1UcHQmGBuFuWGxVEYy4kHjujGkUhy9E9
7vG7zf5/OXwwZ6fow1ztX1FTAK2k5ykJ9X2iQjkw1CsgSrMDggk1aie2kuHDaAsy
UYj/bwpWMRIYAcJ0Q1yhVeParv0qHM6Ntp0TgQygVln1ZIB3t5u4w9NF9E5p50lD
iFkRBy9DN4H8SQFuRqQseg8a+0XNfzRQAnp61BUs+MqPuCVJUCYeULS2ikGzlRY3
WRUrKB7UiUHG+7tOzRJ/5X5PR+xtvPZRypQOUpe/4VE/i/d5plm+btYLjEw3Li0L
yd5LMO0WiyykQbnNQTfE6Oa/5lsktlfLtFY0EzyBza582VkS07y8P9ZveYwu4QHS
W/+yra1WGD9QOgly2xUPP6dmCbzPvBmRhAqlIHq72ZyHRMVwxt1bLE5CluyyKVe7
JqK9RWch942dI64cSc/ayLjEPhWcPU2/DD2eVtZiXVzfKlybcj2Xi7EAXjNYdEc2
m+7UUcZ/BohEoIEmludu4v4zqqcC+bTqXD3IT5a4I9mGffRzpgGrIJDmKjJvch5F
RHdZQ15HO7fvnjwjBl33tq4cTLB7Fodpz5HXclEqX2jCArfOTB124qCkJfirAH40
rKBhChBz4P1Zk3TJXyT+840nyzmepHJMThYu9eIFa5GFmOcnXlB9x2PDoGYMv3t1
Q4NGagWWasMpRvDvvoGhq6A4DKP1dJj3CUOfB2b+21y/DOoiD6DrBUcHSe0OeYBo
NCOjDQj+PR3oQOv8zL4oeuh/TRzW6HmQLITMDR2kChJtEiaSbXuG23Eyv3iNLJPR
/iaiojWInf1CbfecLFv0WH8e/VWKW0zRUelAckHgyeF4gHxb2OrDUHqeg5Yf6TBT
pfvV1jYoUOdM1viJ6rjY2uwrmFoEtr+EPGHGFaj3kpZYQaUlqFwm875mueNPO5QF
7iVbcIFdCTEbAyZ8nQ59y5ZfkELZ1rhW5J/r4LyoIWSN3TmbKV/2323UmM2futDU
ttpMm7aDzoNjJWfGdDTrZwNr6EqLBW8uTkao/2Swv+NnZPRHby9pXNK76fS+4lot
QTjcMS1sIyr6LrzIq8Sp0wlw2eEYw7X6cimQLCe49Cq3+iJgJiHczKAbLlRAUlbI
9VSfGFJvLarAsd2I9ZvuJijRXlWTElbnU+tYQo5lhuM3BdnkhH8gYN/jGn/PlBm0
RdEgWfus5vRV/SxnakDw3Za+WBMQ55MEvdD0bD+6eClJwxE3x2RqL+A0YZ3WwPrC
Pb6Q4fMF6jatxBJxW0QPvKGpqmqR2BxqAZwLt5ArnsAq/Dq/bA3axh9c0wVKDrcf
vWJUGjaR/P0zd+P2J/HZN8HG8ndgRUvXDO1UNndkLoFRFOUi1oUojlnpVcPfOanS
AGX5SXFyn8HZAlVwIedJcunaPzz11UDsFLa1Sq1ckwJQE/ynjfDFoJDroD/MfNn/
LwVCthlHLqXb3TRDlsgn9Q3T2Y9Sw1sWZt9NAsnGlUsvXVPw0962nMoXuYfDDngS
N7qNmr9InmBVBawfdSHW5OlS2FePZDbzXzJ+BjZDN1nJE30L5y1H+xfEBdKJjLfp
0+S+4NleYT52i7J1Mg1ImobZojonOUvCbUL6OXXce4Y8uJBnVuP2+smKCtueyrCm
z/xbK6AK4ioRBn3+mdD/DbG2Hk7ids9GdHdIkX4I5XBe6qvOptZUyvu6EPBDxP4c
Wz0RqC3Sq5KizxmwwHwMOIptpT8Ghs4oa2wzSINq+qDMPTzLW9S57w45Piv93MK/
VZ1higqoSV8UlC1Bb65m4O/oajKP3H9bCy2/E1AC+wRbPOO941L+EYYM5fBbrQaN
HZ9OGDDMzJxG0+yFpR5RD3VIWXrJLWSYvMzaFScOk8o3zsvVRSgNtpFbHd78GonG
MgP1cPF/Cj4wjuU+7sglwi0IBWpWIipw04JRzR/MI+DQOS+vgQo+dGQyUPnqTDnd
60YySqib9PL59eGGm4tvcMx/DbM2iEZsOR/5eNDSu3+6r/924niRtpRrNf/7jGxm
6a2AZXt3L6JV5JKZEYrFyo475wyJ6Ph7TwW442zUTdLacN4xPKzpgIkNyskaB2e1
jIsxHd81o2x5EjealTJqkv4d/8e+FP/UWpBIE9dppkc6R058y9NZll2C8zHLoQEE
rTK+9FI9XXz+TxTRZvhC4WGb60HxGCDit0QD8O9th2Cix5fZXJ7vsQDrZCY6yQb9
GrT18hVTjvzDYP6xW2pkSf6h4YYpgT7Lcc2Og5vsE5wt7HlaaKBRs2pdsRofrFmN
g/y8+zYEB+dRFOnyWYqV33Xyj2TxueYaNIjXzpjHlDe06P74frswhzzjdwkY/Ja3
Lg5nX87NsBPxfk0LMjTc2DF6CIX9wslbIqpbw9tX8u2UTWdZ9h2XoYJXqX5xl981
5BsN9m0hShAnuXFhScnzDev3EXmRjurzBSOpYtBafHIHHIkTu8/QVIgH+put+DS9
+j+GpiXZIIsE5w6VXDY7Ea33yFvcxd/HiAS9RIHJn2c0oQfcXS5LhDjdMWNCKEXV
fCNGUZFe3aFsnHhyhZeZo/SW5r0SAlgflcCb5ery8BLUkdg2w74p5jJs1uCoVycm
K0IEIN1nVZiP7iA539GuYEYt5f1Dxex+hvz9DKfIQFnhA3ZqDvSkUojmh9+PBlT7
hRxuCXZ4Ois6IUgk1YDoLkRfcVnQmNJ7lPQHJW3gkTpcpcwLioxf5NKd2bbTBIJc
atymO5/GnyKF730kvyj81YkR0cDnpOtqETiiEMeRyEHm1p5djMqDGWLUqcf/Z6BT
qXxom6NFv2YbKnoOlUqf3bySmbPHOjjIfNA/dIknX2Cxnu1VIvW0oltrZRY4XTml
V3LOycJpQC+ovApVysCdpIF5Wj1uDJ9f5B5XtkCbfo+zdm5V5vxOodlzKuVcb++v
hdKlyd0G5CBPyfEif3e5l3kLUM0WZ/Iwindvz+WrYWE8sx6rMUgYZ3ipYR6S7exg
/ejKtiu85d2/Y+NHBtsJ6EpjKg7WuFoMYgS3V7BQbI9N6X2H6jLfmI0t4aARMm6u
ZMXwHUMoYe/4M1VN4r4FKFggYC6iH+NtbUpaMeR2iMfzF6NuragHVMmzELwakuW9
V08Bd78h4LaeN9g7Ch+U0Df0D7c35mvGYww9OAzpeT7CLzacL5z6VAFeaQCBJ3n8
Yc9dVppAE4xJkHZycNtSPMw8bO5P2socoD4mbmuFYJRtWNsVt6Sxkk3JWcb/OPPd
EvjxSDhW5DB1Hc301T2GxVVfgfu2S6Lq4bv5krE6VKAH5iFUv7skGDTNb71NNn6i
b1wUTyP7dm3SJWX0axZBAe4bnOa3mQI/2L14g82OHcMnBaDKuFzQRYU2pyIgrdtG
H2fku6jNbVXmd8huas9+AZ2ySf+Eh+MkiQTrHCcAvI+kUvoupe6JS6AS5ktGjbkX
UgWPkwQq1TyLOoOgbq/EXibqawTIAssQuj6reaM9Iv0iHI5aKJ6k7xK2R50XUSGX
KCmPoHgUesaiSS4qwFPMEC8qwoSSlDQTucFUKLH6vgMb0IoaKZ9s9seT2Mcts80m
3gx4nMHt+T2PTJJgy4Z3YL8LfTldXOfMtKEfRKj73gzTcr4J2H4z30hMbunmXVn9
iFA+6ynKrsXNJ9gQp97617FhZpAAQC1WNwF8XrLZZDVel7Dp8wV/YX2/+8s6avU3
TYdbcJhSGPqu/VCDbMDEzjAHy3uUQykNzph27go8QLSRbpwiHhL9l1WUO9LgdBq+
ADn8GiUo9aiZzSkN/rZCrWqC4dNrgz6XX+Mv8jwmYKij+OAvAErRvJ+hoEbOs+bD
taZ+gVFmXCbn7MH246cAQNgoiyxxVc1G8C5tpOVsY1KSSOtat75dlr0R8dlgMBMo
82RLIfOlaTvQWfKq2c6OaZ4Wq0X+FYynLS6RDMJ4mZcz7bqP8Zh275dnnK4DFPcP
xTUpWVmq7oWz+xDRVmR+qqUCuTtzM2OScngNave2keVPB8ORHZG/uAkvglD5Yhs6
d/r7Bt54yb6RWmZKLgOeK+nXdZgSSrgQCOXXF8GYQjmk+Z3OWUKVjWy5DTYYTbw+
UTtPYafqZw5iYomI8ZPn0/BTEDiPGHtFXQ0Du61ywV7BK9//XkxuL8x2sHxqLyl4
S9iIOkhB2GlOmoOQ2VHYb/wWI4H/L1RBko2cci7AMd2RVUUyW+JX3ld3Qx4dqTJh
c0ox1KZ7ecNRpgdVTGSL5w+FEamc+Xd8hpv8aBZxalotCbsSqT7OgZPExpOVfrKn
aqB972+6iK8ot2B91LdXfFLysH3Sg1hwYo467Crl7jdg943HPzETCyj+ymSnsgMH
`protect END_PROTECTED

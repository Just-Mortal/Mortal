`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+y5JJJklJ3dTfAw5WmA48qlZ9EjzPPf9GrP37jSiCRJHQJit6k91Ryh0Yc1Qwrt
NUQVyFLgclNh06bby521d/wXIRMKKBETBHZwZVZmvN63wg/UIO4qt9aT3sukAVSV
5ZVD5LLdkbluhM49gYfyFKggXSr/BVMPve2s53d4kt8xEbErLs3xaSpTV4E1WSR0
C2QfmEeZKO38sJWYXvR3JTT3xsQP/Q6olIRsynFT07UCUXVTkK7hnbGUZl5zjbjs
sPe9Ncinql2yJMzLbItjsd8aOO0Vqzex+LeElpbh0/s1RynKWH+ke4rCsB88U6mi
pWSvXXHPYyu+NIKRCSp1IVu9BpM9AXnoZx+A0P4yMsrwOA40vcn1qGNfaMgXVVPb
+3eVFXl+hPReY3l5KRb5v7OlTbkABlXS4yKlaROao39cbSwJqqk3zCy5+Fk27/g1
myQKMQCEL+hsWoYBs/0emR6vMxTNztiEYJDiP7SgqdjNnd9x08xRmD6jVAfi/vDm
J0Nm99SMlYo+IlY7LSnrtaq3EYj64Rk/iiiiQCABFv8YaF36/KQhKPpbMwvVAfI0
mpzFqSeZlYhh8/8U89VwLeIiEYl3ziIObiwLQ+DZfhubca5qc6fdHqPQQczZ8SiP
c3TP74BlqGw7e6wYb2b8e9F2/VmLJzDgeMPaknFkTBbkupGK83nFAZ4MyH+/Iy8E
+AzjrjOciZVJmB8ZY/k76myE8eYGYHcE4QbGKNoee3fj20ME72xAVrGIeNd1L6lL
fNqwP1oOsrpMiU+2Z3PlIRpse1H7S8BorLylh8yve0keDnmcqXT1G8S6juaPQ7lC
5CoS6tW880U7cuP6YRfqu5vNylOeCASJzlal5hBqwvB1D0AiGzmU3pVXD5uPXrAe
31Z4+ewbUX0lsz598lFFHyiEPZcrVd68YOqxt6/im3AWHFC6j02WG+pGgBYbHq9E
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKo2URZ5FmEFPdz88GjXb1IfX8I9yN8SkswsmKBViXwUOCt8dD1JDUYg+M55+JQb
Fd8PxB+sWGmEDWx9qU3i7NwYp4Es/gUONw4Du94s04f9I5BeYgX24+bIhCjTaF3Y
yy0jNtLfKPKZ9FOfvQhOHqrlvl4+3qN+Xdx7D2jrIwRMDRGVGzp2bPCzqDHPm6jX
gCEcPuE0fe6eZ+Mp4zZWfa7tpVQaTZaztzs4PyjGwCS3Z7NxvqTIDI+sE6h49IJ1
WoF8wDHi0C5pEAkiMW2BfLu6T+w2JCBDQGOJuLZ3cPMyCUq5RI9tGK+vvcjOkLTz
5xXgFFrVp4eI/ZpVJQQEXw1xfBgRHxN2jcArdGkfIFK2JB0/IT0WnzDe3EWE4jy5
OFFD7ozrtIFTpQlsZFG6iPSlpLoR5dXZ9eGkIu6dgtCqA+WQyoGqFk/SmHf4+wSq
oEmJNlTx/aoBBz6kH4PthMg8qWj4EQe+A5lBuE+OV51G1EVgqVczV0D1xqi3aCLE
2JyTZy/Xho/6zDgXzMOJUU+xF1HzEgrhdkGDuxjji0dSsifW5InMnvLVntpWWB4r
j6seyjM432vXqu6UWQGkG16iKRZdj92lTpE6ocPvnWp1oVoQSiV+EXLdnOBxyaqx
3MpIRtJGbZaPV7jmWfxSPlUZqz4YBw6Qqjetd31Nuy6x9DEVALNOiUwbiP7Hdpst
G2waxGlGEmIxFaZl5tQFd+pYwZhmc+epWB+r+BPr+QBpxBAZtVlOIhq1DsurkEmW
fJ6ytAu0cX+TzNUTBoIqpWCiNK2rurOlq1w2ymalorwdA3J8zRvtzfVO8kAxCjaO
lDGZAoCb8FxQ05VFvT3nxH2zCVGbF4jEBJkeNG8KHqf6icTH4KddUsFPmUEl6+8D
UZiwhgCWIHBWL0Q/oiqLCSOfDYhG+EghOXR52GLio7992OQJ/nxzOiLUTB3h8c3g
HXGE7kOUEZu6VXA1sgWokp82VMGX5t4yi/M3SVCJQXElkH/xoQeLXq9mWc13+Hpm
pj5x062bV5E68+uOpoFXqRxCZ1ekqDRvdsznHyIelMEAW8h4fW21iJ/iB1agLIE9
ep46IE57g0MgJJwE61xrurJ0s7qXIUa0JqIGMcnNGPJVZQn4LD+roNnUHz4eGd+p
6bRFxcXkpSk9j8WbnRzQyzhHV+L91b7hWSAUTAErRaB96YBOXMb5ZyBi8tziX0Mu
ghfeWEWZdc6lzbCGfYl9yheUvn5aLlZ5x0uzHUqRS3pEm9UZoVCPS1Rurs9EasdA
yLvAYZ8Z8n2wALvmQGTNz8T6iucA3Y/ZCyNdUyMTbGA2TOrkuRBUsJ2t7K2JgTLJ
acJ3F8YQZUy0qH0lUTyat7jaCCBf22TOjGfZDmULfjFcT28mCflbUJA/LfoXgCO3
RkARRCiBqJ9SC/2Eqc4NJsUBYeGbUHkzLleLBg8sxMmtzpNVj6BnyC+oh38npAvB
xjU+aAJRWWir8J0o8ouB9dG1j8CWlYZ+zNo7eq6kb4MkjqrIxpJ8n9oG8qi4hKIs
jiI7M/xVaZ398f2pcUvYtjLCZ+mPsBTWihs2a+s4ximyfdG8eVQ2fQFgXMDLELh/
+AreeFZEsVoRRlvNQwRKhCE9u56oCPyND4jEkWAbv77k4K2p15i2kRpSG9cBoyMy
Bjpn41wpjIRgLry05U35rT6VNh0pH8vVgjRTq5y9oapq3BJB0ubMEZnp06M/Aa5H
D4IcUr8sOweeKS1k22sKu1Nsjo2WCrliQDvFodkLFEm8aQxnuY3OWv1QDtoPx6q4
eYCjpKjZmBePWTzqzxWAwhRNb9WlNJ0lx57SFYLVGSKoeOex+BaAzBYsBJTG1vXw
dszK52bX/8OEyET/GWpHshI+ESScm4ECfGqG4aE4HE6ui45cLjOSlfQFKhlepdE3
EPduC2ZK8jK7Yow5WmZagKzgNwRp99GPI3tY9oihhnghpfnYv9uk1Dlofa0KPHqN
IjZ1RgelFs91ylMZyTRwJ2fldlHsE2Sl3s6l323gMpwk/24LaI0VXNEXQoYuRjK9
HFzLpMHDPnIPw7rH0p/dQLBNC9CdNZIyekR1Yvf2qtdH70TavpLKkL1/abLMh9iS
WAYPCgfNiWe3q2Vof6yn+5ARyqoi2rSUE7acqoVtiNkY8KxMJPTTr6TuZS+S9JNZ
LAV5MjYuincw2u8UvLU3WFBvz6N1uU5rHll7jdmqm+liazyGQpUD/a/l6862sBL5
p1djPoMPVUPVYhb2k43o431an9IqjxLIEjBM9PwqQyZmR5GA5A3RvdFTB2qpg6A3
YuKQiaJfIoYmgI8UeyAi2UmZ3/N7QrpewKScTrnOYQTndP/XG2Cgbq8t2AAGECAb
REYhWckhlDNvuMInsfyPu46UcS7aYKtnBwBjHas1x4Yc4gybyGD8LpYvSWla28Ks
vW8v3zk8imFhGgTcdcCbeFStJsQSgwMVbE5ZrUQRPy+VwB3EiBRdOk9EsjTqYZQE
LPC9172EyJq6DbE0ED3gdqHzK4JSR0xdoXRCPTar1afXPxAEO+tKxWk6GQp5x2tp
OE5Q15nCpRoM3ks+o+G9HyAVNWbQwvsORChnqB9KNzFQOfRbYGnoZ/WvXb0ObQJk
z5UhG8U0WbH5b1ZptwTcgng3Zm/dCQ+qGxNay9HYe81hE0QlQ5iX9amSqrVOVN7u
+0yGJzbFzx0XniFx/0AKnMiiAMWbmGG9PW/SAJacd1CLb4C6YZJ0tuoSlfuW3gbB
pm9C5hm95t60wd1/MduzJVmyx6tEN9VAKFqVfEixwssSch3TMz4sWslfJk2xAYMK
Ik8UqHPHZqOQSfbsUpf3iQhgAfrvS/zkzlnLeA31/489LGngv61lUb1cHiEBQEpu
WzF4E4E7WAKg0kgfwipRTyjXd2drk07t5Zn0gDk7rqoiMOIPDivu9bANAg00J3k/
vKtF6tEYHndChvZwGtAEVA5hvRyk+1/fkxYOQBpeQc5tPOW49T4DvFMf+w2639Es
A433lOdbb0WPAEYTiguimQ9y7N6jU/sqeh9V5HmvQbUJRTIk6aPU6MjkGnW/Popw
STpDKNDAazdpviHcg6WJeBUNwEKZZFlkNDnbM2wLv+pGTgEiVWQCEAsoLfrCTJCs
X+IRyY6QYZT6VcizhZ4P4HU8DMocAIqm32Ivqc6z30CdIzmrRusO0rj46jklz6NK
PZWY8pYrZL6U97BrBrzHH4UvV+klZrbjEuJulvI2N0xxy2axe6bkrSZuVB8KSH5r
5RCMvsimI9Ww9ywR+FRtyIGnRgodzHddbObl4Y4HZswSxBKCvbSfcgvUyrd6z/S5
AJTKN5hSlXuXbxOK8wGpXIh1w7MrSt3kXaD8fuc54SQh4UkYGbfiVW9QkCNcjdpl
qx/AZF1gDxb4/sweszMDBDefxlvKALjPexwp4kYULIhIe34APUCK5RVaRtBntrVf
MyUYqdSrSdNGOkCSXFlQHwPP/D65pWWZiO8r5BGmXd104BhjGA2m+jAU6/kj2+Pu
5eUVr/WWUDkGuxE7FfkTCN8UkRa+GlmwpELUAG+mDtoxXcuC6OId/iRZijG2grNF
dyQbnzOE7kq6K4gJ4CueoWKwQ4yQFrnNWGHy85tpS8mF8sByVUATlgv95xDA555r
F+s/wBDud9nwTruqfuLTimi7ZwidOQs6lk7M73u0BgiG6IJgweZx4fl+dkCO5oRY
bLl17cfVde7OGCbEWnSFB7dzDEMGt70hD5BcyfYYO/HoGrbMQCVn+Im6AZ/gQHdD
cR2Jrev77PQpb3+i5Ayn2XCIaAI2pMd4eDAuBZgoQ4KNZSF5/MrHMGuspA0uioLL
YJL6O6tr2f7vaTIpTzQlhMQSYh9nlbVVXbThzMPbSuDqIcCXr5HsNaVnL1zk4g7d
k2PI6cR1m4FUmXpQLnLU9vUeaLvYamAvN/N44GRZodlFf9o1G8KzJe1OApAWnNSM
xV8AETSumvBZxsyzdxZug+J0CmGaf3F6htMLifWyWCK4CVHevmknOBWdj3L4l2Nk
gT85tuOkhtkTy2Hfb52lSu8Go98bdakPlKE5//6TOQtMJYuTg2t0iZ8uCA8F8KLK
iVtbp8fNpLVvM8N4A+tikRbCSpsvgUhiGwbkXOHwK8G3KT0D9kkiA4MZiXS7bcXV
jDPNpKv4Pmj7fc3FFmrZS4Lu7h6S1PTH9lf/L9fdVkKKhJplDQPVRxIQ5wfV2bhO
iZl8mvOzxH67LoW0swLq9n2keP8II5R0bztRzswk4So6kCi5D814NmNHOu37s9D7
tD5YNptrCXWCILpzApzEgM6KuC93H/uHAxM3cXfDU1YcJGVckMpnhaEXFZZXzQBN
zjog2NwU/LJsBBtDs96Ci/02DZUn7UO+JhBCDbRqI9ayzhdpTFI1eUPMCtIutx4S
TVSwyvUJ03R4n7ECrh7CvovZJeh/V2JT2ywsWkvSjdWylQvfp/F1hk20d9ozPDPJ
kIqrXzVEclMCQjs2SJuUsrwguOndY0RhXMlgJGIwKuEA9FI892pU5HGnz/nt2ch6
cTkiB561IFgxl965oa0QkFUQTDIO6UA4ZpSglgtcy5R69dkkXp/GoSrOYqwe2sCr
1wijtCkZogJZ8s9vTSj+4uoCWbGhn3W2yb4GUeAdal/CtyNS/3wCo8clov5Wv+51
nEGQzFLPmEjLqka6rbrF1HaMc6ZV1v/DdUk7pc0BTsLiMXLqcSzCZnj76/lvMtmY
XVgkYdPuGB+SFrIwfDfiRXjkMTHxfRtmR7xQUf4Ix30yW4pCKrbTDfHHOLde93Jz
TVbZjcyTpWIBtNaLVlXBGSoivQzo7/EYC8hOsL37YGB3hmb16AbnxTOb/jUnhmwt
heKsBT8I/YuelfHDHQdAcD5/PG5GcPMJw3SK5JSAVGFP8zA6P3DcsstEbIbCmgvz
elzCmLvyFBtDKVj++N8J+LqzQf7C+GRUuAvr8dv5YAG90QwpF4npPfuVp8iP0BAL
DD/sAO76xGqOf8gW58b/KJZUWwF6wb7cXjW097HC7uOym8oYO8IpoBnYNHRLJlHE
pxmxuKo6FF6psQIhu8JSA1FsGigutnTkgaG8LvKpYgxe1YhFxhIkq6N9g9PxCu1A
7RsYDsr6LRBKE+a+ofZ6SVgENzJ9UxzM3GkRJP4PieLrIONOUve+6F64I/t84TOa
X2R+OVqLO6ue5tuVfMqVAmfR4Nr6S7/ZQlkKctG16XIJjFBbiI4ksV/zbeu3yzHK
ctP/I7EXBCCqLfR+/DTF2V9PON/okx79JZI/ekZyVGh5JtWlhbMrpXfqxcS1coY6
4nAsdgxMHxVUZ0qwCpQIlR/QHdKTf5Dv+94u/ZxI3vBAwjnPOS4strfivD8HMB3H
0bYbCWeZmyVZfcwlq7U7x1kjyiBxd1nn+yyg5XrMjwLzzVWTeVRsO1bP0K8+Q1XU
tGN00D3QWFJm8nagF2zQdy9OqOFOp8FTH4UVcEUc6V+hlyL7B86tuB0YOH1FmsAK
bcX5zF3ZE7CLA7GORqOulgXweZDqxJgAtyY5dFHdOWxdxFi52zPiCLRVZBiXU6mA
T3edaCqPbUzVe2DxBw2QSqbaqwPOrDpkjbsX+IWg8ZMCyWPXsVCB5BAHNoz+U8/8
EjAAjdhbjjc7PImy0Gxois1GcmuZ/IVBoj3jmbS2OGT6HHm0KNdvV928qxmdcTND
hfgEJjESqHvOioR74fGib3x+gz6ov49GNL9RztYZk3pC6q9vqlr5HyClzwrKBiKb
F4aOdYhQGwI0B4WCwEk5YCbd6PCEf3VN1H6+JKp0mMAjTuv/wv+0D09SMpy7opdc
l0z51GcNVMEb5q0T0VV+8HGeXA+RcSZvgSlKeHb9R6VYNL86ZiR/5ikkshOVHhnO
ZaOim7tyW3GpNm2vwpl15X6o969naw/9npyWPDpD0al3QMrhWkxTB+8m9YoRxr9P
8qDbDB8OUQdUpbZ6yfkXMSRb+4Jn+23Jx3/TbDw+km7QKyi47M2HUaLIJ3/7P/XC
WcLCmWWnp43xi/lbKdJ/8lLTV/wA1+q2tM5CaZh61Hjm2EKGIvNF2XOgRgxy2ixJ
8VvX7O3ODQc+VnifLGHK7SmS0LP80oSk7/xS14AMEpd8pNbNIrFZV4MgkHCAow+P
fLKRZGhTtG/iZltwo0g190FNSyrbqqq5nENTSjtazVxEjN91NuptwEBci+ipopZ2
8LxkP00ZAgGWiRhu6XTYgmYX6NRcv/hbg1f1rQoKfWZ7FgQbIa2BCfESPmquLRZa
+Xc/iMpx9lHDv8rMTzKzpd3BFfM9yinsmcDyYAqjb7QLHK/ieAPSsgKs19E2Qb7U
mZZbRnGcI7EHOOzBNN/ShjSCoTGext0stH2Xd9Oa6mkuRJ+Jk60zPFvJ9zB1Ys4k
J++2RmMiD+idpiv9RahONxQIwCjtE3QUTm2kjYNp+YTyvngvJQ/nwe5PUxd94sBx
f7qEUGzh2b6/k40O1sV4TM2ZNjoMgIZEczP6qk802VodUlxWSayYa7WmbNFsNuW/
nIUKnSdIpAR0GKLi6VXdh+bmhC5PnQ6jrHV4jTSHJSKLqgTTt7qKY2ezKV7e0TN0
1isRMiA/OxNMy7qiWlq5q6JixGSFWP1LTHB3ZJHQh1VTBceROPS6LFwZuYcpQQKg
u9cbNZW/PaeOiiYRQlqYiCyEJThPV37US0OG7iy7Hme0OMxCZH7Lqj3fBrbdoNSS
SVmzIbsBV6JRtOziRAH9sLIc8uiRAlUy7Imu4UQy6mBFFNXxX0Z+xkuLr43X0EEe
7RkjnK/ySRZuvDpNXUMa9jeecUMl12QONHRlCSoPMqSc/OFBCzZnfSoGVpW925pt
ontmPNEvIB46jPZOXK/WgMDVax1dNHnWyriwcgHZyo5B57QtGC703ewbpfX+BnFv
mA7wMlgIkf3qNmbYscILRd3lWTJJgaCp3gBuaaZ1xINmmb8w0WfZ+rpktKFgkhOV
SghCCcojWBh/EBD8kGdP6ni/jXljhhOXifTMJ7KodQLlkT5vpPs6mjVbjfW5OMkl
cpQtqRyvV4ub3wuvtkmEpOxHoJ2/DC/T0MOq7QV4NTplcbyVSGHLcOaZFZwa154B
peOeKKyN6fXkHr7+a8c1ebVZksiu7rjnZaH98qBxCFgHVlyYknqHqfIpFkPWNv5D
qHXZQHWbbEz2tg4dvM3PNNpzxiX97PXABD1mH84hYm1hFxk3edENFGGGMu7j3dEh
9b66C3ftk0NWuHM17JaTdD0RGTUk2GLG2Vh56zBPWTKHs2Gorg1Hqz5QhFyodMa8
KzKQ0BWu4vHqN7MHnBizZ7HD3G1MIvPW6zISA8x7w6QyZaTaoLQC4QIhNnxIJ18t
ngRUdWKXX+aNCJdaf//6j9XezefbLy+zwf6/WrTJxsG4N5Uu/fdxhMka++rD/e1M
t839khLyE5lAafx2sWgOnGxYzzmvWfZLVLCQBu5jtKk6s12Ss6Z1U4AjI8eAqpO+
Z+8quUNz7XECzugfKMd0Q+Wcdb/5A1Gcg4LZznhW/99fh24rFJQ09C0vWzQ7eShX
RDJu8i28cQMaJDlMpAImTb9dGTUJFn4ix1FB0eI2QO56SaNFyJqKQ0vbkvoFWVdt
03OCD19lluLLboFLHJYSLUo2fnCw0fZ2zSMUylN94JiZL92u6Avwt7d0uCQr/Cju
8lba/ju0nGWmJuYCdbgdKIbuKp2ih8WywPLfWsmGWh/gmev6mVtzaQ392akEGpWA
wdWcLEUWsMek23oejEiBFfYmgmkSeWLTgo6UKd6x+JtFv/Z4413yOfqR7IwibqZq
d7tJNqtgWlavh4fk6HXoXv824UZz6FECShAtlbqpDu0ScVysOqvbNp37YHi7DSv/
63HI2Y0aJOwcjnB71Vzh2LbDvmkZ7ZfrE5UAIVx4RGpt6TgdOJJwqXt/SdSys2OG
zN8G8IMyoayCSsbfGAWPsiWoLFHRY0Df4urwB4JYBAFZzI7TubiI3I8yuIdFVRkD
950nHIOq3uvMIsy1Vc2d9/6I32HNhLS5S1sE37u3fxkriBJXmN2tZwr3w5fI2I/E
0KKTAShpqX3p7pLaXbzvp+UEAhNqcMOzAUMUH+xMsF6/Mb+PEstE2oj2uAomNHrg
bH5pcf9gqwCcYmJDtHWogkkeccLQRamEGUIwYNtcI1OAgxjWtLnD7Pda5vK3+GQo
a7XnED5g95ffDjcaS+9M7HLJp+/+k2ctfccOToYk8UyYTMySSZzea2Kb+R6DEPPE
XlbDubO1vIS701S6Ia6ZJviSzqnTT/EPAAq1LASiHhYNmivBPMl91boLTyOKAqrl
PrdCMHlvxDFdTSGIvoavL8MiXPZL4qtB5C17LNjGNCtbWZSGAlDwvWdVK4naz/N0
fiYd3A6vJkRbMU1kJQSRvtG/Hsi58a4OaiZGpvl0YOtsl98mj2gwuknaEOZwFHHC
viqVN/iDSUrQeDn9CKg7jlk+13H+bX1G6A9zF1Z2rS8dGUtxT+b1UBepWuLu9NlB
1+0zz1/QtP+knvvzkXf8apv83i1B89CTVqzmZPI+UU7Wxr7NTYi6oWiGEjGbqlEl
ZTcAVYrLsL07WPtiqxZ2XpItHAKr4vlw+3hSPIanWJpwBBx8K1SmML4+uvIvZKYl
s76RV9cBrrkJ5b+8WkVM8YOmh5UCjMCIEJsKcli9ILGt/+RacvmwBE6rX25B/20C
42nVjUwzhlFzWEVqz48oDLgYJQJtkP8Ivnr/apbur0qZAR/SPaMTz4+x+ELu+nxH
tjj+MdxPkONyW3R8jxmvWp7OZEbtuuTKQX0uz90yeG+q2upuTBtDfG9vcO6O0dPG
4jzAxQBeHtwTKBQYIqeNkDLj56LTKYCRIQCOXfCWQVOIXMtJbHPH5jWTU19AcOy1
oZz3ihmlBVWnJ2OyWa7bInj1V1eJlHXNVxBW2h8Ql6j1ahNYu3DNUiFQO32EFRtu
f/hOuvsrMTP5mMZL44YSAQG39+Q2PIn279ue2odIsFzEHmU3b+KQCIKbiBhCe85/
7oj7fy80BL6xMB55z552cwTFfZRAmDDHjh3uJRpAy/sNyckNt076Vvc3qsEiKBpo
u7W8ogxQkn1FRRXxBnovNNNKpqCvpL5rSfmwADP/00cdunVm7qo201ubz2+Zyt3K
voTdAQp/Voim/IuTuosJCC+sj1Eac5oXjVxuQdesG4XtAK5DCpOLUKd3vCt80Pzv
l5lnQ6tpe19wHhoK7mMXKu7DwekIN/+MZDtnPMQwldhTz3chDmhvPCKVZY1Px33B
PNzoAYOxc3i1ZRXZ6IAmP9wcr2H7YJWH0BvFIedF5xc4WCJH8HCrl0v9E1rUdM4n
wJULJjWAFFtA1htCcGdZE5leGGMaxa4s9eVN1q6dwMK3+IQFXSH30jymJ/Rd06KE
h2YwGWX1tJXvPdHdbtpQ4el9pF9WcbUPCFJ9hECdLFOJAwVs6d0FcyUt1w5Ih1DK
bCG4tWVb2RjxPgaJu4m9tHFz5toV61insJQrcniwEnPmKSht1buukxRcCCy1o6kb
b1I96oO2rKjUIBd+k6RhXX7gX+yW0AyomF7FKhJz5MLOVAbdps8xMIqypixY4EKX
hqWCMMwYw2oUT7DO2CTdFnW9z9P/21yyLB0baiEMLXL56mSraDKhncr21bUkM/C0
ONTCIGZtIjM7tExiMCj6qgh+Ub8qhns9cp4yBKxrfhG9kOyDd1BQBL5mjImU/Yhe
oawWPZ0M05yBt4pjnBGcpQVIxHQ8EvbYWMOCLkaK6XDyTMddTdOHE38i/HWKOh75
QCa8dXJzPIJT+UFePlYr2dm/dF3diyN7SD2PkKTp9yBbn7AMJs1vGacxDc59zAqm
+xlS+QYYtP7jnNN0ySwo2bHh8FloPiIaiogi0MY69aSY6fnlPwTAONn4yeOnRJ2o
/1x8iu/T1LZzlcRTi3gjxzhH8d/r/Wio9LAv2/wqIyGgnxMVxUU7IoO3hpoZZzhR
M8dTn8QX8UtcRAgcAIngJSjksvSzfii8pIdzFtgzRe9ewlYBzmh2ESrokfVzqsOm
ZK2lNe+OSG0QAvy5oJkoeRGz5hDVetvoZrVTR58q0jA/CmlFs+AjnHBWDjiXsw08
zfQHndiefgi22CiTl1joiWTGGsKyEGpK4QnR2KpBMeA0ylwhQcxO7nRN6gXw8o7H
f+3o6J1Do9cxxz7ZGwMligGG//2L5D5CNyP2eX+RDEyB43y4TqTYILCVfUtv6h50
HODZUzpevKnNc62zf5lIUHjMuWh1oSUU418/3Haje+uTFGurZKXdgSd+piq+iX/2
ulKAZeSqqry/CybGQM26k9ikqqDw3r5XPretg4rny+k8ioprRvHDjgPkIiLZ+i2j
u60l1cpYqi3LlP9tyLpa6n/v5t7XKnCaxRB3FgU0UuAa/Fns7c48NqNRwRTItvOL
Lzj+PwEc8PQdALjwRPJT9E2/s1JC4WWC3GvQUDLwXFX6n4DlEoyfivbCBfPVKDbX
L3Fjs9UBXmvUz3VmSiDdFq9KOM+4wMuzKFGvbrln1LrCxCpAUbgnH6GwN/5ZeE3I
323o2QMp/u2xeqvA3MnN5+fIAnaKhWFUJedwyTkdOFbdyt4DoB4WSJFU/satNFkm
IMiCxK2Agig8IVjbrvLxeUsI6kwp5Bfi+wOO2cc0kmRtlbazLivyw63ZFmACAkxo
oCmdVWhOkDpaqXwI1owqqlRnPpZjnGsLIi1fRX93KDR5HnhDink8+I2Az+xSZJfo
GW1foPVr/uxdOE15H5CVxLI8uVddh4iq4YIrj8uFYH9i+R7K6hOz8IBC/C1w7O6X
9GAWfX9U65lK3f0cdU7s5rgAN9eDfrJT+O0YSOqsEAKqiKlulH8Y4C13A5oei3dV
6uNck2uwHLGApnQ8WjubjpZnpcUal39sbGvESPlgj7T1+vDJEy+G64xJ8Q5bKZnt
NiGHSw7JBr7j4QS67ZZV+GVZxFeiPpEbEn3+Jmw9T8vpIZEI5Vkg9s0AM/8D+VWT
th/5SkXEN2e/VIPB5eZDpmwwU43fRPVlihoro6F0b2YHHQ+PYlZ/zH3QlnEikuQq
XmOfFM0HAKu4l8+4lyCVOkzosU73za6QAF1nBQoBaUQQNZ6mvMf2aHtzlp+0Vd3m
zkdLPr8tYkwPlv/+LeYIg97VJml1jc64N62bYmaaaVACRyP0mAnT7Qp7IrDw3ssO
i5kU17Bb7X+CpruwjCelif0B8EiopfvUy+lzqSNOCwaqhyG4RwtWeYCIjAL8N0uQ
xPRQN/Ea9od13kHYbdd0L7DFzXKpR8/QplnVflcRPemvf25+IiG8Hjo7N1l2FhHm
ltVyRvDvnFVeNuqKH8AQHQ2zbLEHZFTHfJQv1cOI005TrZDkfOmKQIzOP0lJrgJW
jvUnRlYaBWw7jEC+nADZVsEVh66QUqKQgGotLZ3vc3DNisRr/zErypfVRFqP1g/8
zd8DNrWOPXiSOWTaWb6MFqvSpBwnMzOczOI8wdQENXIOgnsV9SrKnDqeIpPxpG1u
2uzSxVttt0xnFsn8KJQQ7dgW+QqHO6sj4gObtX2v05vKT1HKNM3376TAd0Ahaws8
gQnv4Qw29Tp9Dykuk3aBMKJjLns2PmIqckRXmgaCIzbQDuoTv30aODc6F/WKtfsr
GpRH1B4CVFZZJn/FiEXPk0yxMf7CROMRhJE6ydxLGt3Ivh4crDYwkhPfhmSunVp9
KsckB1ELbJI75njaUXgmVvOdxwz8lDZX8biIUZrn+EcA0haWK4q+TUKqpzq/3MjX
YotjfdvgBGC2iXQW/+IDPkm2KRBw9Bg61buIdWj+edE1FnkScZvOWOKRnhL1J/UJ
hEPgmjBN9q2zKFuMXZLwvU5qVKWYNhPS6sv9tvG/0MEzjSR4/YoO+w1VObXMFSHi
+BwMgANv1mxUTTM2hI8ve65nDrW8gOYljDKqR0AQtPfzlq/5EC8g3BX5c9XD1sQy
effmDmqNNd39BmQAAusooT2fadihwYPsATMTuLOh/gNa8IIViTy//KGNKBuRYxWg
wGFB+S6YH0Tj49i5vCY/z9WusMT99anb3hsB6dD1ow1WbetqBWSbBK4X6WZV/Opv
nLYf6/Yh0PJ41MFtyl1MB9zhVFH2lUlNBFEgZPTefLhrup8JRz8dJPVPjONVNKBQ
AT7YnQMzY4BFbs+gx7fOzDPywzVcTAN/AvaeXjmnkHfyWDRrsxxxPZTI2naUGId9
88hZUijdmlPMVYAYmHQ+giGxUFW76sjba22KkNPSdWyIzoPUh/x5RkhTkGWIrVfi
sDwQf1LDtabakfa+0YOl8rCf4vnivackqW5fuh9C1F9rbmfETGBANUOK28zlMjUo
PHeLzgg69vZt6cnZZAxYZii8e5JP29B16ir9suIueWEMA/+tO8nOAsY7248ea+7C
LiA//3+KXRgPS5qf48zQi0ZUVtEPhNJT/VEBuiJww6EWUVwF50WawVyIWTXSmToF
wMaC5jaVTXgkta0pCattNfgjsxMxPn5pnIz45tvYIA6c3NVqhEjLytOikKZK9nMC
cljMbZwl0+0o0u43KkE3FkiYDEHTF9aX7wTWfZsxQ5+52PXt/XDmbTb4kqBUw4rA
LgEEPJKVHgODdIihajEny5V8IhukZZgIJf71d2X/Q6OW7R1NJPYTOLIJQngE+BL3
cNYTCAI/RgDY9WbtzbASD57oUV2AQLHhBupD5hsVWH6HjM7IhSdmB3p/TrdMBS3Q
PGAtKefoFKmcsz2ZvRK/CswFYAVs80+zWziaQktbZweZ3c8KE5pmw5D6ZDxytdD9
1XCRZANM5h8i7E57EbUS5wFtECPcxrPUPLKqMibvhzjSGq3b6De4B3PTVORuiylQ
xV1nxUd+BYu1NYtLMnubsI+Y57PN8qtJ5RVR/pk6+ngRWqpMiJQJ5HrmGJf/r/D8
tIgdT+YxgU1s1S4+qSEa401FBNAVDwZluM+vb9dLBbGfwp6I3LBV5nbB2iKF7+H/
8sfIWhF/INKbo4Io4RBXWAh4AQEnUdo6hxlYmzUlGRohgXFpqiV5dPEXFu7Zle10
QppNyvFlf0RbFc4jkRihggBcltl01qjxzCpc4C9KuBtmG/rwkFfiesBESnpOPLdo
aSyKOYDQgtjQNMRXOoKiFWJmBQ8dyk94TNxcvBC9NMsXCdICt0VAH6uCsK8pq8Fs
VPJYtOKniu+sWlTThmi8DaI/n3itHNRfPszBdyekkFGJxr4FuZJaIcMXpwcCwytX
wKJ8gyeptNikZ4j2oebnDbNUc6Gq5usmZjb/8rUbUHVPe2J1r2RmvKEas7eo11+o
RPm4t00M+PH/ibmNnRwua0prrFlTlQ/7lyRm2tauWS8Cnmj6TVJ98xC0mZZKbDME
zTamqZYuKtTwDLckBA3BvRnnJuG40MByJnzNTPLcFydf2Ja8HCMu+NWPa1arE7hQ
jjLnUqnuS42n/oMvI0eFDprczfQw3+/5Fer4R9nE8uBbJFGyGkB6Rw1BbIrH7F32
6IC9dzP9YFtjJOqZYeKM9+fiEz8CZTueEVoZQsD5yoJnP/uGdtMuY1oDn/Z13VKK
R4fepDIIaJrF6nYSdYpYRH91ctq1LJbXRalwryapU6jrHBW/5onDGd1BCCI2Zrsf
EiXfXveZYhiRT+bw7cZlQ7UJlsCJ5eOaga8c1fn/hXWmUlwA3e/7ORWhm5Posl+F
yJUMz/d+7w+23p9AGxv+L+K6yNiskCYcyg/A5Tf7V57aT6msTsAN0T8EIs+IavWp
YMwpN84GoV+h/2qOVrub7LMVtmB5FOTgznwfDjEL2iCFSz8vp3QwAxlTwFlWZcvH
x8k7cijxWTPe0nmP8YU4Mgb8znPKFYJLtRL7IJhzJQ6HnAKqZLc8BRgk26Hk75ha
d9DFPpk3kf1zo8zuMSKoVTb9qhb6893WT7nGOWyGLo0GjjO9J+1ApvTChVPOJIbV
krkPdU94P51rW7XpqQwsjOlLlOzX0xcgeC9S/kMsMY0NAC9O9hUKwABCCQFCzgYC
F/VdemyZ5e2MCDdDxmwMcVc3uvHf/gqhqAxer0yEzp3uOlzdiJ2FbkqQowjpC3+I
zpobgVTRGIa/F9c8sn6aimgstcFi9pcOmrfREubfbazxrdJaMZobzlAvEbts3398
3JOv12xE2QhjnuV6zBtRCqk4Doz9JFsSF4CxJVbBXOPmBaDmFYb/GSd+JF2lIhQy
HRLN8oGc0vr3FRmChKMcBz9FhnOgXqyS4cU0YMN/8GHLYYO97JJlAVLK0VSTmOMg
O0GkOWr8ftF3SW0Ey2t16iqzA6acXdL40w2hKyzGxmGuEi4snFTF1vJPwRbzw6nH
MRo9ouQVFtzidwBaLwJjAoEni+X+yrIQVYu3SwJ8c+qX7D3nB/Q0fasg5cSZ7r+p
pmpM5D7GRovpJ7MHH8qEqXiub3XJvO1GPFI7JBh2dJ/VgWdUoC3VkNq6lbXP3Uor
gBWN58DPqqtghgU+Cl5lm3UufGoSn01wIPebkLpI5SYpGIxS60kKrcwXv45rdJfI
0iXN1jNm8z2XMDXloUTwQwN/XaQO8mSMNOQqEheY4LOUB0dbypmrqt6bGk91SABp
OZYJmT4G0H1RiFwSm0V5fdtPAEbn55R3kZbcCQ1UNhby/q+am6LhpN5ww9lbPXUB
VTPUDBR+ZQ8uSSvVN1jkqm7XrD7VBJ7AQ2Kpft2wCpqj9FNPhupf7fj0Fu5jXt3s
paOR02fOuNRr8m/8hk+IVXj1l/5BbSHmEocamFBkyyNus3S0qmSqyV+JNA4nDIuB
fNdjIAlTej9xjReSJfV8/L1KeU+JJM14mBjJl1IDzbLBL4ZJMCIzv4PytxieCIz7
BdskbboSnJqGdOeAxZBD5/Nv5y0lKsCcA1XsK4de1a47BdF2mlTJfQIKJ1VqjWTv
j5Fp8bzersMai39juZxzuln3IPMH1OtVkC4dQRXrwqRVPvrj76jKhkhu2nbrDI0i
+eMg+SsndyXyRdJnAt1WQm9WJXsJTgN+oKcMxt7snkf9hRbQKOdTFMgV7Xo6/14E
hlhRDmfJ5RXAnqiWC/ij24aZALUn6Mq2NCCzFaTIErlV3yOrgCntJm5Z5uXQoVro
zM6a4CUnMvqvW8A8cIhaAXDTUY0SOs5KKa8jC2YvSoX+RMLT4gwVUCbCPfJ6W1xr
h+JWKrxcWAHBO3hPpy+Rt4oPjga0EgNtnp8wD0wFnFnk7sEwqmO7tEckSH+VuXa5
Cvv9ndgrTv77PDu762UORYichPN/esGRwnnqHl0xe0ucIVPKyuengstjLp0g2fm5
eAqJvsRDgOLihpYr1y9BYiAPJqvUwxdZFBOX7I/ErbmQvSvnb1SMZqsVi+gwwmCm
zsUwG4z5eLpVQVCbxJVAW6IK1V+VzUGTFsrL3MrBXwiuW/+FAx7VUAv+S/Ojt7kt
97OcZZJeZavtNLhyP1P7SgcXj2gdUQDAHDgKREsIKaYbhxUzLuO2rS2CW/wSPf28
LSBn6CC5wnnuB5i4ZlH/A5frCi/fvK0oOOp1SxVIf9VOgFfRLR7aoMuNxrdLEMzt
lKOu3d/04Zt7EqISj/6rBwQMhtFrD0M8L13NKD4UP9JACz8h+hdyKsFgll8cS7Vs
hJvBkjyO7Grcfl/0E3Fl9P8xLwiIiwfLJn6J+mRByiSyxqQWB5KnOqRibJp2VZ4t
nbI7CTauAE/omtaXu/3iA9xI2PM0RBcnaTULuT2vgYDJiEIa2JKZTOeVWiBJ5bz5
cNo0ebtMGsQpcm2+5aaX8Qv9DiOovzL5z+k9BR/nTS3wAfm5wu2t98yAwAylseM0
1fgSmxKJnVnQS5bo6z+cC/kYlB1rItljDXY+lSKE0nB1OfcerzuXTl6GzJnblQHy
fY6pVQRCh+a/Rn0I8CWfKhAmxyP3yMfkZAvonpYYzzhRxuT/M9bKCEmo+mXC8kbw
3P2O8pJiXQJWES712VaQEJgKVhUiQdcSvfPVxSS/iF5A3HaH+DW8Q9cjE/JYm7Td
OZ7opkaDCY0r3FlPL9oZR41figC6TmhHhnokoKdOkcoA+6s2gRbHWU2I04SuSX/Z
7Mt0MsIa/PST6rSrCrbiJWmAQMviJVav+IcWmuij+7nhhTnzwi3HOW7pnxdEt2St
2ODo04nT7qFOTJupr4x4PlbepQP/bW/mAdvWGXpjG15lw2ouOwBaRMJsbGVhaCuy
Jvf+bPn4YI4syAIF64xXBSrskUFQeCXZmCKlY9OsUOrgAaBWOKizwQLe5IzzLVjz
aq93pbqVwTwD/HN2a/tdWlRC0enQZdcdfciDRF7s2xqNKzhakVXaJ3LokOZl9i0D
lpFKBZ9s8TJ9c2jgVxqusWio6JP8Ctajo5azRSagAbqXZ6vrdmu0r0vpAW5dxZhz
qUEKvwbDGh/vSJjy00ZYDPYqv/ePJ3LEij5LiipM9luCYieQ6ceIILpE0m5K3sjk
lKNAWz6E6MshPsgGHfNZXkZBGvVQre2i9jTIE4zTorD2w55whGToEJqoaEU4u/Kk
mF4QE5xn65mecPJkf1tPXfhikXHYwOYD7JzaI4vyQERVvD8BgJeuBBJlTUrgG9Mt
yLVzeYxw7ih5HwP1hDin1xtLyTBKrWwE/Htg9hftm0gSehai7667eM9tFqh90ctt
XP8zB3jqO97ZYh+cgkiyGQ/7FZu7/7pFU20wKemJzHsUSQBPfsA2oPSlU5ItCQm1
Go2Ytj0LRbNdGEgK6u2+9pL4raAvMjvdoBrCNs2WRtbXX1hWTNkZT657NMNCg8n3
sGXPQ5FlXYygTbnPup/OQl5jvrXeEOtFYmW1No91RG7C7TsKaeTP9w4EQrY9xGxj
WRaJZSe1RaVgf5//Cf8ZLJU9VRc/C3UGslWqOB/je8W+IZ9jR4q8aIa2dbG3kPaV
Fwxn09uddegUV8V+V+YmXV0rVio/71GiwHpxfAGtNd1KGrqYOKojZ+uOK5th71Vx
lsL3vRPdmFGU3/Acg5zxcDxLNyyRo0kLJ963ndRlq9l29REiWWjsrfHDgsO+3LKg
0tnIwUvI4TwsP1SxwsYuHvd5CvYdhjSynowLe14Md9nJamDZmmnDxx8sh80ETLLh
i9kPY6ivUsNnV9tcCmpZGommZtRzCobnShp92efQRt4p4jn3dTkIJP/S5tzHzpWX
iNjBaf6HY5UY9IXoYF6qmuHDZjM6PkeP61P8BzWpOi+Kvap0kQr1idU6mmQf6zxI
xxZFWgisgM0ZllN9s7dvym2RiOak+h681ep0syPp2HkTiKy06EBRlxGVqAvVl/2K
bwhoV3KyzIeFMHGwaa0Y38gnkY2J/R/osyFm+3bp3OquoGiJcWL5LMWJOI1w8SKK
iVseXJkzYMouVQfLZpkh4Vj/XCFsfIbn0dBJL6azOoEyoFlz7ZGrzS06vODI9wqK
fnInBntmqDuLCjJ5L9+4WR9YC3S4Ta9i5ySlSwGMi3ghfn/AeLYbnVprTFHldLS5
+uzEKi4JLSNQmIkjmbagiUNOhmU+hOqYarI0ONcG7RwDdoW9nvEwMaWe1WZghEpz
M9CkNgeGFnTnYeBeC+VIjMXZUxjrExy4Rsj1kDGaYbzpkHcnr/4AREVsSlyaQ9U3
8Y0iZXqItqo+u77WW5gb/m+n2R31Prp+Y761drH/eYJOLDa1/aMSy7wWSgv4veqJ
dmht7qtgMP9CxNsZ0OP/JnutwsV75V/xkAjKW+pnPAGiDaP8toI70YHuojDnFhf/
AmkAVEktwui1r+dg+pk4RBA7mh98G58pcjQzUiWUUzmFEK0xhH/NYR26Xn4c6Auk
iyOO8EohBncqIciGTs0KzntuKDpiRyZc3YlJdMTfgwQfXSlt4znUwGyI7/TQ1y+i
1RvDnRTU78gwBQw2kTDbQ/24OitycE564sScnWyZKi91m2FtCcIANqMj6y3liDV3
58rQH60Zj8hwNjX8hqFMnioRJEsX/vI3bdaCIiOudUgf7WOsuL3wigRd9bz4104J
8spENxjwwqx+KVhRf26btv598/TR9P1aiUduH2kS3q3dhzixjJB5Z+0XDMKghy+O
f34fc1QfVZ6pRbYob1kJYrqfH9lKS81myogCSqo4u9oOmo1mSUYrci29U6wWI+qR
RLsF9AhMw2RdSD7BKbDQMN3pWw8MHaQgy+MaYT6cISITmFdxPMMFsHmE7ePukBGy
PEMwGbxLsRxFf5c0UGSAg+DpYOa7QKtr5Wnrc/v6uUZMxbKsdS7b4rM2KAXaqWJW
C6UxtPKY3Wsn1D+XW7Tw5bRKjTzIrwpDVIRTtwFFYf3V5GDefFbHInbjFKLiD5wD
Hc9bHFeQ3RQsd3JBJrpi3+ZZjaPg3xjVUOEBBS+ZlD2ggJvTlXqvYOQbFtoYZAH4
AF3ulZUCO3kZ5eB0pQF8ifPgZ/k8+vCy6gno1q9ONNpoQaLhZOvQ0HdbfXjxU+T/
22nuepna2mUi+ij42RLEWdRQ8pqSieLsWPdTT+ggQgk/W2IFiy3V3Z4bqfCYo9u9
lt/BDkOWa6HAdpxvVO+jOgjlg8JnKKl28oD2Ni78r5rtiSlZbamBtUjsMvWLNdDt
kHDY4zcDU1rX6Arnzja2h2k2ROCoLjZLHnmK0jUOWyNG7B8hybcL2NBWJetGEtPN
SKSrKqjb+Biht8j0lUKXe9enINJ9xUNs5g+/N0lDrVb0Q/8JxTqrYjsbsTvwEYZM
pot4H3vbrRmV+T2YelL0sTt8N4rfsjKkiNlT8Wq1PlpyGYNekdOOyt9rVGi/327E
YG1VBCcCd9BsXuaWBd/ewRsxD4GFAA4A0yid0AexrPpwFstV/U9FIWygpKydDOD4
FoC4d6xDX+qWSIGY7CJvIgK1KsHPIaSJKoutfN561oNPZJZBb8z2lpSvys1keLP1
erIT3mhTdvOHINZvloyCj/bNil+Z+GAVM3IyfI1yQ7SJmRnRCO/5pEz4tsB+pYCy
rWwd0Ds+bhxJDe+DHK8AgkH6+IBWR4q6x3S9u7poQUIOc+qE2pDxE6m42rV7/zEM
NLAXitLtHO2UOWaB0mWUPwk8WrEIMXaf8ckTQF31SocAo3Bl0jyJRwWDXfb2Q6qr
GcmyNmtgbP6aew8zXnCdsuLMxTTh+uwzY6m5Y9a9T9HgQHPpDQ0K8SP4s+HEFVRL
7CG+KMOQsRNZ68yp4BBPu2VxlO4hbRPoNR/o9kxtxrVqmttrLRYO+ZxtYWMh+nZ3
N3U5uuA6W4TC0fyVdJYGg07Rdh+HykNSFksP1bIKMhnybRUc0I2Odun21MnQ2t51
7OPhqmo3qWKg6b9yNTsvqP8OnS95NDwK1ZVmtJqIfzFF10PCWPNrHr3j3gqjKNQl
3+/R3uG2BfUWC1kCNSG5p4sAsKn6kTKSRZgR5DjEYnQ6QhshTJuh7bwGo7XlE9rt
sLmHuBLLriuaozjXBe1TI6C0umCDs0/w0j7WLeAnLJ/sTr8RMiVO+TW8A/60oD/N
Pynadmw718M5dBjkzETmllqENQig1l4fxHj5axBC9ffqpkalNI6evpckl1dp5l/R
vWUW0IvqD0Kyl8i5zKaJS0Ckx8hYPpgrCERBC08jAj3PWQr6MOH9DkEIjUuDkD2Q
`protect END_PROTECTED

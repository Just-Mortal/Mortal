`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jG3CJ4DeOBeQtnS5sYJH0xuAeIMPfBkS7gBNbx3wl1IDbhTlCgEpAoeWY5TBGZjp
wE+JrFZJCHqj1js+DYAjFRaWnFGxaOCfY/Bx/rmMct1F453hjhylXLsECFfFXABR
Zx8u/eOIWUg8hsRsVM/Dc7f5diAAI/A5TNE33sdM/hs5/GaTR9jj//ruMxA4Nq9O
uuSLOvGpDW05hZMMuB+b8piyR90G7mHeQmjCgLLAb6gDRhMbA02hBBXC+FlbteNf
wa2P+eydjZjQGAqG8Xfkw6ytDmbwLHdD3nOb5GJYt5WGLmJ5pXhcEYRfN2vpTele
XhLNF2jYk7ur835MADC4TRPywe12JYKbgLmPgA3rCdQkX+7h0FVLPfIYD2OXZCnB
gibAnX8VSvXwRL/+T2EQnUtTA9KMSoKXHAi1JDQRDzu2tSt+Qz1w6xVKZoiSo4zo
H0BU5iJe1hvolBDSnnokW203K1QK6Ck5vw9LDTfKCRN/FFYARyoUicYVGePyCRpz
hIt8Yn30hak/II8yHqTL1DyOGFyvlZeCe73STo59mSXJQ7I1YN45U+81eO8fo7ff
3s3VqLTLx9RGYLLHgvSc+5gjvnhf9He4JwnTJ86IsHGuPTh5gU7tQkPJUcH7+B57
xU9q6hBO8A6o7nyY7gbXNV193E41zc/Ey+4Yc9mXIElTC5u0tUusLC4/ddVMKi7J
/tGTgIStC8+LSyTktpn7ukYjCE/ujUWhm6c40Svse/cAnuxwjRSv3e/6WY0Cjcr+
4UnztnvlD/MwlBnnmcQd4fD1n7UjZMlLGZFJD0e6RGCMAWU3YzCR1ACA9GhQlmc5
f7kgqEySqJ+jzuA6OxvifiiMtuSCAl/SttEwuX2oM1z7y3pR20VenEIc8TTCbuD7
ptuGLfiotJzJRplm+QpFx6Sp5We+hoLdeUMiIHU1MYocstQUBCk8Y3cvzqQ61fXu
HC56aS6z6CTwMVlELndwccXbuF27hl9e0ENrKzTL/Fnc9jBpdgNUrbf3JnQeYXUv
dFffcw9xOPdIE1gOx8FT8QiX7sMPYNj2hCaZ6zFHZGlJ1nYwyt0LkHbU5nzVAFK5
CQCDd/9wrBbs5ciHN6Oasv2olCDSy2LfOj21SGAPV8rYZWHLS9t8mmrlAvyt7GLq
+NUuSVdRbuVo1qtInDGxZDmQMFW3zfvXLIyaiorBNvnaS4pmscCUA1nJqqyqLzbh
fTg5DJtk7RpuFmirkPh6F0oq+K+r1UJDZGkyTQwXQvLFGBCXB6+AIlyxi9x898Oh
G6aZQJlCjKMEog1T5RZVmgyAXud5qHb72SGglvq5na0h+fwUMu/HG0YmFzGIRnJ5
snA3/5oWgyJSWPbviiF0t2z7cRTSY+j986BKYjzVTv6Le161zmJ23OepDbHrsBeA
R7qyIxv2NUlw4xIMPTLBmnSUhRGRDNnCe0P1RoHKCmkguo3GeFUiTbg/23XRu1z7
Rlbp5k22oGp6pXjCb2zG7SEVPQCK7ldLf4ziwyGCuulHbBiC8WrqqiPyC0Snh3KS
qzGXJp4Q385e/YaWrIyqEJtGqiFA8ExvfCmEoNSljysmpk1e4Y7GzFQELTksRSvN
ksbuaZUduDknd5H93yzDjNw3dv6UzTjE4LuAl858Its=
`protect END_PROTECTED

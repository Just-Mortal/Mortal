`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ncmGhE4qJJy08MkvenFDkuCokXOeQLHx1M2QNaDL+vl1J8Ugp+bvksfvbPze+kD
SCtstMOBwj7tSClEnswhvLcH5p0Yl9z50WH6BZHpFt7ZcxnN7RxMq34V2LeR8N33
y7mVyHiFYakPPm1TTOSp/NS9R7ZFF2x5kKtWW+zqE1odIf6ru5tuonXi/H2mSN+Q
AFYCUodqGXoJ1bZLsqyqvHArRXG8sW0A9L8e0Uxq3Wit1Or4Wi5FxAI+rghiTLRZ
UKY4XsI5TDnHzcGSKMQQMN80dzBugt3aB0/hAFjOjRx1/XLAtTmXBwWF4Dsj88Oo
Ir5bkQmBKU6idF5MtOXAY7vlEwCMkVst7CU5uD2muAt/V461o/9KJNS6MYzbk27w
4XZdmPEsniQ8QFfFIJZTIU3RJAL9+hkt5oLt88fWF4FiboKOGX6VgOGO+6qegaUS
kQxBbZex5HGZG1jEykNRbzDRHxW1zgmrbujcdn4G5oOxOp0CcJw+nlBDajxYJIhF
c+PyAmWlZGy34xtIwRWiXdTdqI/waZuKszPjSicpTT9ok9pPw9fi1D4sO6sGllID
Isau3rIJgN5IbopgV4fpYYImzRtUzMiTNO5pOfpqHJykNT0rFNlF+K88NpVHyLTt
9mBq53GNTvTFHaf2FN4yLfYg0MTyi7aNQnIpS4slj5xuBRa9d+rgbGcOLE7V8qN1
+d670bPZ6EcXVg1hJZ7xTdAeaMVKmvciZnYtujjPr1AYVZ23G+DCA3FzSQ70RvyY
dTBosbGfXVEJvFyBIM1uPnwlWCV4vPEHxJOBqA5Frn/lut812c4yINhFpxW3HFpt
vgCn90TfgA67yO21YvWZNtSO7vVWj5HASmW6OTSdUmxTw0ROnw66LmRt0O6k4lQM
DuwflYkaOLYZZ05EyRefhUwwUkgRlnnPWrB/WubygvuYirRIFfKyHAL/vB73CmrI
7CJ6G1lQ9PGjxv0xtaDyEk1onc4sSAMalPMt9NjOxttYVLzoFIfoJhRZ8Nn9uWjA
zTj6ULrNjKe/J80e3A2RwapXVgJs+qowDpg6+9pMetM3KjsZ6upJYU9Z8MQLet7j
bbfMyGs9S3HYEwegHla3GCVdIGqm6Bv4+AytCYKgvUUcOgNQPUCeV9I8OzT9UK/Y
cxIEgZQAsLFhj1r2Uoviu5oITLJ3ieMalwnSUgBwt8ARvF24pCaPreAfxVZ3PYxh
0DBWH8TbN4+r5qZjhB+5DOT2tLPkbC2oDI0WUMI8QCEEcwaPdE22PXc0bnKLTEHB
jmRIyyCKtvtynljwiOmi4mYnwXQ10UjhUIu6IWVFpPTUZV3PpZuho3FA2+XRel3S
g+LK0ITTM5Pc/umVXNaUcywYxMXAV5ubMju5+XHqgad+UFnlSBTP/7ZmRX8Jc3ta
Eb3IeUijSWtph+dCrpSr+S19vwNvcMf7u2xHmZyBqpjWxlGJfFT+9WaSSSAipJ4D
aKcqvMqYQQRXXoVsXI2GUcRwkgFw5bcJeHDXW7e/gNfJFOLWLkWMd4W75JEXO9mY
neey0nEPi5DPRVhVcEiBeG5r5kIVZ1oKrYpCt6G27pNFspeIWpLLpJksskbR669x
D+gXMNeeccH+f4wJN1+vaqOS4xAJFxUXkL0vbU25n8AmrFsU6FVp2rX82yYvjbaW
/ucQBiXz21Zp+uiphzvcBvacXBfu+JOO3Zp0duhgxRaP1V3bj3/F/dmk2ldXEaug
aG09r4Lp5CEJF5MufYgtk+u96Mer4IZmdn6RNdyWNwGZm1JQ6hWqqsTwNsGli6ze
i3sztbQC8sJCsi/nnFzB8CmWmA1DP2zHE50mGqpJu3aaeRRRqVoz0U0b5fUJ/4fv
tzvHwm2ZsAjoKcRjM7mnVbOaIAirS7vowv5pjqoLe2YGegnG1pqaLmCR2R5slAhm
7hst+ifNd0x1PNMig/aj3/w/8U6eQPxgy5LzMpOshmAsgr/w6HLidh8haZJrxUnJ
HET98LOB+eO1QoEL4SFtraQNPYPIByUcjgABbiHvkB3tAc8NXyYxVoe0WtchqLPF
Od1TjaRyKPSGiYW7XwROkVt2n7u5FrOpb3i4bT7+KhfDgH8EmxYwM02YBwHwY1iH
2zkemu8wYATKb0Ju7Abvei0uFPwNYDplk+HjcT3zZcHe1v6zrlfstPFpnVUZ0IWD
F/4YLpimA6ncBD5Bvq7fU6YSUeHG/K6IWPNiU7ynBo9JO5TSKUk4pzqVONj+bmW3
r7RMh1872ZsVq9fEGx804GHP6ShygYyg/26IWIiPTTGAbKJvSFZARwf06GcxNsac
AJYUvBtgTwzFHr277B/SG3kBPNNXRegAJl1L2ooU9k49tsMv6zko8DMjRD7qET68
naF4a+GfCD38o9RsqUTFj6JN566TaGbc03g+NF3eIGg=
`protect END_PROTECTED

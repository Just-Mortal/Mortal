`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgxNn33T8J+Gm+A4zhkoEFqM0GPoH4C/fDRcvcB5Hk1lF1LRGuH8f/LDDJmW6HLI
xhNyYWlRT06Q9RI3wBUp/QjRetTA8R4lVk1VCazgGUUaXck6PtWrIBn7x/q5XbrU
m+cLU9xedYqg4B6evaY4OmJer8laOqwmTQ6MIKyUFczBroY396VYKoAM7DWGePLG
HeJKFgYDyI7PuIsUBnZos9av5gHmq7dTKRWv/N3lTD69clhltONBQbzapCzPsq/L
wHPptIGsRFXrz5TCUxFFrpFEJQcUVQfT5T6qTHhhhVpsB7s+jnloA3l7Hu6c1fYU
6nOeqnTMKXLonpua3R6Gi4Kv5P+atLW48DIhrRaBnPAVcn3YzFWp23shr9iLQkaq
Sr9gP/0BwzBCtqkpPjpWvTr9kVtYHeUOkiiOwOLO1J4S/WWla/5zKkvRXRWtuqVD
6FF3CFWshzI/wJO/2qxh8iAAo8i1o+E01IGpgoruhTg2bwiArlPHwtPX66dnv4vR
LP/eVq97Vqf2N97kPnH552pjJ7db+T4C7UZDU5SpVKSH5Rsmc5NHbw3EV0rUaZig
35jNE/39gqF47gJhajdMvsFsCvgqX2wV0RJ+/8otPaLWCuMj6HLzT35wMIOHm0vD
asyBXB0rwYQgLUsKpXq7TSENBdOYGzeTcsVkug6dMgzy3Q8urK4KUDpAJMq1aLlF
beaVVN1C8JB1UrjutxFEnpNOK2uNVctFo7HWxJBwUJc552gO4CFRN827tODirmoC
sPg4ZjNXf+jypBvSpx5nLYoE+RJii+pXR79qj3JUWG4aDG/4LulVnpqOXQHd9ym2
RFmZWNiWlZyY/OCQs/1Rt8ZN2VYg/fqVW/VLQvlk0KhCqG5HOEPY+R4nhoo5NFNE
uk9bq1wYNzFsxgN3JLZ6uC/Q5Ph+/7+0FrIMkN04kMh6A4x1+RZAthLQ+GKsAbHA
/XwhtMx7uWreOoqFM6+1qCN4pPcAl0bX2hIqwR08MGUjRyrzoaEUZkNvUKNlMwHJ
Gfjpv11SSxq8EACeu47CHlN/qxhX5q3Ut8fppoQKyC0h//+saZ2AfjvNKipQPaco
pRlA43+A5kPx7C+oPzdwzDCCmzdDUOLDIu8nzsTQM1kXf6dgaoWvMYMjisLdUyVL
U5XwRS6MBTwwxIgA89g6Illr7BPm6pcEZR4wbILHBnjCLVMS1t/kDhB6o5M0rIdG
m7GUBPmHUcLbtPOMjQjn4F5oC1afYMTvwRV8Ylr0HFUf445j9nLuaGcPCVpFlXP3
hc/Or8nxt1xHgLPmxOESinUsr2iBkpUrY/1BigS8FY4brjiofv2pUdoeljkBYJW+
kf55P8FkKcqE7MfqzilBD+NCm0/gtzGiR3T5AYjBVJKEeImSCRtBu4nowj2Odjjk
CYEO5sCUo5yXgXPz8DsgiJK8vaRKpYjNgSfUO9XkeE8kB6zbZqNV0n65nFbIIhdK
LpgW+0FZUM18gGqEcPENRdpZP+d66v93YU7lWxl1+iVo4YrXLUIJmia8Fr2wErQ1
pVPd/2v1Fv7MqV3e8W4cX4CYql9WL9l7vJAsyOK99mBde+va9SftUq4mhWCSIJtV
ffcV+ILEXdinlSteeu/GtOGtSyQwB6qbvifUkD/vqsBQkiVR0iEb0CgHw+Qwe5iT
6HnFex/TpaHUSuJuroRBO2Wt3ZZG/X5Qt5ZMt9diG/SkOf0c7uCFY/L7iMZyP+SS
QdFa4mzpmAVE4a3ipEFduqJhWR721C3EBvyloOZtRRP2cXVg28u9b3OMQkE8QSrW
EpHMDgC3q3bqx9/iOXBXNihuKEsgzYWYJ8UfONMSahmJyGIsLPrPs4DjrdZ+/mhV
GpSCcm+UlQoi9QI1MiXWKs9udRYpCqP59m2nO7Qov+39JBSoMVAFOJRHGPo1NZEy
spzWNw1OXwZxbOeal+kQCsSHHc+jO7cuTQOMv6I52kH2ENFoqkYJgnRFLHcBg8T5
md4HmMWjWG+tTC/8rBjYbh2U4Dd/rNzhce1OETTWIzuQWhmONGQocwEQcogr9Os1
pS3b5oF8hvFsO8V3mgbpxSIbi97D2G2tdZcQb5Nxw8EQFFiYlqwp0fk6RQG/SqJm
tG2uFbo9rLLM+gceTHiCBG4XMRtywPjwkmk9z1x9BL4ZKPRVoaMJ4H0PCJ7Na/pP
AYrYACOJdUYTbdNJdQQnVDxUCWFsUOpytxg4eKS+BvJCK8/k4lJJeuWuTZkxfwXB
yWvjF3u2pxYYsi9yTdVTVNkiYV87UBRC8pR+S+HuxXlk5UhkaOU50Wcs6o+wpuXl
raI8hCi076BH8Np0UzfjWUU6hSCjqWa7535OKsMZV0+C14pQ4BWPvIMSwFsoF3bk
NfEU6v8vsjiOwp608tCp3fE0/npKyrM6PqIF2jJteYdbwhW+sTlwiyfI1CdeaLln
rb5/DeW/0H5Z0Xnkj4eBS75IOlpI7zS3aODXsIt5C3OIs3yhn+oS6QxrK20FxeeP
I7wiQFjg5U0CieK6ujH7gnzwcQXcUqCGXigCIIugJl/74qHtHGpefJkyvgk2KUk5
RrtboiDwzCBQICVj0HmGuE8B4VJvYR4gmlkUiiR/jIiFwEePMtuui/sEdP+W8oRL
paFE7r0G2/cWgyJMJ8106LUE/3N5Bknghaqxl/BnjpAogOt403j9mhnT94Tj8KfL
e6AzA0iSOzXuCA81lSOxgWB91HwA+7itmiBLO8uLLO6dC6BI8BDsdnQq72n6kPrc
1orLajOr7YPRPBAEu7m+pAGnqK90SenZKRhTHXMq/Z+/yupMSyHuGIrONhaUHPTt
E1Fw3m2Q0J+RJT6gTRZu/GBuqEaFz5G69JPISqbhRYqpvboxwzb/RkdtKD6FpFa0
di+7ydaZPjJtKLDxsLsHoDITqzDAIbJD3NPF9ylCnT7siBbnFlb1rmAfj5J1NYhG
qyW+IKtfB8dmVr6tqvDbtz6BRc9S70EP+tFNM16C11WsVEf+HhiiGj0YVez8+GnM
CzhF/ra5m5ItzS7f4f2S83i4bWJRPVHx58Dw8tGQ/n9S20E4mqHiNBX+X852hptL
M47uklVgnxcFAkilg5aY6HQC/N44CIv5p9ABNKpdXqcv1Fgb/LhJ+7Rbltpi0ZBR
zymNrCAwpzjvLcx/FJhxnyt0R5GsxY68vK9TjFbnXVLjFLtc3maSQuMWLRP2mB50
x8Qbb7j49y1hBr+8cS9rbVdbisUaSOmHiRsH4BUAqiZaAGvVTcbJ28MIL/rbid4k
nlUmnAwFyxTW/b0VG7Y0vCNaE4iIpi42L9WUPFWz+dIn4RAjVrxsD3+O1Y89z4js
AN33a+d5LZE37f6j6GP4qMYPnkcyhYiX/WuK+Pd49HV6n2lEWKMSDHgG2dYSPe8w
xXwGaeTd6U22ylErhg1BmUPI26oDQXOgXEhm5zpGlly7Xwe67Pj/v6LDHHl+pXei
XTLCb0HURnKXx1u3F4Qca8CglsLOORItdDaivmhOOiB4yLlhUokMILaYJLvt9UqE
9jNE3w50kQnsqXPVJ23MXDLrHjdiCF5HJlKoAvVsICfn3VKnl6pdQRW1ZxyQA8Zv
lpnJwuBAbjDKlk/lJ/cmGzDA2BB01VdjWT9Zl3Uan+L5k4K/N57IZ0NdU4repoiS
N9nLRu/gcrbsF1m9m2I6Q4nFNTKMr4tAkMlHI78MXn7e6g4URfPuidNJWSMMIfiY
WbT0K9RVQuVX37zMQJX8Oy8XJGWBuxUw2QedCk7J7BxqJcCOheGTP9HU62riS3jN
3LJ8TLekHy8ErUmLkwX43aJb4PxZfk8wzXhuhFFyZD53ZFlx1OcC85d3wB0VcrL7
W1ls4Zacz3nPc+d66iXTXgra3XQYQRhsIuVfL301IMnK4yQthvhp4xR2iso9Bn+o
CnCGW3675QFFtLXSsi+dOlZmRk0QyCgGOiP/26RtZyKo6DUfwl+L92ph9IxY+iDj
GZMk4mdVVbtFCUrlOgOpbc25rjiuBl8Cikk1SZuBbOxqXGlcngkhTclM/Tv6sTVD
ObZzllcqxofViBFS54W8kQAIhPSqPMdO1Sp0W78MRhHRRGM5NQrlEqSDMyriixwe
sVBqlOwrFiIC0SHQj5GuxehX9mLEQmTCMfsJwM+i0/I9Fasmur9dXliprAmRWVZV
EC5ynIo/qn6phGyIGvLuGkNfhuzpEWVXQy7Frp3coMesMuzz1ANwDy4JNnsb+vHw
mzwOVxlhA7013uCbXIqS/X3JGMSd5ec2jsBxFdha1sj6z7lI/Rv7FAWxzV6lqP2v
6hH8XyD0OnZ4QXw89UpgoMxuPIPpPKxgm65ykrdkzg64pfoaZ7hvaAtau91yHLxO
l3hIfBgWGd0o0zgh5m/zLnEA2hbwSNrGYYVNM2subnISFW7oJofOIVHlujaZOkvm
TRGPQbrztPRggPJBf0d+7YTadOGQKe7ZQ7bPY5ktVDUTk4w6z7WaOTh98IFheVwH
DzQ7ZOnMjDdZ6EjXb47gmFLV9QCYTT5xsKx+2RHkhH/mmyLONVhxJulWtdaB0V7i
2FBfnRUIKnS9W6LwOiSF/TWKvjrUIqJjmV+e7tEUyGcEg86PHCCMPjRF3fRQAYmq
lrCAZFU4q8FYdAypQU2CxH1NxpUUZhvSsdy/6cluRrGqzCT8QbEVOkg8vfCkr/Ws
ZTt3kkgAmow6Z81PlyQSwwbNlKpHBz9ebJvbvyGbJe2hx0EsEELsU3Nug6tSvIAm
0wX2syEJijXZWyuqe4ndx4gixeeWVRPJNpsbidTprczK9/xsUDrrMEXCw5rehkN5
X+/c9v9KMbfy35M3PaZa0hkwsP1J99YsnCxibKB2C5iTHEsr2wCzzgGNuilxFfEc
IH7H94zVz6+6EQLS3V0OCcvABAR9BIbC7oZcbzjvayOwTJHRBk4yxiLLsKR+WuwR
t2Fp4TzuMYshFNei7FxRemTjLnb1o7iAKs8OLolNTPd6u2CLJAxouarYopiPqgkW
//wURI4l9DUgKVBNAcoWaAuFQWONstJG89eY99W9AWd3iF74Mi82ucULLb+MeQsE
Tn2Q5E4u8jDTjU1DHO0dMy2wB65HJtVbzkykySYG0c21v/iy0BSu197+N0NiQQq0
/aqrnTLXduGSBfVORLrXsvJAHDu+nJeXP4Cp+V+gGJQI0kbltCbEnX4B37AH0zyk
1vapyqGIvneZyaiPC3FVwkvq21umETEbAqbOE5R5ABWvb+EBTX/5jh4gllH1Ab83
mJMNpUhuq1708S2nrutreHFKY3SUQSzJzf/lR9JgcmzuYP1/S4C41lAOhEcjY+1I
8JDsKelTgHVfv2ZKosXF0hLu8GhYfq6IGzT/4TDK2s5bhAFyhp4O6pvRu6pvHbTn
H5BzwepWnReFkUPWN7moO7q7agZv5AERyss/X3hl/e2/a9Urn1R/LcxS/CoumlCP
zuIseN7NVXn3SgJkNU6vJDcRMJrISm9e1VCzvzP10hqvMg83/kjUx4y18EXvWU57
0Hgw0CEa6TS51SSF86dj8N1ZaBAJkROpmEGLhGRqEhE=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZpQ3GTQnP+FJE4G2B8RuWoEA8s+tQZAXqCwd1i4LgYJU8XqxZYogghgIsvdAevlX
D01hZxlyHmPIzrn05z7FA9Py1WD4YQPcvhxzq52kcfhbG0VEkaQSki8zYPht8qLh
MEXqVQe2chvUTgrDzC6CrQKMVxnNR2zP5NMzEc3Y8Tfj7H7caCXuyVOTINZezGQH
Ob+gB6cc86lhrvxPc8LckG8Rk23iROMUAu373TMi/a0PNr4RTyrmD98fmH3GFRk6
PYQdAjI/hPe12C7BMb6b6k0DgVVsTwjaBLE50Oao84aX1twBBnjkIWVYtPwtVZr0
6N2aJTBscMooE0luwbnwZuFwQlhxy5LCOwhg/awl3FvF2/LpoMk7hcX1lGhYvksz
yp8ToYA6GXsh+qLppAa7A8VCkTaecdthz5XGncO39i3v6+bjJTLZ07FD+lXGe7S0
MNLWMw1q/MEjOiXjkkSDl/7PJv0SJG2ZJoyeZaMOZxnmJ9EiihmgoeQ17ZUSqG+T
VsSNiXslRecXyOpMS7iwBpK8cNo7hYg0LIWUh5ux47zDoxSy64OugVk/QZehy17f
nHphbXkSlrhy8GDiWI1qrEdINc/kH1lRJxW/7A/6xC2gZqjMLmEbyvTYrua29BgY
V1eqQA/y6zBcry5/fGFopYd5ISIxw7NCYq0dj91ANLs9r+Hswx3WGWZWsG9S5BYp
rQ3H7QCjtRXvSlhgJL5Wo25YKm6qttjxh2HgXr7GlEcQvXZ19dvy3bjUU1mlreq4
7+m4RtNJMoE2JHanv0vYmjqtuoyovnJHGR9ZNkddluoY2NGuyDo3kyspH+On9Yoa
SPlmCL871gJ3yM/JiXfRopXZ2A9jIYc/acPnm8MrwolmpEmsRKBiYQqkyL6ZkQHG
VMo+YooDc+1lnFtZFzJXUPAOZXbUb8PjfzRFAKw1scI1TZtvYSqWTy+qqAHpRxBa
cBmItSMZOssVDsyKGfvmMDsjJ5WzzsrurJHAnDbm8GilAAlrO9ie6glKHqd9qm26
TwGA0KRNprklPwdKSWr2Jb7Keh31y6be7OO1qdm9KWveH4weyGXwPotwE2CRpcE4
TWcbmKK1D5jPFYGENyHr/B9q84foAhCcsXEtPHmxEmJOGXmlfzQFGDOlRK9GkeH4
hFFpwKQ0qU7tK19WTLny+i5Yy+x1g/XnaIHKmYmyEMQC8/isdFool3RnyYpPjB9m
S//ciGNpCVN1bqmWnncHjw5fQ++8jdo7vZG/LQfm1Y6KOAWvD0h2/4UVCVAxMOZo
nKNg93dQO/WWC/9H9RbvUSd/bziySnlUyUJfzfdmGRpCIjlDuklJXjV4ON2szp1B
I4+jE8bFrMKnz1ts4KcFeqzzm0n5kJgiyDGqTbCSfiarfd3A+9r71/MP9AAVIN0N
pDaKaqXEfBJu+sGYV5BDRkWzjL/1fenRU8lDYk1+HzXO3cOs18iA4pdVJHf3epgV
cU3WvrDguNOf5UzWIsWZUPrCXe/9zhfbmhMm7OFTGwiDcJd5upaJ1XpCBcD1FlFm
sGainM/fCKRht36K8FjD/sxQVqs8PAJv5kuMvZd724/N4HfaO3e+Kh3gkQYdOOcs
UFHYezoK2KyUnH/LlobMAlXsYJUgjx3lo6eOk1fFKLMfq5hp3DNoet9Ue+M9S+lM
Ij6aR/ZGCkRu2SbzYphWIumj58I16L3ci2MH1FPD81l20gUNCxndq1lIPZjGB/Kx
yeNHZ2pRH2aAPG6ZsAzZiPxthuJGLmGwnzvyh9qgxqS7sv8SriXMPytzDRSqyKtD
KPGRfL1v/CqcQiuNLFttJb6yZF9ZnU+JdEZ1tGkcxSAojuXbYySBM7Ezkq38aMno
QfoKxfEuv1n5xQvAxLYS3nlIABqTBRBMG+0gPxL6vAkL9goRq/KnefDE+xuUZZXS
/R3uRLagB5no9Gl0md2CsYEa9P0CAIWdQZhsPNBRh8JBcF7D0oekvguN/pPva0Fz
gd9BEPOoZNBYGQqFlyNLLHlVFSi3+Z8VyngzHjNkluE73hpSvoYz17M/m2R3dfQx
ss7mIV07lISBvMjx+f8RcmkEfgAtfz5nwr3wAT9VUMf4MtPy16ZxcMWpHEmUYeMM
SruAia4Ud15n8HwX7dA1kq2nObrKsMIwUHX7hIygeqrkMQOX1YAKH7bVEJhptrpa
+vUWfDIPlN1wCTL0suxlPR5ey3KUBkaU3ZscmQT+bhFTMAkYzTww+x8edOX9iPAV
t4sH4x22sjRKNxfKPDOxa5E9pGwA9ZxNdh9KsPdaVJPZ974i3r5lDeVSYgngTe8n
QjLm3aYAalu5VrCbJrQEIcbvhpU1BgV4y2OpTDpRgvB04hr0/+Dbazm3TloqJHMO
ZAK5ezwHQAG0kVYYHScueVOO0cls+aMZfPsEMjZavfQ5tFK0BVm+K2FsYcCRYUTc
PQapoDiL3+QzkNTT/FwJINMeiENqk5MskcgTZpUiNoSIfOlqJSih3Kwn9v5LSRtk
dUlJweOMkVjoQKNkWAmx1HqLruOiyn4pBBsddK9+xtz+nJjaV1Y6iGwhzbeLxzA8
7TCZxaYf2ZS5sTZ3De0Y6uB3yNdH2LD9BCkoKbV16BJ1KzwoLd5IMIzLEV+iRS4w
1sFQfGfdunZ0w3NTUNloC06qbgJ3X/gTA3myA6QvKiW0ZNXwy+IdxT6DBjxln4OL
BCKTUm7swg3TOJYQ8o2hYO177Gm4/+u7CXiBgh3186os3UlASAkO3GgLPXKhbNun
Xnzpr9UVnXz/shUP7gpRrPEvJ1wkVOQbGncQb7Cfjila+B+/Y7Do0dxQAJ4NIqRy
PZJgaFXXSSXJ2sGmyhLi80vSOvi9eUn4K09TQrasEnYLnq0pJm9ACybJr+1LolBC
8DCGkn2nVuCQFg0Ur5A2P6Hng7fEbV+5Y/kTNnIrUMUO4l/4oxk1mPu9SB+AGn3P
yx8zOkmudjRe+PSC5GqheB7GruAnc0gkmqsGUkfrQRfdh/O92JN2Nb550t3zJhLM
uTtQMpAmUWNkS8NOkTurLJpXjp1yGHgpVpvW0iQvwU7fzPfSHM/NdgXYF3ywCLzo
u7MX9idLK40juYlbc3sjpudSRPwKlFnwLucFw5SRpCnB8BuHr5NUs+u+nK3T1IFd
Hq9vfICVtAdkBeZff/mo3CDbCjqm+kwQInv2aDJyIF3imllOru9moEMeBRL829/Q
5M0uNPmuMvH4paacMF9Ql8gFkrV53CV2fOtozhIHG76hRcGCqaRGj58O65j2gU/s
PmYbfQoTXAhCxnbk1Z1YuI0CAKKzwspgBKCprqFddVPNXLd6QdM8CThpXdRp6/mW
p52zSzuq+M3DfkXYMSPAz2WKVC6VpJIxAJkl30o0j91odZkryN3mX3+DYeAqql2z
LYaBNpTtURjmrB8+qfYhbpAmSpnRpDlnokTfLboqmlmWWtDoeEDHbDo2jZdDt3K0
4MscPbC7ZlS/Kf1lSfl0WIuvWr2k2ZsiDS9XLzKQ+hd46lsRdU7U6HHhNIjDgPk1
SY4V0diZOj+ZsAMBHn0iGgB7e2txrWfyMJ1XPc9Fsx+OYGvHFGX5E1Dw3aCsB6NF
tvn9HbtG9YbwTdmDKrMzkig1zgwjRocawVTLujQJGdab7JH3pXFd4xd7iwjzOE4i
AfMgZpOiETRAUtlsC23kyuzQaXzNQ1Mx7LpSbiZZRy8vsXX4Uf+LPS8v9++wDgX2
BroNwD1Rh/pjA23YiFo4xngj9ytUrcEJMhhdWIVBgaPMOF8PZi4e6pDykmgWP9Zu
cIZXZDyMlouFeEE399zTABTlKwpATTF2qdUN3189MZUYlijIAoTuF+Et+AVzyW1g
EpE0oQK6DQPcUXosvpRBsk9VoqvAnO+mKJSqdOf7lw5/NR4lohzIcHkCq6xSsz2R
J+zL73gAdB+pi8tetGFJPwJ3i+WneXw380ClF/r9CryyfoBGEnqFQuyTfBwI6STp
o4jxYre0hwOtJ4bCfPqHI5DJEWn+QezoxR+z6r/OztVIDcbky1hn9M8b90nNVJLn
1AwYuKDUL6V+6y6b6cO8jg9OhzfzFMLKPHSnFifk7teBtHUtoPSNCRjpt5CuEQNP
7ad0mflQuTz7gcH2DsBHnjca7rTcn91G85UjHbrUJ4svYiaDxR26GzdPUCPVOmf4
yYlK6cA3gXZUvgC4X6TaISZvI3qnlS26YE9afkNooJA1W+RdwYVrE6jK1BC71vDj
zUPw8qVU+hRfiO+yzTMaJGCDuVVsVuykO6Q7bFy5suyQRZzKThPI0K6JaX1djDBn
ayWx4s47o8iYtJau4GOmDgdYMgBJJmlJmMWGfndOA4E4eMy/vGTNgptg0s0ufbb6
nVe+L7QzUrvLPA1Z3BhVoTxtExEERGfb7ZH8zTij94OoUHpoU5V5s+6mLFUHS4bz
lGWAMRVeUbLuCtPIxSesYO47+3afDCQtcc3QSXbp566FsG3xf7CMR89dbby9Ee23
YjKjMOhIwUbzXJhmJ3R+gpfAFY1J61WvAYjtmu5oeyD3tTl6R23hbQI7UsEMikjk
2ZshFMNLF8jKS7TrNkzQWLI8k4g+VS3RwlxJWdp1TTZsrmRN7EVFkTU9LYMx9drh
1qiW7+/5K884LS6/VQ5G9I7ZIx8DeEpp5s+BxhE0Su19LCMGTMQfyPPw4/OERQx2
NfJKVjE4r4KInSHXoJLnquh3C7aG4EHZIO1TwCzRWAKav+sXnaZ3/AuRHQAOJDpI
efImNkxTiYsJPDPN328eKGTDumXcNW/fC4OA3dkabl44bG5hiPRhCe8uDexo0Vm1
ss0yQLaFuZPM3EXMV7fXnMlBK4NhzTZ+H+TVSRA3cpSnFXWWpFz4lKqy1h3Yq3r1
Dx4fSwGwTLmV4Qs1atZrX6deRgGLYsZuaD5ls6rVbD6vG2/Uisa7MhirZIzHfeAL
ZVuaiLH5Ls73uEk4KXWpqtfqHw2F6XaqxLbY+W8E1+U=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frrpOGYfWxYHMBHP22DQZ8osZIuSaXa6bE2j1SSa9gqOgvtTBJCUdlHs8jPRLrUG
jpIpGlm1NHX0tZdKamXYqi/1Gl33l0Ha6igm5P31T1rFT7bgcwx/mb5ocicZCgER
8HMRk+nZ70i1vtcbtBqH95vQ3dSu5VcThH1YXBmXNeeyNp8EYzSeH6yiWXmXxdoE
L48NboVjLsaDFmvdmjvrtcABNPXy9tbsbJZ70uqlOM05RsonVSd6kkejr1FlsXSb
c1xun+nc2W//W8vGgzu8y7uTLm6bCgjYrXTtbESQlMoxhoA8vyNoL9jzVn2osfEG
+93lE/D49izJDv2+z+pvyoQhN1NaW0IUGYpX/2Lpthp++6jo7aJPX2fOJfd4xUy3
PjR1MJsSI4BfFZjJj9puZZPyMjT6Js/eRe2b2dXflNE+53LSvvjwXrBhoJY88Rzg
4Z/3MqxcTtIIV5D/+Q7LPMvXyQmedZ2tOfPwfbqkK8eL/uIUP2DtbbDh8oYqnIlC
UZZPCpcJrRcItnJSlVlMqJo06/dBVtSvtEDhw20exg5fKnUgWQt69xwi676QDR9/
RoVQDWy9ulC+2JNnMiuY5oQryUc+3KpNhMvP+PmelmYeE9PKwe5bfzZz9aUfHz4Y
azlMF7UsnKlqvgeF6H+Me9jrbsknjX59lbTz3pbrxGykAojI7vSjzUy9ncNNxdsv
CYTP0iNa1Mmp0tW6XymaCqaRVmk11YA65cSm4gyczMPfmWGrNMx+ROJ9iUTR4K6T
N49P2i+m3FQo+7EToFjwGHYdcjDyZ2YSn85u5AXid2JWYigpQ0BS/8tTHvQeJ+Bd
C5Nbfrp0MDD4H8sWvUThAJWYo8WPPKmlQSirCCcJBi+HTmvYBIw89GW1cF3MnJvy
X94nzLOeJMj2IPB2KYnZyi5LpyvfqTnhD86Zkws2PJWNskULViF7P84opGGBdqQG
aXgG469Ct+rfoqK+qnKt3DECv8jnBeMD3LGk43qQDB1TB2X2zcX5n06ocmgtR0To
3hmoBG81fvkznRIIhrKmahLHXRkVzmU/VOmhk45Fag7rmYhhb5e/86Cotfhla8Cq
9nSOcsq+y6CT4dyYL2hsZM6DuQIlI9ScE4Awx8Tr5S1f/uF9L2IckjXsXy+CYWdx
Ww5jxiYwHp9LrSXMuIbRMPhtqiW7/CMSlHNzBpMnMHd15vNdAbowUO/LmJt0CWyT
lehwM9AKORn+CPpsmnjGqVPSxvaHs0LHp+B9xyTChjSNP3UKrFx9pRo/Vzs2T1dN
awneHf11fcmDAZB+wEu3+KIRnMPIc4kZ3X6fOz9pQdD9UErg/tp3Y44sw5MoUw19
pwQWmOJ8QhWq+du+MdegHRTVd8ZWDKpA0NV4x3epd9hfn1brxJRRUex+wDHcBysY
iuEQJ8hCJySZJTWUlvSRTfIoKqsbNxiwvJf/a4dpv2TNysJHmOUwvmPgUAnzuo5P
su3LNLfMI+4a0RTKdfKJe45LRyLgA/ZBUn79g0iKnEaSSPljpKuouP50a29FhSEo
Xm/oeu4nrjfd4nYiA+QyuiNmZHucHAmlDFJK+25OHEHoAhtNGove0TaToBnH8+KW
TB0/fzh6NeYiCIpStLpAhIDrH6r7TjOK+NMQ8yz45f8rR1DPzGxTcsb6KNiLJfqr
meVFl54UZVXpweg7MxxtaQedMLIIcfPc3K4Ef1daczN0lMOaQGbQsBDZy42JHUsY
MoJAtvTCh7DTUOPaiIvBTAm7NNs7xfn+I+TK1xicnsZHnerQ1H4REXT6t8IBAVQv
0lGOcEQ2HmC6DSH/SVlrK8Q33+vRzcFVseHzJFBtGtYlijMuuq4joc8ko0t6xaHK
G6YLf/+/8RBP+PafGEcKPA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwOdonibG+cehHkgUDHKDc5dHkJspfirphxSe0WQ5Ax4j75lm+9cVgcG6cxQ1Wvb
j9LBpRpSl+Zs1mSs62Ub3WIPpErPE24SENWJP1zkYQn07KD9Q8cRKECMadZn9C3G
ldzqXY0/aFmk8P8jcedSdpj9O33XX4Kpbt9r1lYJzstF96O/9foTzELDncWeicG0
V5hET7Y5GmaVobg5G5OqVEj0BkhnIkdSks5gJJuJH9tQlQrepiMPe16XznamuFdr
ms1RBrXNHGyvldS2LtpxItMpTlLr/UaTkqU9Hux/0Xmb1HG+3T8DoM1j+PrvKr0S
owrBLg30zQx37A9HuVf4OGQOjC0dI2CmJo1UZf5He9syTE0jtFmI0vUW0C9ExleO
AmSLuqwovLyEBf+GIF6oQbd1XyBrzFEB2FQC97JDfHQmCJzn+fRdhG4xJRNbhNo1
f9X2fnMoAQmgCdCRlWT3JwGibH+TR2d8Eo7LKEVGiCziM/fJciACoaGZ+xMzk9GF
DSgNivaQ6MWKJYaXt12DhQx/K39f8NcrTQBs0lvE1rCBZJL11YcIfe9XnlKFEjy0
eVhxwcBuOsamRw1IwHujxUfegXzNxFHcFHZg2lPs+r3QNZHcPl8NUwHkVdu4TiQ/
g6Arh+EknZI8q5iJ4BQq8xLS2kGoowFDjdHaiDHgkh/7zH9KMiuCxlb19NxRFmJI
fO0y28vfDdk6R6Uo9w1Hw6qBuacz7AQl0s/pCJPCPsl3OUrjBxrn/eAW3NwOsdw6
m+yitXP3zl0Z5Zw2lidQMamD6x7d8uOrROQBY6ZSbgZIA6dejne4WldKHo0QmWAi
WoTO98v+n9tVI2FzcRhtwFKDmpmXVXfeWYR+/I6kwL6HEkYzhRCsvVn6j980dzGS
50dV1z6y8XQxyeJmBPGk8f8NuHe6Xb4nGGD4bwYhK6UUESDGz4VH4WcqdxSxGLqF
0f8x4enIEaWNvqC2m4s5LY9Q/6KkW/pzFhJd7iHZ6G3JW9FCNrR4Cz4YE7TFDysi
ziQEKR4QLvsvM26ODL1ieTfFKr+zOK4RfGd3bK9/XmB+DZohiT9nzNOBo7Yc4bGe
SO8adbjIZfkIbeRixvImxXzdudgfZMhI9QBVLL5Q25GEpUNxkpvcLqdrU08TDkxF
TJldYt5rJkErvdkFxvI62DpccLmxqSXQCpYLCiy23imN26PBUjT3HYTD3SDYasw7
LCQ2zegVh/lvNBfba4yPtPdsEqmN/+afrdGXMvtRob/W4evpV1goeLSfsSPvexO2
OuQzrLyEx3OEas8TxhlBBbAi+YlEi+p9Gvlq6ktbt7L8CZZqNyUIR7o3WMRHs3Wa
tr7HLAvekcg0xPg5WC5/wGrEN72aNr5wv9lZGTg+mnYHRIf1Ve4kwkKMWnIH/eQd
QfeFfeWtl3AqB3itL+ttV+9H66XbM48IQXxgLqKbI/tk+fsvJfBu+WJnkeufvH3N
rM+/CA/pp9rzdzkJGLOpXqQWztEbqSXl6bDexyB7NbKmyXiyQectEaq1lsbb3cII
YKoa5JC5EtPD1zdn+OhplOZLpLBKTCTI87SK6KmMULWi0Pu/BPtbKPGZdXkNI9NZ
/uYfnXwAHxkSeZx2QG55Dca84cONmjBfT44jhGzVqkPUP66SGbbYAQ8WbCpSNmE4
YWQ6sRMy33kC9lXnJJMFFjnXn77zeN2ixL8fvawwmys5b/9uuPWfISyXA36huWPw
X4YQAT/TfYEGOQ4smLnSltjru4reK9qoEV3cARvGtj336CsFCQ0M7GOL1oy/SiwY
gaa/qYRUezCPMTwUWjhFe1bysmSCVXWh3ymVgsVJLeo1H634mAbYzwuKA7aaFv2J
KquEi4pJobrXFZYe+R+jE9BmnOrdTgXkHNcn6yX/4f2mjNqGw5oHnvNirtzUEP9V
AbNnQKMy3icZKMF6UICvz0/wSTJW/ElSrRECzUpKCalGY8O+q46Lcv34XCUqNwgT
MCFtmNm1Gczay9QxE05ke+duVpXeOyZirfOqyyphY9KJDCNwoHnfUdLTN47KF4jm
FFWBso61RtkW7rK9EZr+cFJIWqHjkeGihnZoCcXk1BokmZ1BqP3C933/fs8zECFm
DeuESg//o3mBQqBw1ar6/f8XmoxDDY+r18P9p9pvLyXLmH4PLmhWG7XtDKeIM6l+
rADuxLgt5sw2BYiRLhcbh7GsOo4rIXklwR4sWpo/zvRCyUIuuaOHdFMRIuPKNqET
T/m4QmObIe0gR6A5YfEXJm4l+rjT7d2eh/dfx2SwasZKN2jlIvRUurifTsUIFYEA
LOQb32ROYLWjlJXEGcKz96Ty5n9xoSX7qnL0oIR64dEDAt/IAuIlUKwKdkAIebDe
UthxSHW+5AU4HjEZ8suuXTrx1D4yJ/IGZ8v47RkVXtPbRXxs11DYKmRDG6b1NTqs
sUdSPGBXBqxSgbGH+YArjATw8YTRQiRP7aK5EU6q1E2eWU4I97Dk0NrsUCKRdUR7
ND55JAlgWU1J/HEjzB/530E9vlHzy0XfyUAwf+Ur9O6mijIpsodJ6dWnVNSupt35
epsvFAZ6MSDK1OLonH4OohGxqPRm0r1ipZkS8nD7CFug3V9dMK8djOS/SW+NDOZt
B33yFV1zJWk3TZA5/bIkGoSiRG8m+WAkYeW+ilfvibsxyKkYQXwE7COFypGHlO8j
bwIJQ/oqegZ9ycU15nTrg5uBaau6RPjh0XN45VSJ2bOcBENfV3B/hVAxTJHZIB5K
PACThXQ727KwbpiscdQRMrs1jHQ0N8AV7cBgJDVg71QyxpH0QDsfJH1b/PdJkVu3
j1V9rpKNsO3UXKUvJFZkAfES8jPMF8CxYLSkezicGvX++MTPzo3YuWzuXhTyE0aW
P9z31zFQOLxcISGVT6KW9K6WkyWNFaL8R6Jigplu0QS9jL9kaCXIehbRcWJzWMuI
RO0XjuX7VbnNa5DZffmZzW9FI8wpxJqXVh776IQ5WNl3pCYo7cICQFVXWV6bPtXQ
ShldNDdU5wY7WCG+IaVW6Z0KJJk8Zhgbe5XG095WGDEw1BvN9NgnbagSHz4KR9Th
36fMSe9Q4KyZPNdF96UMWSpuExFX/CPUyLjS3ERwKKE02PJuKHqy5cu3do/+r5MP
vtQtKZTnkNa6poZpvf/bPOgmDyu5HpHp1vdHPLNuH5TJvwbbbwaGTQ62mZ9/Kyrm
XcZJ15E+8AGTINtXgpl4ILgKiBjB6rkE/xgSI8V1dZE7Z/m/ozUgNfrYO7ovljsI
IjZOWNR2cbVqwCbls8Rmlheflp+urD/iJraI2L6FjHDEZM/lbOwJAZb1j+tUswbD
1ELVfOD1x7leVH4UNyY8Uo5gIfUHofHVg8mxZ4ZFM0Md+Ymrkz1K2IRCbMKB+jy6
CzRWKNcBVc8XuqaXZN5AxeEvtJJuN5xTbb5bPN4Edy9RlZ8x5//S+UD7CIwoAHbP
EYJabJRzZNtBqHCseuhBBaEowGfyjmUHqFjtnMfYzXPxAocPsXzHVtLNjBwccd+T
kUMiVBrJe4nf7ZnvJBLy4dxr8n7KT1p02mztQ587HtNzX1lYgm+yl0FIfP8D7onh
pbG7yM86eWDhxT0js0/trWMH+dcGvSqRD1FbvLsu8rGwlz61dDKdEi0DlDrFaamd
kecbKStLejmMiW0VoWNySjP7DTyHiOQ7QhMh18j8qJWw3tO4IAnZV+baZ3SkNIwX
kA70eoAr/5Q/0uCaGTVA0rfZ71GdgyX0/xnY03XvZVwF6ql+x6imXGcmpHG5wn1w
YLTFKUZhN57v2dJV/G7jnDuVtzQyE9laF+LwfmgHODewlKhPryuRJtEE0Xkdr/QC
U7HiPb2AKekNZm8aptf3K4atPxUH23xeG+YDLqx1xaPXV/FmBmqrd+ubtu5qoxgX
mllo3DWpixcfLiR5iBmMHQzlYTBcqZ4XIAVhTXu7C68c5qXrYhloCGkmI/mCyCz4
tHPIrSR85Am+0ezQAZmGE8phTPF29+vUZV0q78FWI5pU29EDKmfY9OW42JgQnv+Y
fVJfABrvd327QLpqoEldqETYr4Wx5VeN8E4d6QAaDRYJSf8Yip/QmB1wblPVyI7b
9UjE04DGG+o9XpCYIICOaCHMrEP5WW4xXCzxbAJbaG7N7blGPUnTPEK8s2Z6MBnC
8IwZAG/7OtnCvm+n+okhR4q/lTN/iKunJsWPjoz6mR2WV0IA+dTSYnGJlPK/O+04
IFk2GsLyH9uc22dICbGl1ZvhagGOycfxElhIGRQXuNBUnYPcokZ+A3fyTsH/rj0h
Z6DsUW5hkBXWm2hRmUrXxE9THe9pnnyU5QB7xy/bmhl3S2K1sPSJXUjLqoMW0UQM
sWIjqcKoA32HhkapcgcEcKtNsIAHkE4JqQGmXyHQOrOxmJ5rIJR9o1168oXX9Tse
17a2RsobH0LenHseWZBmWjrsY0iVuN+8/Id0Ek4DfO0oCSq2TQy0wA6U3pgfYYoZ
BmU9DkuguNAGxS7JVsfYoLYECmgGnxnGJ5MZOIOGIM7UANpY1EXRunitRP1IY1Tl
KMvh4N0sUP/qBY9LFJlGnv6PAE+x7IB3eJcr+dMjsiL/NGpjz4Xcf6pSSarcEbY9
cRzbsV9sWtnHz/20R7cA/reQaYHiqayLJz3VLPy66D8JQ9xOZwI//LYYsLACmm0/
4t3rkc4DFyS66umFsopKz4g/NBDxqTNorcL0Pyyu/uvWqwybA9oN5vdGA7Cv27AK
winh0ZfsHSGDI5GCPLM56Kexpjz0xcxqK4cbUsyqVEEacP+qKsqru9ELxyVtjjzI
mgCZUI/6eKtRizqF3PF/xMicXi7TR2lCG9AaPZZYTKN85Y0Vty07D3Bi5YtpXiDh
TPhEuFbvb9yfWr24Kd17LZQar1sqe7EBo8lff1twYx2d5sLLUJEioU1vuO0JfkN4
B7vyfrRofV261oc5dn4u/Kirude6oKXHo3FNXUB/Yt52cKfsYy4JC2tBLP+25w2S
YIUyhlTwIgP3/zt2xTk7mvOi0hGGcQspEW5JL0qreADo2t/8i9xuv3I8p8opivx4
C67PcdZSH6hZvXD/BN1wW1Pxm5mlk2bXEIYoScrhW/3FXoTX81ySnUxHVqs8IIHH
XSAEaqnA74z4tsied3/5vFJC5ULnwHf+xYbVygPXO6FP1z9yXsMdXGSlwnzhpVIu
4Elle59ZXqLRdDQeQh/GstMiU8G6qge14aNsk5O9wQUOuGONe228X8AScai+Eiwp
A5L5PimffiQRGShVMGJ2l+aToELIFajJ4vrPkT0rkxdAVKbJ4K4nzoronAlXt/eB
P84Bpto3zDZEy+LsirIZ9nv+FHvAnu6rgqR0WMxvTyc83VL2a107VjUoBDbgLp82
pmtdgYX0ezzbh4qcimiTGFZCtABmy2c8a5a36+1tKHyvfhJ6MGBn45owpXtLHQvv
VJdEri2HYbIPeBNNJZq536Nm+VR3sqpRbezN6+OKSLCipqLzlGAN1x148La/fIRh
yjdST/jGfYVrzCTbvdAgGXe4UnEDZmORyQfe4zFiTQ16zjkGQjb3/hRyWwGIqyyY
RHRMlLDq5oIkkVI4Bm1RKc0YbmtkBUo2RemlKR/htmukYgEQlb+Tm3LuhkQfF5Au
bgasFeKddcs+SGyXRb/IXEI310yqeeDZUgQlNdrSO0EE72dCJyYKwIAwdXGtEKDY
nx3Yl6jP1eEv3GNsc1E+Ss7jW0EnPegQ6hBD62YHfV567RWU+Bt505czutfUSJw6
Fo4YbTqnc6n647qbcb6xQqpYdZ73bC3bcVmJoVSHCZ1/f/iHxmSK9ixtQMWFBwY2
GX5Tx34Tkrs+WguSDVjFTCBsNL2ce6bMWPNVSagfXeuXmKS3Zq9CjDVBq5p8jDF+
IFReHXzNLYnMkWLwO+lMbeOfgemb2w/BrnxRRSA2mjlyb4ntvvXsjh4HbyEp3jti
6ZDeXuoRu+gwCKe2XukmBCNKvDGb3xnexvxxMzRcmc6g60VKrv1SSDm3X8Xro0M5
RDzdcXGEl5w3SM9sqhAgotQmT0X6c5SaYXYTu2aFsUS75YqlzwG/1GSuWB6Xqizv
z2t8f2hdvy7yP/YHXkGX/6pHbXMW4kFjcSuKBBJcFoDKYy5LXAbUif/WfSxzTKfU
mn1wOOJJNJg1JuxeU2tGePln0ZYubVpzH3MyYkApQJgf/RlS3ZP8oUv8+cZm+RRR
bJyaSAG9YCdDspk3e+kfW/tuXKksFg0ZBVHz5twErsNPKPm5iw/oftHDveJAAlAS
MigR5GmnkxWVvJNe0znloUIL/KVqFKYEA7UjASIyvcy2ZtLiAzvtoKisILlPiWpa
qeoMju5LvpP3cLkZz64vfrUsOrEkz/gfoRa5QxT6SFG4CTyy+Noe5YbR+4/ejMRx
i6CVh+yxdhEFh+tGp19NP2Md5G7pNCPxo0Bhets6g74/S45MD3GGEs2etrpeetQV
BkTmQNC9zoRhqOWsoMfuo1dRhYR4CP63gmx6bl2BKe/h5hxm8RdtOqLvPOC816Bj
WZ9eJMeoEKu6MHk6K1orxx77T0kKu0QDuM47jcPKQuyrR67hvhBZoJbv3KsJm21m
5XRmz3xzaz1wTHouN3W4YVxYy7iEihsyCWjTuBlPslrPVg66c2r/bW/tRxEfwm1i
WPP0/yfCIwsohxAS5C4kmUpT7HU0o/QAKRFYe9l2wTsocCS0YU9puT0Fd5jZEFAU
tJydhOGdw1swwyCtLh1KxNBI5lg06Ykokj09f4c6ero=
`protect END_PROTECTED

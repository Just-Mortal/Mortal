`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJeR5CMoyWWrpCZIvc9blfwALPxHXoGT6Mp3NfyQb7kp8bFiHjzYoywHPWpGzteE
HEy9WeUE+fKljlVfhbOl3EzDxWKdzXcYopienl/9WH7M/IxTUMaM/lzzWhkKXUUS
kDr9JGqm9GytUNo8UZmzhRU6yPtPIo3e6tYD5FeMBQdW1iQeuntyYsMZFwnMSLJI
m7rYXMPx8nR5mTcBpnUkniP5rHrf8gzNF3Bd0Z/HiWcrYlCj826MGGjkqHVgEXiR
fW9jriGxQ4BTT6JEdVkuaASDxU0fuqduBlHVXTrVPThb8R3I5ha6Is2KhS/TWyVL
ucG7oF4wKWpbSw0bjn1zNR18OwZfH9mAEHWub9llMyFImzs56kcBZymzBr4YjQJ4
YM+U1fUT1FBGakbiUPZ9kgaLPoLIsuwT9gyPEYo3+154bMEYrsWSVwW7l2VOj1bu
iTbz1KNs8HRR13t5o0uJBAkaTpW8rZF7NgQL4wq0XzLzua+KczevOueJskNPTB/W
Ab+burGD028WcEZUoW2ZDg8N3xlRIOsaJOuKONxxq+zzfetwsl42sXcAc/ksJ5Eo
H5x3rQMotxnRh8R4Z2fQoSN68HpOV5tiCoA3jeqF1b3M4RWdI8Njw5XoxbPxOzei
5TbEry9qFcupqa7HLWPj8XSt1jyFOHiC09oOJBje7UHZcpamxolYeXypXa658A33
JtsrGJx/dCjiNbCzx1QJk9YEi8mlE5KldugF2uEswvh3M+q5LC0Y/8pIqYzaAEBm
t9vDW8/NFYhB5gqMykoXZwmfIeNMm21U2Jq+AmIVoy3aYdI6XD77jyWrfsyE8dqY
XH3oIZDM6Y8upvp+DXiWmLaScJ57UHc9qFnMTGDLfyj4W0LkhI141pJepZS3e/hc
XmCbkOvBvxTWr3iYkEwZ64q4pwZ0yahO5KjQfub1P+xTaGyw+6iOZqqZK1l1MV78
O507J+XqXlsVgnFIFpINSntnz9LXvpPCuEWhOfM0t6VvMxOEHNMFpZoyRHmPeMgG
ZlUfzeaL+aiCNWd7/bPqVg6wYfV2HPWBPTwI7gNBMG5iP5IhH8peZFujqUp+3/SW
G3bcu7ioi31fjSo/ciGkeHYJOnCfouOB+KHUEpJBlsnyFqRML+QeMwErWuGAY1lJ
eunZYvFX1++NhDOEuRxbI+t/Rn5X1myvJ+A8CHJGIxeOeeCwGXcTdsA6BAgFxPWP
Qu7RE1MNL99CCBqtUjn+hQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fcLLMPV2HuFRDNP8ABJY6PVbVPb9EN6IbMQ1W1m22AQsE2HATnBUKXbq1rlnuk7B
p9D33Oqe3lX9p/YN7BKH+toAyTxiT1SSt3nF+bKSjWh8FzmS4YWGVillugmu5U6Y
zDIQ4pd+IyBF8c6mo7opOzHtSMmBvJQ4PZDVtCn+6pnrDkC7kRAMeqVC1k6b93KC
Rz36ZCPc4Vf6x9WUTeqkRiPxcbNQKFw3TE9XZosMrm0JXein9jc89RD57z5gs5Pa
GVKkusY7qPygYUhaBHmt4YJRgSba6XE6nc4AsDFtHZhPQg5SiU3Y54S5++3RPAty
8uqJi+DPYryDGgbev37gLm6HgmOliXuDmCznqfM5OTiSgkVAEbg3ihFeAbHPhkTV
jZRxsTPRqgV0T108FMuHChxupRxFBk05J5W7EbqmZPb+1uhwHma2Cv2K0zbl01Uo
fm/s9IYhJbGkkPHy37Q/pTwN1K2ot+phLK+NmyfjH/apcsrJhC/eps0C8qHbD66p
hLjOgRVrOZRBU8uYIt+TdiZnrACHap3tt/+v3wfe+N8xwbXCUlggTIl+ULneJIsv
zJgiY8fRey3RnlcPDfHK8w/eUF9OU3mAv56Mx4N+dxIvkqUvH8UBI8FLb6q5Iiem
AqFbVXgcXu2miBBThdcNaHKzt3O5iKnIyDKW7S9RZDkksXJwDKp1OKYW6nmpt9Sl
VnU4HHyJfLV52XpjRWXHWb77ImxswRTGr8xqo11pqnbBfB1qwKq/FleeIyUtoSwf
1Jv2FM4ebz7fEBh4fThCKDtFizScP0fmTxc4lqOM2jMyuizEdAmV1UdmsiukOLnA
Abevl8sgjUnYX8vD1/GJyHoo6f8Zgj3Cu9zPqmKSrG8aeR7aNgoFjGzWatPnm+2k
P9KpUcJZyYOnkjOIosUSOPrqZfDCo9LrEGQqzSrqYUhPbL2JWaX2aaf/4f4Lea5+
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRlwm2HR9UT9gvcKDstjSLkwzQMsAVwBAh45GgZNlBtLhexGsApn8O4TXjumPALb
xDcXgXkFsMuZt/2JqL2KQpebGTazHak8151hzyoXlfIsgydsBmwBmFBSRhpiJXh1
VqSumdy5u+4nD5kr+5Z/w2G7LZxriSyVkJdEAebO+q+nxAoBUKkNaO9wegiS1oEC
i4d47ctfqUeAWA4E+pu1y2v9cR1gbA/pQ1kynH2MRhCIoMUjDfrGPoZp0Xgsl++J
sC7JDI1DATgI4PN7ddVdYlr1ubfCPWkB3P2nHwlTtr5meN9Ec1T9fgiR1JH6HPHm
Ne2zkNB5faXErQb87bEfqUJSQ/ba7x/BHvo3K5lvp9RbvIKzpuEFpptom+kQQCxX
c4sz1DFqzxODBQ+7hufednaDE5XRWajq4N3ctmyTE9sOXAL8FcPhaSyZSPl5ENC1
m8753iw+U3XpTBKRzFbZrZKXbQ9sKCADTvt0NLr5S8b2EgKQ93CHqGJathpu00Hv
fKu8Nmd6gsWxdfSQisjXy8RLFsaMtu7Ke/mq2iAaRIt4SxvjrQvU9EPgCNWs4Yhv
aTs0A5AdozNEmHDqe87t5mS1jwN2YAz8CBP03siyGXMiHAB041mendth4PAUtLLJ
SHCNTPYb9UUKBGQxuxMezTiw56dDZlL47WSqJ09jGeQT7agWEWKN2bGXX4vxqab1
9Ld95sMr+ceJBKarssn9DyZa466GlzvaFuLMsCmFqGnP6t6YyWGc+ZGxGdQN5RR7
pxhYphn73Cna8vAkCbCnXadzcYGgM6yv/Br4IkcLyI+IJPgReDfoMDAP6DuCM7Lg
qvcsZa3lR9rZoD8PW4kpuhbU451HZIX6uMA79nd2pEqlTV3icWD2bYMquPGbwzn5
y6b1uOOi3kJQjrCdOzhz8d+gGpBQX/HqM+5s3swJ/6yeJGmpHaoDqme5vDoMrqGl
+a5PP8fb+zXSjO0drzoHrv8rjw3h8amjIMhrPdiNbvyeuZgztBod2Rnfv6gMKU27
a8YIkAQ1/gx1kmzkJZQ+KlVTC+TPXGTB6ORabZ3iZIlAkIZoPJWjwiX1kIWRVS4Z
cOx70LOz3G+3AYlqxHaa7BEQeVIG1P26gKhXQg3Mo8AlaHBww0ax9C0+WnGwEkUK
o90KfHgf1HZnlLUDFcmhkwspPS4b9dSijhAVNYynKnyqE8FiTL/mxStBe1kpRise
PHx9/CimFpFkemFlV9VjjSk7d872f2ObDMR8lrNbbQM=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CECXACjm+3UQXLtke7kQyU4AiGTOxUHGplHdETd1vJFvTq3rrYnMl2gD+pamiSWn
f8Up8QDxdY3RWWgENYeKugM1MO4FynpLvOhreRFq3ZoTxrvi5Qj6fY7HmeXmyEzj
eQEFk7vGihnA+Oyp5WaWtU65Wexn9tvd75t39vnjlf/QyCh90NWdvFhQ6hbvneb4
KjcF/qfsU84jn730C3V6k5QRHPfh1sSq7wrDN+Im5js5vAxDia0a16ZFNtFzoM5S
lw4Jba3Si3M5JfCqurWmuQCkcix76m9t8NW/tZdB13hiBK6D9BHM1T6FJN8KQbJy
PgtbhZ3vZFgonHYLdTyVvtFJ5J5LM5TNDttjPaK08X+eRSiEfKFuYAFWGSiVl6NM
YuES2mePszca0YxqwRjR/vUV41hYR9xD1UVm2rBGtBdCTa46bpwIsyq7qYWe1KMV
zXqJYE+dSPw+Tpbupc/gU+uJIQzkiGuS4R4ooZFy6iHLusTZ1UHNPrLiOAaHn3ao
lfpvcFWnhdD6AeVtaOsmIceezTSZ39Ql/8PpfQUdWcD5R9dBwEX0AFYz4nDNaYVY
ii4t92J2pICY4Vs8pALeB9yDDApZB+q011RLaQoXaXFhVYujFnAKAyljDIDo561A
1drN5kWXuWdAVfTr0s3VaWSiXgJpkZv4yUI/hcu/m694yLuxbghneBrZQ8HcNVYj
dUvQeAnW58hMOYbb1CHLUbxnccbgGui3muwJBIfuXKu5dVBLtpiUFmubSGCj07qf
PR7kvEPujENskxXohhkh8bNGgUloj2vp5OXpF7h8845hZhkL+c4BeGB5HJN6rNas
dx5zQvojlS6MNBfw0wEM6fKnWShR2aoicI0BOmv+2eCgC+dNovT5XStt+wLgrE5X
cpirnAKdA4SkvEwy6aOoCbFWSAXeJVoB4d+2KBgK9QFX4SBBFseu+ihjt9i1BxWs
hY+0nRQ1f/uZkCyftc6X8yAZlPBjQFUcYF/JvMjAhZ7Ro1gBRgHSeks/kSZHMERx
iSeIWDdvjdHhQc40xvE4cRdSabNhvmLGPnvpLtc+2i/Ta7SvqH4RE1dttziZunXW
NbgJdK5kCglgr9GjOZ7ZalGRGkljSqTk8MECMOx0PQtM9x99UGcwcfcDEpu+mY/D
ffYi1//jv6YJR6xwPm8u+0e9T+B0FfgOa+EC3ftRGQp4bVftGg+ZEy67jzhf8VnQ
+WlkIoXsum8WfM3TO7qg0Tx/UQihA/dJ8pU48cFgIpGHHi9StdFVK1LJmGqvhOz8
vf1R/7PAME0VJlabT7PnF1XQqBxP5xYdY/8jxcZuuItdGI/n9TTNQxc3lN0q/9sY
0FGitW53JvUyq97jQbVrnJmS4is0u0UyvoFIYJ1R2AbRBzjID91xPe9j1TRTNhnG
li0AXzmaGTEHJRSRKUVXX00YwJQWOEQtBInjKzaAAQR1pYegrY3wmwPHK/6Q4kRV
HCusU+XfWIwJgeJqtCJvdrt6hEYgJWeOgpJf2IPemMaC9Ptvc5w0GVGRE8jP3MOK
AswKEMrty+O9K3QStoKZRLxhlLtIesa4otSEU0gjHHBTEhjSTmVzi9buQTlXKcKZ
A8iDAsy36R7UOzaORE3RyzxtaEL6RxkWqZ+H1zyGoFop9n6oPVszTwuo6XpQHVyf
g7hAavfXpOZZVUgyZ91IrbIBRaSkj5JdtW0OpwsrjqH3f3NrdJDS7X7BpBU1xCYa
TYV3iX1Z4KpCAu9MwXWWUtejZSau2pgiVtlOMRuIbsN9YlHjUX76s2HUFJN6oP2I
SXtX9ULwly7bMb50mzvwVG8sleU9xNQ3lby8BsQhG4EDwQAi+4L0bi3IJ2u1AuJt
RX/gd1ohWsixv/M/1r7QQU9nGUJweCcV4KUVEAY/PL49JDBjoS0M2oYtBA15ndo/
hc23bxpXuTIxm1YDEy9rrKmrCdUk/7MuBJA6jquUpi3MDpnY+UMIhdG+NU/FNRz/
CYnR+ehAQ73aPt/wXhzzGrVkJP017Y+tXRRIx8XxbOj8oiZ5FSdeBkA9H4e2n2aX
4bvy5ezEk2slGDHGI+cLhS2DcYrn6bpOSUIvhPS57kw/L9Q56ZvhFfjdqkgTy0s2
/ASZnCIH8+utW4BB4HeHtIPYXUCdKjW6t06UYKlktbpVEn/geR3R++giGngO83t1
QfULN93wcXKYE9i6vh5duwMMRjlPjtIXdu46+TWUK/2oEj/o1xKt4LMD2AUnBtBN
FnU1JoN6KlCS8hHElPP2lxZJ8BlRA9yPgdTMaD7tjGcLBsfgwzT49plyvfr5n8QL
imOtBM5oDK+JX4oIFmQ8fcNiklz4H4GzgUatVWnnavzrOa/9qryKMcIuFqBHOFvt
mIvnkZlWNRmjCeMQ98BDXoG2r/A3dJWDD//oyAHzYFqcnJbXxxOFKqBJfEXRX5+I
gkburnlKY82LUUXIqc3gKnzYe0OrEutx5Cd6fgQAEd2dVRLm/OxHnZPkoIAQpKVu
bYArh2WsxNUxTkDjo2o5tku0T29m/yJX3azk991IONCXM/174L44cMsctN1ofjTE
TTvHbaTRgWvCwpDTZ4LUzFRqQ0MnBzJq3nPjqvWKYZQm8KesU0y4dmy9R4tmkYAe
vPSOA06jGfj0R4UEghK4jzdiNasRUM87inv6bKMBeMqYtXdT9Uw1AQt1k3i+V3KR
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Be0n4X1Yf/fTxTlaaAbVO5WHyzmtf+PHAaD86tRmPQoaZ7vXZHDHC4rWkWd0qVB
vMjE0FcJkokqj9Ez6EzS4zMgqSSdI+W8kUxQWxpRkkaDMm/YaXTDjBaLE+8qBNH8
Tb6DR7bJ07Ks7kXXKARaor3Y9xbBPEqYTrftVj1eGbmC4yP/htJCnFLrkDd8SHUE
YhXRY24auzyxGmtWorkU2hL/Mq/7UqqR2u/pCk9KnVRmNjFbQc78L6BxFM40Txeh
9JpJwk1EzZMD+z/peBjmcwiM318iD+txdtcsXnCt7VF8A2/Gzxqhho8Ny+z04q9l
uDw15cW1SSbBdE9FBK6d+UzE+MxMLxpJHZZlNEcaS6CYPLjky7RZmxTILbvJwRgv
kCwBWsPkNVkHWxsoX6kQDYBJAIo1a8QB5T8WD1+nKW+1Gkg1CUqHXTR4QuwlKLf/
2AVVNR6Py5/SJ3IqerArSR+B9a/gfR9PiYi8tqSvdLmLuSWZW+RfaTL+xlnYDFxV
RJRGLzWK0IBlcmXUNwcZ/eNmRTCeX2HqdvaQxZDQqBxdWE7IiT9hRRDFwHPfXMXh
V7cxcKpe/DO01pmEOcFgOQ==
`protect END_PROTECTED

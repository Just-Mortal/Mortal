`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+eo58CXq78jlnnjnsWerqW560aFofUgnrmActI/ET8jJiRqsImm1nOYU4ofIQeK
Q2wuVRucECeKygXR9iNsoQLVm84a2+aky7Vl4RKln/iz8DwY76crRdtZiV9LrNz3
UPGEXYqtYziS/7I0SmhbpJ/qDq1/Gdvqhucn64wypRRNOb7WmI1hJGSWkC3lqLPa
FRc2LgHbsb5auz+no1rnVU9JgsNn54pYVgeAufp42Di4QEwQaUpLv8sRK4ECr8Va
m5ffRBcrdSshxCzSbLTNHxggWFrk4apZqHZ5FMIHBKZLi9C2bDVL5E1RwVNV251T
ePYVjpEiBTs0wjCeDRrRJvhAs4i+2MsRQGmrz5Nbv2NT3aLLcdfZZFVpMu1j7XCr
i2gisPFXPIYj9KzlEMaOiA==
`protect END_PROTECTED

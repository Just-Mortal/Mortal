`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrrwNk3WzSKnEWoUt6HmmSREZWQfLLZ9ms88afde4vvLmmaSd6W1hOyhYNDF90NO
spezU094Ljbq3Ex8yC0+3YDBNaq5SAzlVqUuZZS9hjjwjAzzFcUAilK22ymagX66
kaJ4AXR86/kUNkwy6+L8A7kWKnr0sY0xyXWi4yGcOE/tUVIMmdCOdwZruNuLJjCe
KnLpad8QVQCh6yeMVEPeKcFI+fSn1oDsvmhgx9jn3Ug/YuuUzpsl2NSe7i8r1TiS
udEJ9znhHw02CY+jV0eYkNNGxMLtPjCbAjt6EXHLhlMoViskZb7VhoYGvKW4Tk5T
EoS2owLtoBkyfY4MLs5V0vTvot9IGoWUx6WOKRbFYe5i3iLj0i9QRNY2YkWrVuGJ
mT31NIWxp5HVUuTW3rcFP10iYFss77Vhkukj2kOJ+0PJc83yxvM/oEwhozx54YMs
ILGWMNffn8Nnjzz3It8Iw3sOB8aPisBdmGD4K4h7xsPWyneMMqKRd0sSnN+SPsBx
VeGPl56oGuTb/qSWg97p9ndS6sdADWNgTBHWFZU7roLxdORPP7UPVa0QgOX5cDNk
s6fp+wziI64iqgv6JTHLgLmMqPGjaGBXjIeBxQndtOimQJBhAPiU54Jv9dCCxVEd
3ZUSyTZ573G2HKeaX/rOxC00EBnNkX3X24b8+r1JpRgtBBJxiD6wyGgLFp46y6Ww
Dm2SZ/2s/W/jKKw5WAUOuG/C9cIIwIclzcHHSjF+2Cs7M1jCzTO41KTqACb0UdFd
rdTzl4THlqC5dKi7UCmTykayZItsEoqTfPRhh9oGvQQWTP4L1cQ8PnenUGITZz0Y
BDIfaay4Ig7e+YoLz9cp16ALJg1NFbRx+8+kW4qup+oXfl5/WRjJf8VQtywA/KMR
`protect END_PROTECTED

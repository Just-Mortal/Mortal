`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vps/NB5jyaVEDikk1hcCV9bTgfhQr8kDLQnqq/HwxJl4NymYBS7a0EvxlkqPicIG
PsUbfk2txKUnJ3wp98R7pTFZZeChpSZVg72LIkJcSgCaDbGBO5/xxbkk9OYp4F9s
azijCe3+AqgA0Hl2fgqDt/eKI65Ba32N5gi4CKbP4BpW0CTZqKqTWVYNG4l9c+Oj
BFEOBQLESxc/OfC2erVr+IgVuU5lz8gZVpkX3YlaCZkhtaBCpr7hszGBqHYQ3PIi
lFSac1b5EnBLjdV7Hsj9SDFFCHKM8I3GpuZvM40ZealVxGCRLnaiV/iMvcy+N+5C
XcgsPULhLLhyljfQgkgNPE32gCB7b4VgF3snj3shxA2tq8BFqOk0WPOJQzDG9T0H
1+d6xBtYEjmIlBAVDCLON/luGHTMSaLIUBYYY0wagdQpedWBNJy4Ty7McpMHcrw4
p9xq+CbY3OWo8KdLs4y7jJ54ds78Kizw1jG1FhgcCzyqyQyoDrXOdckhvUZaqvaj
xu4SzNV/jyBiqkHB4GIftmW+VPzSqnGCfi3rCABhfJOvEOXPj3PNZIPNZGWD7AJJ
pdA7tIIihaqV5qLmCtpB9L74lzM0HxNDEFMHRMUkEomx0lEwmxUOIriCrj1/5Rn2
/9/bN5kiL3U3gQtgngH/f5CMBojTP1QuVKg/+QfHyU4PgcnFJUe3u/DRlvz8savu
f6+rQbFH87GJHWtpW/i/Z5tvMHvd/xlaAsuqcTXhR/HutR5etlO0oX70qxZoU3f7
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMLKPVYH+5XQeLDAeqV1Wv0dN3tQVD+4B+cMDSkO9UVcjXjyMZS1uRyyuD6dOc8V
Md+WAXwOlLQ0al8BlyJCtbp6kiClT3RHzAVTykDbooKCo2bejWIqFteE0ChIfAth
XLLh7JyksQbT/Wlmor487O+oqhXR15k0xfPihvEWekVurT3Ryp5YMBFCDnKVC530
a9MecFux0wQKZ7v/9WbMavDBzuFPY4Tx5oWWOyAsu9YB6vgq7oDrU4qJipGjsxwk
QSZAb9LlqOEbeaJelnqpKSFuWNfiwQFRlC/cewzx91T0cbx/q7wUqPnsrFUydpTm
2Y3NjRpC/gljDcxmZt9Pg9qQeuFYfTbBx7I9LyyoL+EXSKgQqwdO7QVGCiPGmXMi
4E/egNtr+x0T0cgEFlfNXFe+AEhe5DBqjcHST4FWzfZkN3JvG8ZSOLQdcJbmNoaC
0jGzeXQSHD2OE52sY6TarfQ3bzXDYv7YFc97X1WHQO0XDmvghK0yLa4lQXseKxk9
WrHaxhQQgEKPAeaqpmpekEQsv7k/B2bncMvz06wMjA6wzCmGt5L8viKkoTRjwW/d
qzY/W3Eq53fuYMvXHPHJDAEQXQhOAZOblt/GM+dOmknkHeWw03FDViKYxnt1AhcO
WxPkeuNl7je8UxsQeT8vZUxEjvAsDK+AuAI5V5V8E7MaW4ZWFuUMm4sU6PKtvlXt
3kVP/b3TA61EJ+Of9Got+fVhNeOYtw7QCt/lclyau2c6oEpZaJJhzOc3+dmMZP9l
dU0w2osjy18DmPTYswBfnU0pwDDPgFKLk/3/dhdzeCjVOx5GvbRS0ow0Rw10WUQ9
WWKY5xGMh+X0wv4xMqVDVHyT3XmSArNMtv9V883T7GT9Um/qDJkCgh4Q3vhguBKC
qeBrz5pDTNIGGAm2fcUVGrEQ4NLUsZTt7SkqcP8DQFBFnVEBELgQxMWU1VD9Z3MX
BbjHkfZxxEIaa3orHF2+GNj2x/Ro0pT8GHcZieGBjwSwzdDmFyyTBszm29cVfz+m
hXN3VUB/nvI8F7RhGckH+Vbrf65quNdSpyNsW2jzLZSjCmgWAwRoYemQ0BvlWmcl
nXKdCEVfen2dDt4pksIqLE6L7bfPVaqfB0j1YPJ5hiwzahx6BzpP7B/wcKbVzwO6
HaYSvbx/YQao2PgK7LxlhmnjoUbegPDbW/aNUf5klQWZMvfF80MelwPUJa69VwUp
symRIZK1ZelPyQj2O0XX7Nkl4eekK3VhLGxDsEPzLN9Fjh0PV2jaV2GKlZyf9zzc
X7xq9nAxkOwz/+5qXROoL2cNnAoMKXGEq/tCLf/RyyE0sZkbf6j/zTri5AM3cy0/
zR+vxfifchRrFx+fipjImg+5nOFEVHs8kx8UG5LyhC578DjpAuIV8qVCvJwGmZ1s
XlA827/g4cJQBxbdqF+2P4FWIliiuUsRHziWIMqRrjbWuebwh2Ud2MctIQ6uFRF8
`protect END_PROTECTED

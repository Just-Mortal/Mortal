`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q715qF3OqycmC67cTp7p8IAJoOecLX1lBCHM1WnCklnGDJ1T5cQXUNf9A+l+iJ0n
u/Wz7w25F403a5cShQeq/PS8QytCmHfWHI8iWYKM/f4NU2Pb6YnRce0YpQcEbvts
4X9+05dNOX+2riV2UXmz5KVwUiZ9ptZnC1IDt2KMxy7uNBlaKwMjcomnYe2p/Iv6
I50dDzfY9MFrPbVZBfqv81up05WfBOWYlMzWt3fovy/OjRgawJc9pVndC7RGnKao
XLbbelQILqn+VTRhHyQiSObwTBwXN5HMu/wbm6P2I24o4T6NlTfPfijce2bNDthj
vsElXYLLCxQc2AQWekeUXxeanuJjjOrUVyyRu/tWjJZfdLCHR+82NlTye+b75q61
HOCLVuFeykud65j5j7DUCbubMjuxYIN8W64AxdcquqZS0JVY28BcLd233e40TrFy
FpEbuEFnvi1stW/J6ij5C32L/ryhb2Ks49/0mb29D+v1dfEGmCZSdZLN69RQ3yag
Nv6Mg+FI5iPsTx8s8owr+H/jJk0OHjw930A2UixrCQDgLDJTK/LnYN/l686+wJpB
NBnvzoJQsXLFb6DIER+RHgpA8egTkGfXoJXd+DCvU5imUO7z4AdThxu7c43Q6qZ6
6BqeHUgej6+lsaRU0GL95SPbVdJUAOSx9tDbx/hjyyQJTPgw60xN7uPYV7kVBNma
m/yPm8rvePsXByMPUIolYEmAnXzkoHHkUO9rOiX4nYiM9Omjg0PJOPtxIiP6rI23
MQP5EQLR8NEq7RY0zFZ+icJVO5+4ZqgVwHGlAfbmVFT/oOYNOK6Y7xHOOeGzCVHF
4bzwx7s+WrSYgxTIy1ohLRVgS9sGNO1jFgw5n2z9Ma3F7P3JMnrjBC5AFPc3gs9N
d9Gyqn3hZR1GoWCJjybeCLjtLFkH3qKZwc3JFZ8mW3COCZKEwWO1whgOZozeKes0
jac8dFe3fV9fQZOS3w1HRUAjtHD4FDze+ok5xq+fF/A=
`protect END_PROTECTED

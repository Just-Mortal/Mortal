`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4M7p8lRbcM+xd9wMwaiUaqqDSag7v+bMt8SxiKEqzZiuU1PFMQhjM62aXSAgoT3R
n1Nny0w3dJAnPXdPkZI04XhvSiM+q/WEkSLW9CCdje0rQsGzX5vVvmo+XglxIre7
oxAFK4K/qRxDSwUf76/SC3NvkxeS6jkhC5qsvNBCseD1BDOuVEI0zy5XmyWJ3nlr
JC1hqJ/Jy+R3osL8B8BPzyA18eYkZtE+wdxNV4Tp+1DfxMDBiINZBQTNNSoY1VdV
VbXaPEhyE2jaHIX4h1oh/g==
`protect END_PROTECTED

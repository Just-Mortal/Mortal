`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETq61VNPUd2f7/gpfEseGI0/XMb8BuZk0YsBCOTosuk3GCmocIGmRxB1xwA+0MKc
EPtYYaBUzrSFBCDd+T8H8P2PWM0FuLvPYGaVWMA++TO3QbIn9TyN1pudU2WR0vaE
YqwOG0LQBw2zUeZUMZI+1NTF8pBNedU8XXXBEdhN4xLzw+drqbeuPgmkL3NWcbur
9U5GMoF5ksRcWPUMGc0Gh+fZHf+P7Zlgx3bVWyeUC+eS8nq007y5lca3Ng2lUPup
2616XjQi73VkXdtAlT2dfc4GDYgO/VAkjPlo4OlwDdv93p+TlwQXhZiQC5ycBmFh
PZ+Ffj+3ZpQwOSLZ3fGILN1q4/++zAUKSREUx10PBofTP613Nb/sgZy6NLDKP1FQ
wdOMnqMIKdh3SjVSlTF95/ciyShZy49K9NBFITPROc/HWfsdXo0p5GkimTFavT0k
KwHylWUs/vSsNm68VvADiNRVGFHkDa+NWkO1QXKDk7CGuZchkQXw4uucOqADMz/n
Bjc7UvKhKl16hylE1XyyAUuof3WhN7aL7225TZl5qi9EhbkdoWX54YgMcZzHxZBh
zkcKVvu19h9aHXhCnMriZjsh0i7SbqqvgJNjBpM1KtnF+2Q5hb0/xfLJVJwVRW4L
rn85iHAPiJoPdIpCf6rgi25MaUygQqe1l3iH1uGMMqH6Dg/ziQAbJZavKKxNEXoE
SDA4aBvLm+AQw58aega6H5qxaMOrTelhvBRKq1ZQcmmgsv3X8bWcJKFcCuUGnoL8
4EZcSQ8Gx5fHy+/ERuNnGP31Cq/HH+rX1VgKGdK1KKSGhKw25GysM8Ba7gsVeU+2
30oOamM+iPwlofb02aPTvIRlG+UGeyxOK7IKv+I7s98=
`protect END_PROTECTED

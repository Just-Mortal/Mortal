`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vv+kvg5ibnBllzW56MojPDLU1fv/GpsiG+Zs8dvqagwNOwIDuUHQpxjyxzCU/0yQ
3Rfl3hpiJd59n/AXCrTQXYehiCB2SCeBPh9KltYL2ebipf98QQ5KNx9U714AHiZv
UeYyVk8P2dA0u9gEyMv3bTAVYiXQi0rQ+VYkkVt0tDu835CxYsYzaOZwMqDPe509
mZy+XRIHqp0tbEh5C+632cHWP4Tnlys2+0B3GSLiquIR7m2riDd4BmrTF7+nJagL
7q/3FrIqCi5QyD+yWuXL9I9NOMusJeJWvc4F4D6bwJOPQttAQYsyLJROoKbpKyF5
LmSOCkgUcA8dEhk3bJ5AVWfMg7G83Y+VfnAI9d5Op5y1QK7Gcy7984LZBcGNNMPT
0m2ts+awPkBxHea739Cj4oaP0X8ftHMHNn70ZvVgtvK7W23pU5uQk9RGD243sG7L
izJEyyXC5wky8Wy9XOLDkvFHuLC8irJem8nhU4XDtLDYnyhpoYaHhobPCBfnIozA
6XSaRJhZ0WU2bEJYxU3MSL/Q4Xbu0eFK0d9snalw/Tx1Z2EPEK2q19HzRTfDUatv
ByJXNTb221Yb/hdLDEAgqrVUlc91fEI7cwaC7XHomuUKOu4KASuVi4PhDT4BgK7S
2rNBgZZjmazMqbJfBEQjb7kPZ5eUjQN1A52OSzCEs1EV5VK0qO0tCF5p7R9FnImJ
i1kLIDr5fqevA8vq5OoPQEn8uMgdMATOGSzXQ1IAJQux9nm6Jphfy1cUCq6rLBEj
3L9cz/xys5LKxpHAABfnX3X+zOvgbxZrEg8Qfrt9TlsyU8bhlOiD0/zbhxO7qDws
9SHIdjERHRkIRcEIKm3Q3X+/ka9KJLtkO/NXFQDICvGKfnN12H5OAc1amAf9NLsQ
YBxnP0uugDdehCBVPsiqmMX3qUang9WxyIJK2Gr6YtZ5eIpDRqcfRc5GnSKMrYUg
4MWLqjxUExrvo44zI8ovrrNs465YsOB3lZ9bbyPe3QN9IIJdenX6H87gUAtgCByK
33/349bU26vpxNui8kTjg2vtgoHk/N2a2KKvUC4jSa8itu2rgvRYph4/tlVGmolp
HQ9IstHtLIcwCBNkdTGw2/KoZ899abK+vZO6AKF6ahfgGSbQ2FI6+bMliZdMzwFt
TwPR0UE8kGaEYXmRWHYRi4KUAoadvs31ATLf3mRWJucrh88hWrvANMnMFjzEahp7
WoAsGEJFPUL+7uXWau5iput9igNJViPu8rKcP3jQ61eCE3gglegU1LfIYp0hJftw
DBhCXEPV2POihlfC9DOepUyeVlt5f2qxEQWIBHF20opXj8mpzzChYzVgbj0iC3DD
MNYehQ1wqmnTjvE4KmWKTqJ8MO/SRIrIMSEFaahSseLcE0acDa5/GNaJzXGAWvXV
qSZzkYKm3BSlNXztlTzMg2rZfkfpZTemiZo2+8OJlV7o+IS6Qn2kQiFB1ZzXqwov
khtKZtSHuEElMLT2a5fs2yAOlGAqccCIuYsa05Dtk3B5/KGU457zU6tLeFSYoxaq
HQLmSxuBPDrPjXJaVUXDPQr8BJbQnP8FXRdVrQU/UIp1FmtQv8ydE4uGzG6AN0/7
YmYGfplIaMGCzR53HKa5LIsCR3E0EX5PSwxdV6GZiQE/ganKlM5y+LCOmCm8T1qv
9t1QAq34rFchMkwxPitoaEMFBdvDXb6nACBvapsei9Qz4xVVDSLzfzMK+HQMB3k6
46SNVUyicdzz3NVWmk5GzApNt23AvNbOas64qDefJZrEtfcgCpg6xndciIjU0YqE
J/crOxvQNpUqKHodasikd8fWfXhZC+ns10I5hygWes62bG/an16u8dixE8jPelbj
TygPYajkug3TkdlKGy3QAn+5uVNVHO5sUhsFE12CA3DldTCerYvZ12zjTP0t312W
N/+cz4vIy6fMystoZtWT6GL4UmZF1+Y2VeJstPkynAZaZ0dN4h6HLpP6nEnpKOa8
fdH/e5Ggw8W9sYg4vdewUZ6QzMaj/s1RUaPiM88nmKz9w5+vxzBq6HvYF92Js9qZ
woKDpbmgaAMZeORhhRfaUFbA0c2KZpjWPdsraTAEpFOVZvghVt8MULip0ekaOy2R
1Y+uxRZn/DAB+EKXEAOZXA3UhoVJp6iKyP9gfrJHoz3bKTV/saZaIwahISM0tsdE
wvatr8mCjBtL1ywkMdISW9qDsA9n8UxECSX0dBO9TnEaaSbeqGDsN+8LdWV2aX/M
XkxL0WIcVWasKs7l2m1Eb+057zRtC/BHHkm4ubTukNL0AApQISLMbZbxtTq5yr5/
91ZSfr69XEoSTMUg374n7MkFhyg6Nt0nAkMEn0cy3DE3uBDuMd8aM1JUTJhEcvzF
FuFvjVkdNdpP91LRDJFSN1RWFeYnta8Wta4XcD+5ee0FGbjDTCvA4WTij/CKhug6
CV/IbisVb7zKGQoa1swDlRzIwuhMk7p1oMNGqAKEuGUhOInwBtJ8kq9oqSWnHYHG
Zvqd5KeAsXNNppQ/TaWZdoLZ1SfwTFKBBSZD8payIAQv3nNo9Bs19vWMY3DkctrU
T+V12vNeJwFfbOJbxyioWDzxUtYVQmbZWLjGgqipCsJO0L+PBax5VWLNchNlKVSR
Nvc3MErJWSicKuVMuPINMFD+aLwDwCckayT7OPlp8+hewO3nCx6kpnnGYKiWZjDN
h1s7d4Tz/kLKlMMFdzoKHW/o640Bxa7RnwSr7qJvYXgEqOtR8NkbLaqu/YKDRN4o
SE09Dlgq/OGr0I15NPWqwjl8PeAi+wgQo7rSzA05pbx1HJQgRqY+wtxuIkNNeGLg
cp/IYGiLa+4y/6FB9ahirVo+QTgAPdOTjqaC15Wb8Ix/D95V/hhHRO4SpjOpcEst
VzRyP/kZ2NW7z1rwcCZSbAshTEFANabUNleDFl0Og4mu1yHeCJoryGMG8wVeZjL3
fR+vHLcAv5/y60C3ofNFgo7oXTu4SKTZ+CJ3dfx+tv6DEnzsRAHSFFjHNp+uBmtn
oioPFM+qhBKqp716zXd4wFELwk7H2PYjsWMcHZkbH+1WpyinSdHdOWkwHkLIzjDS
SV2N0hzWjoYan65ZtUYP2bq8ooImXwHUagIPdhqb7Aq9Kb8e84BVbT8XFf37A5DM
dqzcebXk7YKKRNZqeiB1ZZezQJq6tXZa95BWQytMnJPqB5OhDg1Un4yyemUP9WKc
Nal/6DCCe+evw6GmQRxSrNLSHLt7YVRDnP734T9o/0+AJgSUt8Rbnr6FBsDxkU4f
Es4ALr55F/YeSdRRu2doP0KOyVOU6xZfYjfgESh4K+rIl9ahz7lURx8jC/LFhG0r
A0TlMAzoGTAwWsZn8biFe/bxphRHgFmIBB6XCxA72fHJxMAQsT2FbVEDNdRLCoIB
vpCjY9UCfleulyCdrgwCLhPIFJGmvAO3+J+uFHSwpHPQpSBHEhOR5DlSjqgsJLAg
scACvemPsXHytxi8ZaXuktD+O6jw1+2bgUhxog2zFgJNzSbEwX+S9LHkrdR8wo4u
v1/q1jTOnnxnZ2huJYCcIyKrGtIWhcIeqnIk8D3GRrN2jFN+51EzZ2wv4ROn/y9F
7ePzWVoArOsFI1vQCjJ2AdT9BeJO/w8UMDKaIVmIiNRIzOIwSyO9P7+hCS2Yazse
EGTvrORYBDkX5ayvdGkHBryzVQwqih8vOT3Yaz6sv2BSN/1mi2C2h+95M0hx7ubO
wOXIi50FXFA4FqBOYIWPKffQdGSoIGYIlDdHaGL6GzFkb3V+c+4EB0t2aQvPpY9z
UM2RVtMrqvGl4cOkGW6U8aWK08GNxIxwqsWaFzzHfOW2SubCdczevNZpQQ312shC
HswLaB7VUSqsH/KdUXTcPhDAy+JsbVt7P5A3JopYOnWWDu7MomdQzlrJJX3ARJ8e
JgoChx/aDEJ3jBsnd4kLqmekR3afv470GoQ5yogHxBuUQhF4yv4y6rbdlGzAoOJm
EoMl14UwDzqqK9xuUAtvovLOyDkBhCHIocUtHGAO9Fymgolmz1HCMtJwALeljmQK
UbjJFd9B1sE6r37ccpG9omwNQroUGEilia+KbHX0y3q8QdeGEduCz9EsBS2q6CMg
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSDi47r5a3hRiVvLK25xMxP1jsKicceAIGVNzCZiH/KAum70wcHoAeqFF+c403Q8
kZqfkU8SmXZqBTnu+so6CWQt0cPAXxSU7GACXS1QyxvUUjWxkuEiBzPgqNIX303A
ztCkIu+zYesrIRAg0wi4wahHYBkeA8iQmxtgRGgmv54rK4wrcIrBNj9Yt4iTyXCD
iWXwP89R1GO5zd6TnJJvaQwf3rZjXNcG14QxEGxCXeZcS5reO08AOdwNANSuYfAF
KVw1fdtJ4wCox8dW22/YTgXm/2Twg3Y83xKgzsVymb9bbedd+27Ejuyz2gDYG7is
rZwGM6WXpWwB5t8YcKm+Ue3ubBBglhJfXVhA0ZLymcj7phOGWL3c7X1dNjAPMlvg
SqRXXsD03TO0jaOmeOleaO9esOJFVyMYj6xgLe/j+A4WN5npn2SWLquVvk8mB/BC
3rH6ZApBrv8wq8oY//w4S4H2Zpl6okKHOj7G5FDy/ga2gRsBZ4XeAcSlP5JQ4pIp
vUNrcZSACD/gjxpAPC7DFjxE8vYoeKnso0ViX0HHtDjNS+51P3pBXY0ffLLdtjLr
MDJCcSJxVhu+M4iIWqgBmZRiiZYi2Ppro0aJ0YsYbsBp2mIh5fPMv0+CAC5+Y1QU
IO55ekJimmbJRHqHyS/d/DErwFplqaFgJ8y9+8kCMs/+DcI1iSE999txnBSCkSWw
ofpUtYv/t5cP7KOO7YuSsA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E7UXKoK3otWTYOi44W0BpxiFBgMscX1HGBZiZMCX+MfoW/o1uF6EwZLuyshsZRGV
gz8RQRwpgBnKn8j4xYAEcXrEJq4k1bsnNYbBxaMHjugi3HbA6R+XHAFRjINvJx9Y
JW/BHQibqZmGXA/yb+cjhMMazXb+uXyb/olk9rmya4HxJ90N0bdRqiJDxvydFERU
t4+N/nnOSizhNpwUHh0mdYiUKwgyEfjp9dc3sPzLRJNTRNwszADv/ZvrllmMKOJP
PRu1su0Nbc9eSXTsm+QRI34A9ilzTVYYI79foIKln7HWuTtZ1v6A5esJj9RmUEaJ
YAJTaRWqA5WgMVVowINTmi2CgFDweOwNc9TbWnnc9j4hnPjOUWNZMZwkVDmVGUH8
axptnT0NfJck/DzrLcUBwIvhQZ9xck3mF7ZWYa0FxOOALSZ6qt4VgjlzcY5GdaE0
ub769jTMhhXVNd7u/Y5JWVkm11Olhi3h+otJOrrwyKfXwwOcS/flgoHPc1QpyAs+
M6e+INxWGa0vGg01gv3bB8em35/h4bzJ7IAQ5sahdetU4vDjDgoUgMOU+X+vNkr6
8/ffBy8vJ+WDze6+iMfBj36/Gm0rPcXU4BnoUUucVwUjUPHuleJEQn1KpDB4fUYN
EAaQyAKNaOqycHLiXQLlhyLDn7mHwNo87UVgENIAW/UJXmwtfiZLqYs1gW5Kb/Nc
b4tfSP4qmOVyGhAj9U5Ye1m3oMAskKHC4U+PIGmZaixubfw7Khl6/nbaahSOx9Lx
/L/8nmYvMXjjgcRYgJofu22yqVoGS0R7xRfIE8g5VA/Ua/QEVZRUp9z+NkgswnrL
4tjS2PProPHBTmo7nU6me/l7V2kEo3c9DvjHeEREt6cVKCNVXDkEizIT7nTfFmWM
3Dz6XAg+Rnf5zNz4ra9Zvp+p4n/mNT2p0QTE+qC45Px+fEoAp+IHXh2JkchYPjDQ
j5u8u3jfv9+cvymqLxl/zccgQjtNRFgsl95ZBt6gTLNiACnEk1YAH3IH31gq2obn
9+guf1Cb/+B6/8somZk5FMp63Rgj8AFI6DbGF1WpF/CdexZnxY5GMlOhAvB/xSe+
N2PEzfVk9Xu+PvoBOhHLGV8Rb3jBLylO0c7IOc1DnxA=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4j7FEpgbQxqXkMsEZf4hgCbzsBGjgK5564vMiy4eZWHbL2ezmz6zFbkG6soJWKuD
uMsDMsTbCjU2OnrPEVo4NMgpyiafGIGwGaQVcMybPQbYuC02msU4IexJKGE4x9F1
tOGz52zlYUPlprG3T/+urs0n1wZQWsIglBlRAFVy2HpdE58V4JdBNv9HPQ/cvhJJ
Fck6WxBrDTXYycDuoucHf+RXfHrM2OzNtR84Y4+6xybcBCRygxGOLGi4+JvLNx8J
n8c2dio5KCOHkfVsS786QtXnVJr8mcZeJPDRXmeuJuWf33ZvtN6f8j1jboEcy/2d
QGvwGGt9ntDBTedDcZvXgCNirq0midmjPnNGYNxwqklySU/6rWLgjreDjeLI6Huy
u/RoJX4ZxuhbHOamdV9OiPCfa7kPi6EsiL+y50O2ksoYt8s8XVluPkrJcmGW536y
eMtWJsSbIVhPYIl/77iNxu1ATVbNXiIWewWD2El+oU4A5THPQipv3Spx0Vqco/Un
iVYTCrA7uqwNM29/BzSqUMg+R6hzs4hy54cEWriD5ZmecoUPXxmQC/Wrv8OSjmsf
+NQO1yK62boytV8oC7d1oeNxXTVIyIXfHZSQ31e0UdlypNzzM0K/QKdHlDGxJWik
w+gLJTHxn8XoTnBfAD/sW5zeTQ7a0OFVxuPaNT03oF7h/Js2+qsmeh/M/0JAhB4L
oiyjTc323IbwwzP4h86119VHjFPaeBocKtIYCzbl2CIMugVG4W5cOJjkNa490kkv
3ahaKCfOj23HABQ3182bzWl3m9clRRzfQ6DKl4GRq570o/DI+tlMy/i5hgpJeBQd
bk1ezFP1vaURdGiXOhNug0VvK8ZFa/Z4bv/c31k3GckXa0cOKK+tJ+KXmPOkeP83
08EGsgDF+EHqKcrMByFFACryFCEnm/RHDu4SVyNOkMgcrmTIfmEwVj9sGlH6Qi19
BXPsNzdfF3tVVEpHfI4LNep7WAakdOZhBoQ10bcdfrnHYZ68t3xa0iEjtLNqEzXy
Qf7jbKGRl5Wt15Keqr7vJ6RzQ1dqNd7RfBoyKusETF36GXvvPP3WGuGzv9Vieuhs
tYx5cDUgaKA/qu+8slMnwbcvVFv7SRJHBtqrDb1f5Hy9lzbmiLGN5UB7SeTE6wWM
FRX2n2euOouKMm+oXFXImWq1FeLZWPHuJR20ZpiTRjhLGOXuz5LNG148gpjVHVR4
x7tzzSPWTL4mDtadzHjRZ/RWhnchFswU6IewSonsBCapczr0SuW4Hj6VzqoMafEN
O5Uu6FpPq1ggrGRGXTwx+MxirlaINAl4WcRDWoKLM36bPhNBXiyu7W2bGafco8//
/ohyViI4phJ30S/P8hjaA+JFL9dV/yLsxaYPvotQSzuCyyzAoQ70bL1E8gCNLyGf
sD/KIR+4EZepyQznVeKBOolDDsPA7t1QiZ1Dyg2HMaJfaeix1OOn39h1brYlIOG1
pjibLHMfu/AgGghrob+hWCt9xvSZz+8iTpYrnyZeAn9XZX4Zjg80/yJ2VFUOYB95
HIMforjtI2AWFgT2QNn74HME8PXaGyUy5nY9eKN5LvopwgFbr81BpD/lQUEUnZQG
Tkv3WjVqUNwaOrv9KbXUKaRqBirL1a5PNpFtdWqp1UqueyLmm4McJaoy+mtrNrti
4eT+TuwIvTEoNHtKycDGObkhHdd4SxOmz8vdf1PPcywx6aKktqBG0R77bPqvBKhb
NIELZx1oskI6C6KGOBhfiHKvnMwfqHedxvicSY6+2sUqswcDNADetfDDwlot0HNG
L8TiuMSsJL8ymbHo9k5Sv+HpMngpfpuIni6tnBlLp/ZU98DiDi0dD90iElARuwzy
9yxuPaePuDqski9/ksnI8hdcf7RjqkjjypR54fE+XI23Ly9V+O2E9vMQO52HBjY9
LPFZvpNOs3+9u9mKAjeV1vJ0aObjwMocBSuCNmguFHNFIX5pSIokt+reMyKuw7Ex
FWDELvqQeGbab8SKWjLbSmF4Gpt9FGELG8mPIp2LoSSLHGA3GbCS1viJ0FhiTHLE
ndmsesFHeK6igZzdUBrdRq8a0Z27KiDlSY3+jWTlxkT6vbb4xOaY/ZaeUQ82miqh
CoCsb0ec3ObWbSAJh+ec1i8PoBdiB3B3TWIYP6/4O6opU1p+YgkzVUGN+0kMxcPR
nVTzVu1Yl/TLGD4Qn+dmnayaigTi6RdYqPrNDQwFNIbfrQHyVN6z5QkxxkP0gzsZ
eBDILGOLw14gubg73K96gG/E/KpJy+ClAIFSZhmZH0EJOiw6GcJdvw7wbHDQDesK
Fn7EN0nYoMKH5RwGsws1W8i/1/+IAyrN3k9KQcAdACnPUVyIWL9fvbFY/ZHb340J
pN8peWYBsuPIX0Xkv82ohDmRkCFotlUJoKcD2p+UYpAoP7Ij6tDVHG/IIGK5dnAT
5VFs9LUa3K+5rHxUqVfJHLKg7IDtqyiuT7eZ4JmIyCHPMYQPYVDj7omM+UqvvzfM
B8FhSiUL2NcXSvdjv3tmi58q5bQkgCwRETbLsjKyF/HAo2zv+NKP8YieP5HZgnPP
1Ed+fRXNVFRhLvokhw24UMeTm2z8fwhhYQqrdN43L2Tepv9Pej/uXj0cY5uYSptb
SUaq+dj0hjskalXopvRha08EtWiUuEWuwSSgIMZtSkfGMwCwMyQ1M/j4ZDT2P3Pt
CJFhXnmYqRTdbUrNMTSrZicmSfFotj6kxfuNhJw/uvIBvCrayG7vs7RD9sj22xiJ
JybI689DHkuUk2nO0LoXj3P07XXJiOiNCsGq355SAe/7TidvMMKnI9FOH7JOPKqt
zJ+n6cSaWA9f+ap1mzqWgn7hBh7P9VKFdqpeO4TZfYexvxc8pc+rSvI+xQvm+Kwm
2rg+qCLu2GxtI1ONZ2LH2MtvteR1Hx5wqQ9SNf8vZ3/JofhhAe6Igl1AP8ze+AJg
YVpKmui7XMWuoNFKBSTFu3YDsqfQw+TEdK8K3vui43p25bM8FGknPqq4bZd6Pn8u
qqXs5fBcwkDYQX+uHzvrBzN59n4o8lwKGa3papvLYOoMbmn+pC+AjoplMfO/W/gs
dL+srKqeJiHJBYwSJaD+fT++eI7CsVNfX3XAqlZKdzsc3F4RPeX1JMDQJdEXdR16
GHVupQGB40oqF3GQaHe0egcYTO3axppr9SgyIItZhLT76qmpZJS+MAO+GtZ+hQi8
UnsWS7tnbkdn9U2F88TYdpo57tQgAq48T9Y8pWJCOt5j+4mNLV+3u9rl/FSdN9gL
9ObmT/YEeP6VIrwNkYy64JFe85u7wH6tzsw7Yyv9uobxU3jcXtxlEqCcnhyO0IWd
bMuyoGp/92EGWetqD0Ex0+1D5aFPU0ra/JDOmmqCska3HPB3WtKJXSyego2uTJVa
EN9X2XXBmRiza4vxyj1WQyYcZG/qbjtLTb52AIPRe8UJyCsLS8KZ0Rg9H0FtKxll
thtubDHnDdlE99UicPps0bd3Cd4QcC0bBTGZDdLDcCk6v/J5KfTK+VV1WRbhWxRM
jaQJLBdcyZ4vUW2NGlfn5tCE6QwyC+qbOf3YX78lx8pWQOU5Kekd3SC0yRuFSXsC
XafLQmidvIlVohFgceks0ZlTIku0FoPiEbi8ebh2IR7MpxLLkjlZ8/ZJ/hv5XsBo
OOVDLxm9GoqtQPCMx1Xwe6LG0Zbz1xXMdarFotSSxG1xEViXlVZeGX9BrwYFKT/7
BYgEXI9qX+NJgFqSfd22BJ6c6NEViTHprqkDTvhUtNuDaZkbCoo7T7ClEFoiz0ym
7+2YlHUapWGP3D6cnLJ3KVtvjGI8Pke5HQeBxLCmbTPZTcKKfmbTgmY9AXNalepT
LSG1EcF5k8WcKT7/CsOXLpByr6Vq5HWosBHECjHzwmZNyEozJbDSO9YncFFKDkXb
rEEmuVAO7VnjfvVy3tJkwyypWmq5w5UJzGKEUYF757sa3S2aaXl3a7gqGgU9+bjk
wuR7IboPW6y8M4G6c5AoA+lKDg0UOzSON8olYcm7hs6HZ8Z322v4qOz1trUyGIS8
dQ0eiAs7TgMzTI1Sf97LfTzXoKrGlGRKvUe/K2KM9r4nGy90PjAB+4qIXRkRriI+
HPL9tFTKftVY4cpXUYKl3HmwsiEfhhL/Q4Z7HvG3FwM0CNKbHatMsUu8ymxclD/l
7S7dDsoJxw36+lJCCNAn7FnLRDIAkSLbsH0ls8iK/GEZ2FkHlnhHY4U/nwv5xuzg
YxLu1tiSUw5NdEvziFWF/zFkjym6hQj9J2wsxSF8KHen9uqVL+xoAc5rg0Y6WR/t
Myc5ji0WXWXogaWv7jdTpDJkfkw4IrsVHyxExaNkvtzInCAWmjyzAZH7QP7ERPBU
6+RVs4BL+hkfpy5JVg1HwsM8WLBFQMLbhBGdLcHizJvq2s6ct/urX26Gx0BTP3a2
5/5UZPtae0NLrmsMicPECrfB7LlYlLJnKDiOHHJ8YovzVB/M0PuvFpNCLOCGw3Bg
bSGmToHUouJ7v5wz8Hj0CLcNj3lZRaGd6yN9Wj7f1eDE+xcQORLJVq7E3Y6R5bAX
6Sj4HoS9yY7d32R/XcDxJbZ3kRZiBTIDRBCi5903ZZZMGEXaAMxdEDtf53aWEgUl
G0mc96FZ5v0PmUHDiYelVV2mdQRuK1zBYY9Tm/XFAyB94Y5u8EdJIjrMYmvFKeeQ
c1ZGmL6tdc4/uc4fba7miCRCtz4QoHocG2xacy67+tCmXrsRoFotFyA6dzFpi3l1
6lkge9iUp/RrSYIKqrajKZ6Q+DfdaJLX4IoOVpCxyzQ3ChwxtDjVUI1i2Sbzm/QN
JMhpOYZlYN0U6KDVvs8g0BCicgxB6ccSVgWQ3Ya8JhfrFbxymrUaimBpUhVE8TS3
hrVZyz1RwLiJnSOFWYOrsOvfMuICW1tZcZtHkr72BVL7b3GiIbcxTGUYAukfiMzG
sdT/TbqJ4DxZStysyZwD30zwpLgTDLpVyxfG6DkG99VJKivQmp0EvNCKCcl7LJc6
Y8Nb7STfp19IrQKgYknFMC049LugAfN+KjbTWR4gWoxQR+750lSUJKjMgN70IiCU
4+DbE0Jr4QK2wLzhs114ptjD8Epq9vTkXm0mjtjOPSM5wXkwSbkdK9x1KN1oN1pm
l58svJcjDZ8eb1rOXLk8RNknyHRoed2Jkb+yOUrqUwNOjShc3P5O7qo9alaAlphJ
kjoQ1R7rAKfB1FC+ZrZ/TxGpY1BfOzKxXoSNf9EU9/foNaX62Wm04j0SBsh44v7e
hNp7bNK2WSfRamPRAN63ruEAqtzamsjztXTZs7+lyDdSuNccmA9RTjT+UvKNNJD7
gYul6XzitAC0UBzhIvUUCE2jrW6X4/0nVcGp7c2/Uh4ajPQL7A3uToCChK31TU9+
OGWFGtUlA5Eb+93sfoQQH/hI4jngDWFhuvcdAD0jEUnx4D5aooGF0oWnVjaD0btJ
jeHuNg/ZNg1EoLGxTN/WJWePCe4i0e1ksm1S0WBAlVFiUfZV/nrC/LwsVHQB4uZB
6xgUfxv0Cd+qENiy33k8627JvEXwoHipqTNzUq6UcdIy0mCEy36eZYL0TWRgrkWy
TB1urF8XUwKs1juZH2NExY0cIKerw7X6H/4ztz16wuzI3HW/AfmYVvfntPnDE/ry
U0/m0aUN9RCS4dx5GFUgJcpixd0aHwv909+umIYzNrP9NzrbYLjeg1mpOIWuFGQt
8xG2n4ymV4XGKfloleh3TJB6/kjLFJkM1KpUcij9eup39yJuKzAGy9Hx7O6j91xC
Jffi0Cfm1hmGZrgmd9ViIpzd0UBmYc+4NBhupcHGIk0hopEEl4MBpxeoTDFukx5H
Rn/v/nS4ISFgG4vjdJpI+u14UXl7EqhKgtuU+B+FzdlSXzzpCtO7b4Sw6CBAXzA9
MqMqmKLVbXkil7IspiBRexuNYG/lMY3VBULu0Lqv22V1KkCETn/2TLORpQlm6kO+
s1WfOLT9C4FtkRWoozXuINKyYTm54AYI740p+wS91p5xeWQFrW4htkCV3GrEB91t
Ei+FikHIaFAnkpF210wbKY2kYk+zt2LUQwpd7uiAZMl36TYK4nT19ucWyDV8MX0A
XPe+DIWZs+9OTdn/A3dow6SlIVKQgb1J2+26KGlwPrP6v0pG/Leu8WjiPjLHcGaH
R4pK7eDxkx1VWqN8XQVuCNyNnxFvwNJiMmdQXD0enkwDk7d9guCca9Ruy62nPZnA
iTJnn7YOf2zjCD7mgFnzh+/kdYymzvuM3eMQsRmlSeKNy2BniZf1M6DWE3Nl94c6
9Yeyen4uWiSPrlylVi5HZ2XpSV4M1rSB7H6zkFmgCAqtziPt+FLzLHVsxnYRlh9s
efDjV95PhsMyKb10fCTtnetCDndE6kmJP3hImf8obXoZsioWjlDk43fIXMPvit0q
iBBFm/Py+cn3ROyRfMtFyeHNGhTG3lcwZYFI5LBKHl0wODMAMMV26j+aBAkQjwFX
XAxkO27zMVoZC4vBxSKJpybVG63r1rFz16P03yU07Rk5tfLbX+m6oY2BH5wfGFqX
McMTYY/SkwcLCts2rnfobnshsDk1Cewl45lJWWjSA58XR7JXmpNptN3UiA6ZX9/t
XOVwOvMFEdVrOi4+/sDra4M3G1DU9Beb7grPuBxTJL4UPqE0rUV73AVL/RgFGRcS
N5MKXD6fjufI/LQ5KO0UHJk59AiOmMoXFH9kmW4CFbaDbSXRDB7NqcMq/5FXDGHe
f74xPn0/wFf1suC14lYXvBxTyGSTYzXwsChMbv5iOE/Zev9oNn0JCgd0O1xMji93
Q+eNbAMS0LdSwvm31lcdTXhYyJzHBjs4PrnRHFPtwXSOsobnmhcoqqbAUx2XL4Zh
jHJClLgesYgVwINnetZ5JUEIAmM6XSUirVvpI1z1Q2bVv/bSKccJVVXC9jDa8kDI
TfJbYxsO0vn3K5M5btMzOP+9eTmlqORCJ81be+XeM9MsdNRzMWK+vEyHrJ418LKF
ebNYRsOIbzEdMEK2zHJmNYhCLr/VAm/DHZ+fIK8anjKQoMPZhmEgoca1jLEcpigL
155JlJxz//QOB6MYSw22VVZLxVkg6LC6PpfScyJOTfp3MebPBYr9vv64ud/JzVST
bpLx/oq5Zqesl7hOjMA4XGoW848YfKuPfHBxgdq1tG7dFSA5SSYT4bF57D9eGhKr
ZEGrEfei2dwBxMYubyM3hznRnam1qcEOh0DJNKc43SWV5HTBFEe5eeBrwVbgVCTh
5+MrOO6Got/MCGSkxfy4yKjQTdfKmx6hOPl2GZwXHwE2Ij/O9A2JO7+L4Vl+PEl5
anN6AuemVo89MlkAJ48tI0xL4x+cmpJAQAlm/DYN+asR7o6mgvvKJ9J35GJMuH6K
U106t5XD7vZ2M+Yhe07/CKD2ybF7GSG3EjiwRSIa3GyZ/Jwd9iHU4vdz8vCVmYUl
6zlCcLosoqXfIOeldUiw1hg9NEKjeHnouXOM8dvTK2fwrzQOI+msTEKcMijGX3C4
PddKbWJ0ZPoMXlxbsx8WosiM34HT8nbETSx5wmKc3K1wcogeenjo6+yZgxUVgHj9
XQsQr+vcFS07MKnlxeLAaR2/hws8u59Mt2EWJvq3bAoCIhC1GMuiwQtrfhG2ePQf
/+dzNCPRPE+DW8hGF9amychwDz8olWzus/RC7YXXEn4JotK1B8lDtGQZ24HxYieG
NQisC5A0HLzUnxiVA0c5cVvw2itp21nsh3CNnde+hZsX/+iD84gaVP3Fu+gKViE5
66IHHrYh7jNrnXzFiU58XIJb8tnBUCPLhYsR0OVntbAW+HA/9oTzHSU8qeTMwkyp
oDTLgTP27eFBM5pEepH2bk4tlHU7y1mwwtuV1N6PQQosb8J1LQnzbIBQYGU8RZCp
JNn42Qpwh7E+DLcAb0GUGwL+nvjMRqIE1uToBduKRvkGDWWhVr80bZR9rjek5hJ1
K5lDTtpfQUbyV2OGT9qB+6lCiv+h96ElDTenFHaMN8SuPZWJYHkf/SWazi1BopaC
XCLcLwYPpFs3C9Gc2npnQZijSvcK/wVbzzFXT9kwxHm/N40g8dWJgzDNkY1Ob8A7
44XdzZTw1AT4WDCb8Zl/bxlXdp9vsdkum+nVcjvgxoBGUESOW5l69KDvrkCdLY2d
6JLWh68D97Or2vFJ7ja1ZfMtH67EonXYk28A7i9qSJowC0wdDaLaXiN/mfRq4lAV
Y/T1JtCmEZa2+UfpBmGk35On82Udc1mONrh2r8Db/ockiwoljxPKF2ipx0MymwOm
uV4DnjwwOfgqR5IslKUfjy57YHyOHfsDYmwdI6AbaDbRlRvsqFvkW3G/gxXNlReC
BGgE0fOSzpdeg4uUbcB6v+vQs2VjFV1YkPY9xhrX7jH6BHHfI0TuVzRKDw+PC2WH
rwEBdB3rsPQLRlY+olIx5Lu4QSJ3pBGzN/qbAPB0zfCY1iGrctdM1rtobTeAGU1e
Bf/caMnO61sNH8Dy39DoV9oCYvgXsV4VJ2vJ+wTZgb1bH6FePqz/D37YukvpcH+v
xGIkttBTvoVU4o1WnsXgDTwkdZbvRxlwW4A+XfWdHDj7fcCUle4ztindaVEFl9LE
Tnt5PQT+Wr+7Pg+4DC5wwDw7KiuvdPUI0oixK5d/XHRHnXmb4GeANTeQbv5icqA4
3GDfNK3kXZRsEAWXXpx16UQ5SUjIedNKLpdBclrwmqey641fqkBCpGl+F5Bac0hb
iOWp7xwKC+UZpGqTpe+pYNjs53rGjnJ8SXe/nGB+UGXjEnGsc9t8tzeovQYq+W7B
ZF4J8S9AEiLUtsSfefE7Dyfbz8LC7XBf/ZxMNfubYASR5PAP4rR/PZZlVwIhQ5Vn
P2oiayvzc9zdJrNilPszIMwMLEQUAYMv1L02MQwA//7ADoqtrbQwxB7uqkn9tS6L
7VWUAzdhTTOJDAoJuP+alYtkbPiyGRfC7yzZO9AbbBx6nduGzLT2JmiXa8//pJ59
7MgXugPgdxI4J9PnPRMh9cOCEMrg1lqRU1kd3bzcSXOq1njoaTsWn7b51ZVKgn6G
JWShjHQ8TwZAWoKOkKANN4Bjda+lXR/eomZd3Pnsnz9uk3ZKY/SL6GiYSoxkZt9z
Lm/qvTm4tX9s+WMPhVBqrkhipFLuqoQlt90UIUNZUrA3m1aSPwOWa6QF8WTcoo6g
uv5D9tB3BfrBdra3aVuCFFJkKDy5hdduF1ZQu2ySs42KVAmQWQ/pMoNuTUZKKMtC
NplMe9zJIgmxx7PWxWBCoeo1hbZVttn2syDuzkBKMCKnhQhqLUPCImvdHHmf9VcO
HletS0NfJO56DuMumFl98+lDdBZqMlwatDvKNXVMgICoHBhz/S9APBnfWP9g99Bp
LpjAjRNTesOj6+HrzZkgau5/z19LfYHwOoVom94hVetzRPg9+MTMfW3u8BrHFyP1
PTEL3B/4WiKHCUwYC6OQRff08VSlTWFDMjKeArtsuEz4Y/rgbk0WjdBpKDjotsxw
5sMS5oR3MfIbu3uEgTKv+45P22CQX8lZDgzUNtmSHRjCKjMXjYG6osIIDF5zxI7S
dhgBzfZ1fy8PYRmQ2b9xM03yg/Htqh0P9LmRtDIX6J9zKnmNlBOmZ19PbYDemhSY
JSRX7Gx1FRG/5WjVIC4hNIINH+CcRvxh9QB3oBjwKMB9w0H1SEtahCb3pZWGPT7D
VRL3OTRHY8r547u4A8AYtDM/cY7Hsd0l3dVBIQ3wcQXDWg8r1dJ9mbUctdx1JND7
dARj5SIdhEvE9rFrNX8Jrf7j71+JMIW5B1qVIt++YSO4ReMzGNoKwRiYfEoCqJd6
6mhpse2wGgsejgAK2gIgOmecdwVNMOrT7MJmpMB0TkfrMGXfsY3sw0lOJlihj3jS
hiTMGaXM4zrP1B9ILJINTlggZkujYAiCiJO01qrqCmY/X0/SVZPOGT6IJwYS/FmM
TnMFseipL47b6viDUa9rBtbsn4vvsfPDT9M/A6tuESnEoxnyxAW1X1oFohGfRk0Q
E1TMO93o4oPmkctvc0dPps/K4waNww3cTOxN2uw7y0rcTzz6yQo3KzHTIlzdecOy
Ox8hmeUsC74mkWuSt/IJ8tqIvw9L0PZf8t2MT861jv5Y52pVJtcoiA+r32UN210E
VLt1o/t2529QNd5UcL2Fk/+EkZEQfSzKt9uUNnE/JbMWymIL7seVvI6NH8hNNTaI
KlbWFon+hilz4ApcRm6ieQjE+Iyt/QGIMJsZuFJQ2at5LNY9iJQVZPSUIWTO+1YL
zyOnxHPftItF0AaPOtBT8aBuzmPmRPEqDreGSVsAJkFOWIVj0Nq7hApSutWba5ix
R38jtbZ2HQ5YTF2VzPa8qfh6SBLNlEgMua2UTp05vv8aEmTdJ8rs9MpiACFQjIZA
G5B7dCsDqi0ZIOEflfezRS8QQwETnhVK3ht9O/eW8qnzTT7x8CNrQpc10Os/Lia1
U72boRBB3p6x2Z7PHvroxRTx4aTs5JjEqym40ShkJDtXcd24Z/0ptKUmD9KrPXts
QpG5apRjdQd8HTS4wGDC2ThGR5Uv91ZtTCnuH/Uc75ozP50ISNV/92nQKWid40nU
du1zLQ6/EgLypXmdee5E4bXAmUM/3b5RXTnIVp9QPh5QdnRYoeorL71EjPdMPYHv
tdU83AQwnE89K1YsyXTuZGOVJQr8qpCjg6uLLjnfY2piNqE4LRZ/L5I/4kU4kzaJ
g6aPsWuINDN2FJEMMTEFjGHgK5/19dwrPUH15rzNNjwKUYnQvRrTdkCGUL8BIHoF
tlCqNS/rZiAXsV7nCfhsMA1MTTZD74mwrDNq35xgSfsUn4V0bZsxWSOGD7jObZ3P
jxDvuQEtPLl1x7YnoMC+6X9RyDAZmWIJRu9Rc5+81DEp0aHd1Oknqb82vdo+kcHK
dFj3BNOZy4lgNr+Nt5ejV4S62m/RkKbafFFU7/NuSww55Topr73tYhtHS1J3lmGD
UZwO7NO3TTsyUKVUtItkm7da4QzN6QuPe5jcgRH4LnQw6SirpU/gFENpn18CEjG2
YhcwPXMIpUKyjHQInmta/koe51EKC7XNBd0alJlLrkoiE3e4CXay2BB4NJ5DBIUh
3SQx8PdGpcMS4oYyDIM2HvQqR4moM1K4FqNZwrX2G+lmV9cDzLbxYDBGKCtSm8WU
BaUy7WZVZbMntOkAnox4EDvq7+cJvmZPNYHRjVZ3NiCi/msDqqEnlxdyEY9Nyvc6
bb81RGkf45TOr7QV0kvOxm+x/hIrcpwGp3xtO8DvSPHJvhEvJOpCUveDnvDXOaX8
KPK5RTFSPg9sS5h2dV4vRk31RyDTovmi9mqv6eVZvbzFKSTwJi79X1bcXtm8PLZW
Z9MekSUnL54mAU/M52MvAf5hJK4LNQN5+bG0zKHXAh1xdVtQ9+eIS3A9zI6s8lJi
EFEG31N5CePGw2Cy2xKmnYv/eoanUw3qJ5SLqkvn03gmBstzs8KMywb/1zIByWcS
ljdf/INRfbS02ZuFTrkxgUJ1MTgbbJyWneXMuwHQHhD+IQ96xkY/JM0g62lBO/SW
pSXOY9q+3+jQhuIQsKItZswfAspfgfAaMzJT+62mUfwhvxwhPSS99iZ7A48foDf+
+F7+7b7J7dkD5Y/zI1D0cFyQAf/gRSq4yHV8Yp4+PRPEFSPSwnSPQBm0LmuOXX7X
qSWEjfbqiLJgU+jns/ffAjYeQqbftORzdm02QdUuON5p3LHvSSVu7e/LWlOuVo71
IJx/gWNV3zTi7DiWSm6gDXj7hNYx1H3N9OHlzJEfGAHoVAm2iYASpaHmawxbuktG
1H2ZgAtr/Q6yfS9g2XRfUdBuXRK9kGCSSK69I3dAd2xVwWnouHwpXtq86wDN3V88
Pttohvq+hqh4G6+EqF3qza/fwj5ZqUM1e7vdyIpNzDoDGVRZTpr/jg27Z/DcP9zo
ZR3XGC+mbWxnGTuKIHXiQeiWlGiXPrlDFirEwKJyB4+zkxelLNYbpEIvv3JX8Gqm
3jb/eMX82wCzmHvz3pql+hOGKpMm6G53TLaayULduHTpEhXkyYV0RuUcJcObErPO
3A/auDO52m7hFZlMgWkXLFGqnq/+2K9x/dFdQpzBWI85ierPmfxw1/PyWokL/Sor
nZWD8m+e2g5ADsiDTNm7qVf72IKcROArND3BV3MYM78LxqqDoZq+0aEZ11oO4qxH
w1nbFe3vsWu72oWAaJu59KDaWXrUM/HYU752hYv3Jt2OY2Hj2sCq3qiE40EZM4vh
xAP3A694zOwzdG/psXjqxgQ7uk7RHZxCA29rJzkKOocymvFH2e/MNaNGbvuaaVOV
LLVT3KUnFVLYnYbk8iYFt0HUAlzOA3Ioum7ACpTCWxq+JR8tU/jF0yqTvMUTafKA
U2IB7vQgS57xgJ0VJ+Rl35sAFFY/SVqJG4RFaQkQM5Cd0SokE1j7fmHbdJ0tiSJB
LUOBksBjVdYICrmMdmiOxMQE+5EqqgIGM2oC1svHeIMg1gQRoGdWteyN89nrUmQj
kAc94d4wbBHDmjUCdjEApseJ4hfOhaG5wSjGIx+355e4j0cuHLOn1IlDjkB3Vq35
lDt1qPi9VUBnPiXT82TzjgdU1hJamRFo9K2r0hbdFRrI5f/6Ep4YWG9fNE4ujDgu
naYduimj8aoJQOnaIj29mN0jRxjRfPF8dBeHrlTp3lM1/h9yHK/R1nRf/AKlT3wm
ZriUT5coDu21lQo8NesHHp26U13t3P7Wp4x7ImyFbMhIgjLkgz+HoSs4TE7I2U/i
dn7TrxPnxzOMW/P02kYQDGhXQ7sfvawDtPkhIPG0YGHcta0/7DLgqOf0CjTaHML3
AdSSot5xkomZAohBQUjwBY4VrHEJYCx9I55Wfu043JyLp8DZ05df0T3q1Pgi8CYn
FFSb36AICnsE4A/qb4FXio804y5GCXsqqjW//IWb9/wr8KcPVMf4DdkkUzlVdF64
3uiwHeM9SOMx3Dq/2OsUfhh8qhnbTYUCwKkk7Y+EBull655V/IRjfjHILpyv/2tM
dAFnPvk7/Aw/wrk3VYYNdzhDdpRf2qyhKtpbxsjFLE8hWOdZm5iZsSj5ZQOIN/Ne
F2q+OUyD2omCscwSze21JKATu45/aB16DNS210WfFm+gR/AO84rOD/vIloJFTy2w
udKEB25lWDClD0gKT0VkmBzj52v/IrsXFwROgHvDSEZzzkBeWFlKTwvdySWBkm8r
FgLViMfnXcVXuv8fIuyCnUGU00TqNhwPEFHaoCILQjir0UnACupwDhbQmfsPjSPA
TlB/tjqiEOJyIqbl6GVLbrzdHfKdCG8MmvYauExR1Mhsb3LD8/aj5vEdwUWDvSpd
zMYxKABx0DhAd10s3eTPIAAP8yF37LjGb/w2TWw0p1AU+Ubnt7egZnZqHs5w2XYc
mwgTKgKP5YQd0FMqfgw23xjrVARO2twpwIOzwMncv3bNeaP3SbAZStXdGOyU8E3l
Z0gGnUROjEM9v1vjNQJ1wCLc8UFecBA+GJbMdBA5weY8Tbw/QcWpQOES7n8s/pHM
yOoVtSkGtMVeysvtN/0+enPEK1OwKVKcPZ3KkXQlrF25J4hIGmxlam59r4h5JPIA
2DrNV3KxrSQ+Vnxv3MNdD5AjULCumnWC3Em2A+ASdfMUe0qN07gErzuqvxiKzwlU
DuDV5/gV37QPg8nMhhTtRI/wmHDRE+6Kc2vfC3xaZMBZymQKWGC2Qw4Omk+l1WXl
2UjvAjVN7op0GYR1SVfTw4eTJp68UKhfdplatoHv08dmoci+JkNERUcM+gFhdvqn
qJoJ/wDKwOdYqilKHLWnL8qgLb+KG15qAImCHAYsSAcmiPyAfnByb9qj8XU7FV8M
1AiXtYCfvSUyOUTsHmnprP1pMl6atQBe6YyAa6v26woUl9x40QTobqyg/vQJJNrb
QsseC/B51KhXb+ZA/8eunV0esGFwPk0yXnzpZvNV+sIgkcYWaXy6dTLaOL7ZiCXl
ccy4vIajnqZ9zYNP1C30Q4yHWsIJJa2hDLKKbitsM5EjSw2Teu7aGWpQ9B2VL35O
kLc+IevnvL0/1JdmRuex+OwKeq8w8LqaMHjOpK4mFFYhJJjiOl/c3xmaKdvTPx5W
vOnABkDrPMZW61WZDmkyuQ17RWkqN/rEkEe6vIrhTSNJJWIYQxQaLTAzUYxuqiyI
mNIgBvk/CXT8DTjxAb87mByMYh9CcHYhPo+o1j0642KxwlN+JHyZMNHczyVYfDTq
FztnzW4a0QSetgLhk/4Xd3KEuGHkB+JeGT+W6urDeE+aGflz9fMKO/XxvrB+92oo
JbjD2RRH24v30eGU9i3PjqmiRsGQbhc6Gv/dIpN1byzV6ONJ1YYrBtZ+ZI17AoK0
Ho2yFlbs9UfN2uec6bxDDNTThJnKex/fPwSbTePBWeIb/uA1917uAKW11xgteUgN
T7XY7biYXLOugOcki0a2o7f4qCLU950/ki/fIxDVB8raIHdqFAJn+7pyFSBnM6qt
VMEd4u+jh6Vok9thQ2AXU3F3aE951vnZSaYOW7OimqjYCIgIOP4pyn2gNybQs51a
yJDba5j4J0DN1AXZqwx/Pqug3zHFNYiTtf6qsHrUvRGXalULGxtsOIY0ASZbOFsI
5rqhrzEmjhgLG7dBVX+fXRGlpJga5SeJCUlrcUHEpCu0Ddowu/IUV5Sdibb9xLpV
taEvqohi+MbzeBn0zmUrUrBv/mmRT1KWQmt3xwkfMbTpfOeFyjiMSbqDYkGmkGAE
gXygb8mm2FT7ud9WHk4Hd/B0rvYCUBtU67wSydtSCG6TXxihX/WrHYSHl7Ly/vAG
tXYQI/qxI7w9eFMHtR5bcoajHa4ymlD7SEmyToqfqyT9KMhSf7MOlWsOJK43Fd4X
iB1Xvf42Kws/3UO1XFb7RCGLcgQAFfypfwM9cnzmZuWZq8mZo3XDk4jAxw4CMN3n
Feq8ZejUU2Bj2FDdiM32PuCifbL/djv+mST4DXOf4JZINCzup0e0b+gvdZY0gf/n
B0B1D6xXKMjfV7A5iugm5oPwVOn1o3ffJfFljgaqf7qhflzdUQ4TNP+2lD/50R4y
ebEcz7QZPD/Cq0V4Dzvrk3yzrc3Y9jiN+fsxR1DfElvchhGK8YjmeHeAG4uzOtGt
ToMJkI23knfLR7QX0LBdfvzpwVRvzjmkaVpsoSORcOWKsteRsSTlA/TJADOaYvw+
sDCgo8KtdPK5IAxBFuugAE6LyMlC2zZg490E3sujLWCKSDyqF8Iz9llVvdN93sIZ
q9GsXFIDXklIj74shZfUmbF6NGTmIpGMWjnOqWTHU/BxuN7tBw8prepYk9v1uDy+
nMDpt1hPkNTGdEwKmNXeGUFHKOBdXHj4VdIlSB4poOKFe7XB1VTCTyy5JEPhfg+3
rP0g00F8D12sgtNT5UkBZnvum0YDcD4qKHZLhZ5LfMcZtNzp29XTlnTqVoJtvx24
yf6ICa+hjSnFa+NLxOzVxdXae07KghNMM5gbEzXVL+NIrh/lSvKXrqvK4pNWYg2Y
s/MiYbsCMZesJ+9XqEqqH5sEu1tSgrZ+1UZx9Y5rv8V+QRt8nLfjsxuE1P6wstHs
zQbaI/daIQpDGhQ0m/OO2VhJQvoMhXsugXsDAexJbIrkitcg3/XI6StfVSHG9acz
Wri4+5rwyHJ9mbGgHet7kfY3fYBhmKSAQ5dM+o7PEtM2SM2qIBxYhtBpFwvJ5F/p
/INgSg/RTPH0vsmD/vgcAFUsU3cKtgL5TDEWT/OSpErUxzwKUriVhgFaXxHAIzXN
T3JobloJ2/DbqKmDVMz+R1jfs0hr3TzpJVWwNYx6blY3xEwtDiY+BuzvaJDjhdV+
mi1+xzsa28yTQ/GQfxP33nly0j8IJoXG4ZWYVkpNY5NE+1JUZ8Tm2N2T4/+hdNZC
LT8o0ja5cMkJ6r9rXaWVHnBsQCju8V6kw6ldOuT+Q5OJRnlsOctOxBqrKBRrtQ3Y
Pn+BJlnluq0tmMD98vXe+0v0J0K3darzE0cMb4rL5bLrXG56zIl8dMn336gfi9XX
wDsXEdUQvGZf//tYuMSYHdIn1T9zcpmTKKINg4tJedHtDzz2ueczzVZDKrf9MAeA
+ROIxTjq9JqqsCCT4FPPAGzA5fC2KzuZBnsBr2T4ub5k4f7Vpf65vIw4hyiI0Icd
V7VKPkmRoex8l8P4+VJgDmSyrdqQ/NCogriuC/geNgRmDvT8PaXtycKLYxR73NVB
ktgo9Fm7Fu68OHKyOsftGMh22RmR29lAe3zkkiOqLNmK50MNKNoc8fpL9KX9s5bw
wn8mtK9skaXlZy44dWnByWCOvgw6r1Ealfo8qUiaxJewoeN0PumVEtgoxQll3NFY
YCEI0h3rcAMg2osR8yWpmwLGgnhebNW0t+7ViZ1jb8UmLLzW3SdD6xzg3T7E37Jk
tAw+NHZDnTXu8EEQq5xWxOsPpBL5Y93NSnNMcTP8WHwHOnS/zKkCNL+t0PfalRVm
bFBJ3ey35YreA8YmQgSsruAtzMQRT2NC1bkF+pnQG2kdX81CcvRm5yvNiv/LXtRV
XiK9+k1CkRnj1FwmUXBKrMlwKut3+JjFeXm/6y5iKdHPAANRbbTgI8kmHmpbS1vn
6GZgWr4zjlVt37eJFn8HJuOqOmGHwpoyqY4vP2+VF49KYgx42bCN/2eBNUaTpkgk
PUsEbSyY20XufMyPv1to+DIDAZq3S70/u3+kWaMh3nAwsLAb0DECQaGLI4q9OsE4
BxalLqFhXCaY+D99v9fwIQ4prnpwQl6xQp0LZdp0kQdfQ4YeDHqq3U038lNfkSFs
r3Ckf2ISO8F2pBxNCMr7p+eCQEbmIoXV0L1c+juz5ah3L53oib670KYjLywXUwb0
FuPOeu7oLckvcRn1/+yH/p2TwzzbCmE4woGPBbe3NF2TVqX+ezFFo/n73Mf/hD47
mSRgom/sPcu9l1nAoy3P2rMYtJAkrx9tdFgvJilPAkhvss6fhVSE5ugUM6D422cx
I34uK+19x9GCqQRDqsUJvi4ur1txzQmhb93cLZ4NaPm5oA7wl/SCBDeE4z3VE9Di
MRK5LL2yvSVNXM0PdKrwi3IUUlep1ZoJ6n5wZyN42hhYUdN565HKiz51Vog3Y/jc
KOTAKwDXnaFlP99NQUEYLSgnXuse1ZmgmUmEB2e7WY8ajUkkPiAnyFI9YFItJZTD
sXVYVZbI1QzWvSFPRI4UT+Hw7MPoOy/1URDPqtEclsVB7Ask14AKAfkGZ9NJSZ6R
jZOJ5qWltC9f8ks0uB+x6vNmIXhkCnZItR27PEUlOAO/f7jo64dsnYyTTfMXWefS
nDKadVd9qNt4AKhzFOyHaUrsg5E2Q2M3CGVmewY7C+jSw7dwI3YjXnTtFz/uo5va
6+JLI4fj2nLanV8e2rW6Tft7e2rmKFdaJIDV7g33bvE6KS3NtDWsGv9A8jbWjPKO
4S0vrI+fgydDdTIplNqG013bIwH6vIgRUtkvFgr2rAiQDfKvGltOoAL5m9gbl1Us
DULkfBUP2DCDNk0PtttK8bSUVr8NnSRHQIBBgIPvvyCWnfmfgrxSnGpnyr+6nneF
vMHi0DeHDC2L3VUWe476/m26b8YX7q+Amah2UN3HinRMkI4fN1nW+QqDbEhyKWoV
Vd0m6A22uizIl87DwMxngTLDxJUHFqr2kPxU0TdS/MN1ySYPJxcBvh2OjjzytZbD
yNfuz1NGO66ptYF9cs6DTqiBtWtme9xQg1vmB7A9dOw4lwf7W8h7P5G8PEzVauaS
kTScXelwv5tYTrwgwVkbGSYAnuIExqo+Ayh19TYFAc9kvSLDWeC1h1hBCtf3h4QI
hjLMqA6Yz4HqNOjCYy5JD/29IL19T/hUz46VECJQClMXl0IUPW/oeV+7AQ6WAlmX
kkt59Cq66fnNtfmE6NqGJydRfPfc/7rTqgYfDvZmBWxCoQW+7Xncc5flk5FJe14s
SmzOL5gkhuZ3Z9uZNQNdvRlxh0X0MHvo7UlkblByvJZ+BVTmPKNKs4/5ju/cKhVk
EiZ7W17CT+Ua6PPXOihnV+AZNhIATlerAYTV1p3t0Y7+i2Wdt9qlTRmtiPflWeap
7ZyvT7DO5UJ7jxIeLr2UYufLkF6PtLWaxX3gsnsnLquyONlfe1NkRkxQvRcL5gCC
hwktgYEPRdBUyCnVFLhJ1bzJzaofYopNDMxq/TCXrUHaImQEur9M8C22Vf/Y8ILs
LLIXCl2mSm2or8n7I1O6wl2Y0dtuszZ5PXsHNG+s0aKxxsR3vR+Erk2dYXXrODyJ
BWBBcKizJndY9yorYcgbTpIfoVYiP50V86m5dUHOouqRgNQby3i+4ttIdAb51QlO
xjRT6Yq7mcaGuS752HLTHgwyCWBAc9vo9BjqXPumx6aV71Wj9zfY5mPgwvWTSboQ
d199o5w3Gn84RTn9RFOi0IHv9QzOZ4Tpx6AWPZ21YaNRH3UmSCJAxCFTqQkMh1jx
9UklFBZ2xHU3x2XdsIP3ikqiqCUCsTJaGq0hXExbW4kGSKfaJdzvkW+U120d0ljF
zR9/MdEXa7lNNABOZC4iU0ToMsZCJc8O+jhSRALxZnzprosjdyTKgIyuLQEZtJza
hBzShF+9c9VuVNiwKr2qIDsIDhxJxUrL75WVA4XdnmdZwEVYC5YYlePXp1x+rusV
suRFQLGvk2ziLW1gllFSTOyih8gvPQ60RkhV8/vBhJgQ7hof8obTIvEMPjtyGfIQ
OFP9TQui3Ub0EFSitCWKsWU37p1NavhW/FujD0U0PRfDlc9YFtwafag/lHlYbUja
Js7e6RNiRncDVQTIrkftVd8+KEzOrHxaepZ2SLTUH2XJTQ7uhTZOZDAnSIZhLbfJ
dtgTKOVrWs7iDCNR534FQXZiJ+anZhmkKte950Tb44AC61OpGhUhTjiFKohzZDRJ
IJuSfNBqm6p3K+qgy18lfusr4hVtbulf5U0dc4/f5pkSHZmrrv9O7oa5pdeMy6yx
zq6LnhlUjwV3e76GQW3rmHgpNKEL0GUYl+TdEPzMW2dEpVA46fm8OGpll1ASYCHs
cnnhCg67d0KQN93GZpZc/FmIpb5UkaP5G/Qte2PqOKO/WivQahurS8rnmkDCXEjk
sc1uFL1bRkdEfAGQPXUl5p78tnZuXZty4CYoYjXspvgowAwKKE+eThDsT0Ga4k82
TecDVt0x6F2PPU3RJpC2sXr6TKxeRvRGoj/69Mp9N6/ixneAIa4FcfvdUmsbWlmV
ixhReLK5L25+O+SACLKQ+q0pABhwWNlb2HLrr+RutDQQFfTqwraRfi/DYNkr42iT
y+BFOOI1XNlKn54eTBxvMeJ6Kc2ooUyb3JXciZLhY9nbUXotlJErYh9xypa5XBXj
hK5wNpWPmIsHE5IW1vPCPMPMxu2JjLEHF1M+CCowHwNh+8rc2UW3mhQTbl0RibSx
lcux052hU65DmFyK+sEWjHlGze5J3FQD/SFoaiw/nogfXWlWzTvj9BlTLZcYJ5pM
SjnhIofbOLnpKJBc1bfGT+Bcvr6LfKB4WNGGuY5bfzuBuQ1+1RXZXf+v1pOEdJhx
0F42KGTA1jdGiI3FhwuhOOO/+u4ZG6Yf9CgCpSTuS5fcnriA1pFuoUbA13yCatzv
VtgICDVnuwismVaU6aj2QrfEo4fXWISXRJwmXzvnaFS6i2aJqizhwrqEx4wvCRqF
PbxSoJnCPwKFgu3MufTnOYtJ6DNaWBTNfHzdImp9NkVpf9o9e+AwizWqouDqsX9W
MvkMtxuTw9FnQnjx/is4vB7ujgDCY3uq31XVH/yY958eIGLplCXxg015JREVmGFR
PT2adU/hjR3TVjf62LaAuDcp1GlsawCUL/gd6A/+v/hbQKMyQFNoQR1r6/UXKjBm
JXpqM2j++lmtnBVfOwyhsAQeI/FxcJ3PECfBH/3SL1RyRz0mXf4yXCKribtuNy6K
szIybIuWJC4lz+y890YNO+v0CAcJwr5zBfv8meUHE2v2BNAXygloUlEBwkR14P03
dlxcqKJPbUZ8ufJ0ylbDYQE0+Iz9qPD6UB2OdPwMzJc7y1EFsTHPEy7A8jYpbViv
VF/A9TsHV/y69Ql99yPLTBmYospD6HxLQVSlUxObqSTrpnBtOMYRUvVobDfxccgg
NWFXthJfWokFOXtVvRttuLk19PWOu7KudiEnyYqFHSl/UkSq8/AASU5H71iFWdcN
a4s55+w+eMwU+J4rnCuPcTkZSRL9z0Kh39hDyaJYIW08vhxTSuOyhz0a8BO3ty7C
G9azYLPqUiRAYq+TckJZHjnCpncI9ts1aKa28uZbk4H5xyrUFXH8U+mgCLUpYdnY
oOVTwKEDvFr7SYIN3LECx+HBfEKaGlr3C4nA++qGJX1DtKBxRg1zgbRQPbU6k4Q9
txgVaP5KJ+X6YpqwsEc/LN9jFJ9AXQn7KZJAj5SB/rQ95nzbSmxmpUipBOOL4n3R
4vrSc78lpjysYeUVYyt21k4f+JK/zRGz6CEHYaxOj0iTTU4IN1yuxOk0m0v3QVEl
vk4VXNh4+cl59BZTVjyoc51UmLz14v35JOjmgeHNIB/T80s1sw0SpHsxUK6Jyexd
kbPpazDQj7NBtAl4/H1XaE5J9jU8yH7jwkTsCJ8bxcLB8thaPsGSulvedtfxbQpq
G8iQr4YvjE6ZDP/66LG87a+imb2qZlJO7Vf5ocF2Ao3Dm2HIB1qcp0DlnF0xTkhv
SUmdZthcOwSz7ia3FhvvEkOExE97VyJ4aBvPkxAsK5FCLxE0dJ61d/lUnxvVTeV0
alj7K4A8/o6ehJiwWZfRnlf+GR/KyECh9nA8BSNs3xT6M5akh5A+gpXG6oXjw2PW
N1HUkEZv0E2HMWeJUjq/a7j4DE6lSiI0sxSm6+2sdsMiOPN66JRRuKYabgjQGq9j
ENbUZNlDJT8H8iPiF4NR+Jra6QDfFWuFH3Z0orIjq+uUOS6Cwlp86pzG6jvbh9rW
RlKkZUzflgWU3Uj9CHGk4RR98ffwfgLNAUyyBRlyyuZlZeUNJkKfyvgN5tNdEaAr
RmktBdmz1MIUCLAjQdmc1bFRtPi0YZWSFATQ9vicLommOudSGZ/0dDFYdB5HKa5x
ry63gn2Y82JhD/ti/Ksuj/Ib2CClVQZlUEN6tKni8OFKI2TlSq1iCVeWXPewsUKP
jW4XOusozdCTIiWMs3YvMG4BhtD7fyu76ysYSqwkVerqvNEuicWPeMMqHVtdMnxM
e+HHTTcarpsVCZP3jCyCAkKBLY+muupgXE4IZuDZLdxFCgL7Nn/sSD4gvtMqlROJ
+oKL4T6ADqdcURbXBZizMg/hLmq4KYRlL+LpN8+kJ9LIGfC8iOohnAdAcN0ag8c/
yTYrK4QorHXZdJd/723nmh5qdILU0tAekjMos4Ai3tGaiXqPUOsBarqUwYkpWKB0
B/oknQmjczmp2CUwmlSY+ReudmIXhQkG//9JclGm5Q5AWjALNQawGpVavA2fEgxH
j7reCJWA5kCB+0GPCv/447O+1vh4WcoEOgG9u+vJQPOEEQGY6Tq6aea0RIAokauo
lbP893WvcKJiU01bxVefhGEAtYz+z7fMHW8XjihVKCGbjSdXQa+dejTcOz0CGn24
HLZWCC58scEfK04/HcZxdBfgMkSD7gukbZ4LQ653EUUWrP6kCW9HfedlPOz7Mi0M
JQIzNIt54gEOmW4lpHdD8dUZXEko4nbhqNhXvtXDvOQOEMVrQ/ougjCIQZB2gzw4
8ki3JDDPnmVZ+9p8O2IQFi0gkzAvrUty//uHeWoNkZwqHSsM25GSWbFF0b0JqNhk
hyj5o7gnYIs0ty9mWYAalLL59SUeJobGGlJxtBPQdmxgyt9MNKXigUXG5e7zv0+d
cnPAXpSt7xsNug5ZgfN+K0RdAbALS/xOvgufsDjpQuH9A6WO0/6rMvieHMCFPyPp
XhbbFeUgn9ZH9lFpEFSCPDsZY8SdjITXYG9oZ9c1KX1GMxDOx+zvVVZqTn/gtLbn
D6wfFVzy8O5GGxaehvJJgiEQ7plhpMSxwKYhK20+Blepfcs5ojjRNYT4efItZJa4
6+Hd3HyAh6zVPUWtgdOcY6R/yUpTG4qChUWsO9BJxPsV0JTiRtz17rjIQctolqbI
uPozDwSTTOMDwySAdEnJB4f+CiarsrEh5l1tacy+LUMg0z9zWdY+1X0nbG/e3pQN
T5FSs2hZxuCZpT1j7pdEHxggtmthjDZ4XPd/16Cd/2KQrtgXXAMib5zZi/Px1f06
lD2HV/rHy9x4Pw8byiFbdJLqlNtHzUVpwT71dYRJAgsmn+ASNb3a3RmJYjsSHxAt
lE/bHLBsl+O8+jF7FtmDiJr/KUH5wZ0dCfuwrox6BvBQ0i3dT2iXS65s3j2U4xDa
vbVQolnJX8BKsS0imSPpp1dquVy+BEqnWaGIrHEraIr2ZD1CKz9QjzTj48jpH+G2
2lR6kt7ne/cOd08r1blG1+tZ3OXde/CRHlKXNxWWHR4BtpvmyyTPhQKw6DGhE/b8
ECLUWuL8qfcfBeXWcEYhUaVFHteSF07cw38uhCmt2WHD+ZemMg0+8ntjMmYQp47I
RtEvoQ3EixlGcIWS86PnYCymwrJDRf5O2ZUeQ9BAjyaitPXcsE7wCZNzArExsRR8
20PLCkkaovGXJMF0M8qpovH/pV3V4rtpiKXbU/AwchwzUGfxvsS8x2LZYiwEJ3wa
9fyO3Y9k0NvK/vlJm0yfJk9lmQmzfB40sfHRUaLoDRjJo6467QvhgI6mLXmkCvBv
Y+VYalNpa1F6mOeOHa551kQyhewHUs69Uf3vcU4yNrfVdon45iRCs+oE5uEE/6D/
O84077odT5CPGvPBXBGgpbyTnackVYnsvZkWNZy8umkS/PCvgd1ySR1o5HvjEIv3
VLWAk/YVA1YyQSqmeMvkf9P8Xxv1R4hx4b/UDwOY66XtLgvSYEv/mXY8RR13pgCK
L7AsdLr0kf4iiTaB/MvFMvTFak644rkWN5uig2icJ+BLTob1nliYjdWNTodnf/5a
uA1aiTgx3WZUv42SbCBpThiH/esJ3rg/sx9HBEVkQsLgYoKm/ue3FJ+23I8eFP6p
4YfKb55mB7wRnZLLPwJ+EWX63xHndjj49xSlMISuFexZFkKrLTIsO7dv6cejfWif
TBdcDGWxfZsOi6hwacY1DXXozh34u/YDIeghwwtfC65KniliLGxCHvHj86lv1zr6
Avuyp0Kmuqu7c/3Xz1G97wIgzdBBGgJ2Yi1a8dg+/bRbrsK0viUwQe1Z4S5SdlMQ
qM5d9Irrc1sf0ez1Oq16fS+7S65ZDAcvH4KFYjvOZA8lhec8fMPPzpFS5jWqj5L6
5pYSNfqMmNpVomOx1qE5G3r6XxSttkuM9OFk7q8273fpsdfhJBjcX/pzeOvX8AhU
C6rQBAqOCj4jl0bvRaMaYI4yujY16r4WsmskDORfmJvK+/q85gcz8vrCGjmN6JL7
vcwwcWZXnwui5SEgCCIj5bqDpp+9M2B1bDuFlngl223qNScqQT+GNai0m627nQIn
Gr9/OjgWXCl8wdb+YVGH5jCj5VMyEQI7lLmSjyfdin45nAtYRdqrvQL9+QyPycJm
a2LISHKvoLC8xzFSBSLyAf+w3j3FUuPxijkN5x/P+O26bQzCh/qCE6faxN5RqaYm
6i+AHD8UMqllUsBPtBbCxIdwUqCtE0jTPrxwqlZzVBZFXqTtC3qltavWn8/HYpuL
Qg6mHwjvsijwDmpNSygaju7Bj9mChHbxhsBCuqnMcxmcdPMvSsoKi3/SGKbXkiXR
tUc+aKRBfoB0xEgROUbIChNELHkeB5BQOZJaV58Ds/pxgt+HUk/6EvsH9vwLyxFD
BcIpFGZdoBvvy7OYTmwqcL4FU9ncqy05sn3hGHgjHTW5uf7IuXSg6e4qmyEXSDNI
x/KY6ELu2v/4qmS2f2e+UDc078ulDEdLZ668A6DqaUPgf0pehWXE6mUXPhqEsGoL
EUz0+n7nqKTRzIPZa8jDkgz3kzxZMmExc76ftNZNiCR1ZtgKsVIH/cjHI0UpfOvm
uE5UI2IUadbMkL/I4ILelOcqmRtHFiRcz8o9n5rle/RRSYUeCx1tHdTgqdU4Bjzu
RmM+mx6AGExgC7YJHgx5b8845dZJpFypzsXJA+aJpQiGO+uAHhcKwERBszWTIWwE
khsRQStlOV/LAKTP6gSxfrRERWpFqMMk0BK9xzuy0kgSR7q6g9gJUMQesE0G8jOw
WXvvV2NCkx4uVxDHvLpMpOsPXr/TvU+6ooXRXg9lqNNOygMBqPUY2bkx1cNCTvv1
ZF8mGHnBYiQ9yOLKMLXJKB8PDyomVR8IbqQJNgj75CDpEfptf4auxucP2j8Vt/EN
qCMsb/ieOi+te4CDcyURDUJ8/am5zVJfFQJLRAjdHww6uhZuJ9zYrzQbHjN+c2Rn
s8sVD8DrjsqupFzwlFrH9jNBPiK22k91xyyR9zfA1W0Ajpp6OZr3lD50YILgpzfH
32ClmqfJchAetYk0WzYKUAPERDo5NXqdXRcvFQUPcN6/3BuAhqKDhFQc7+ZdTqzz
TezVBwj34UneF7qnYqT4dZcsJQaEJZkiXNdrMMCZ/EBbZaXmlmL9X/G7wCMLlGZT
ORTCUeRmkRXDXFcGaK7WobDjMejXGMahpJf+Qwuzicp2BE35ZBUku/1+oqYAVA8x
ZJVqXS9gJIlzLDVG/96RpTD9yxINF6eRVroaZJrfGz94lxX88OmroOWGnaX2xkVd
u3vn8X82cbrGXZM0chV92XpbaaH32IjZBX5vfgYErNT8edJR3pKy7KPoRlo9rqts
V+mS4G0LAPA8mhu5D8x0JoyFllu0WAXoC6sJ0E3uHD8FPPraM2J6V5l9/UKs7OV1
eY+fJMuBCNKqArL8TER9ucnwIarvFZeOb3LkqoCJnRJu8ssGXR96QgMMKrBQzPl9
6XjwvHu5MQ2unrYc64N+FRAdIGhG7hh+DrBLwwGaboe41x3+6Wbw/ydlAAXYdehZ
mP5uG62sO4vLLP5pygn+19jfoY8OZA8qhrCbLwiEpVXqsdfTPeyOuirqhtctJDC6
4eMwLdXq9kDOpbN6ksMdn3gTIeoES9chI/L/6czBfOF2buSBDhwne/vW0ofp2Zgp
+q4I9bHiwI7qkrC0HVDrOFBTU5QECVeLUlDSujeqzny6hWOQfyh+5BwhYx4+t8si
Gr79Xud53beGj/VJLtOuiUHUnZe/ltxkJd/tQlwuCWpBBFemkAbPRIpq+06AbIyv
/V/2GoLbQMfTrGsCwGY5CF2U3XFfIbRQsnGJBoKaT0OYS0nvpg21pG2lbH8a60Jb
Y42+L5Dr7fYVQ63wGOomIrYs8Lo6sHdjMNYcixa5hQ5HBtXkFfV8cVbbhsSCcCY9
rTBQzyg4zR1iCSAXOT4pGKzkjM9q2j9lhvivSvn3bmufkCfBBYRWf+NzQRH4Rd0V
g6jpD6qpFGDKjNhD1ZRStQKtErY3/7d/S1Z0wYYrYjFiEa4FI3BNuDFgN4U1GuyL
jm/ugtiZkGohbJps/vlCaz7Kd4n+j37RxD5vESGK8lxuQDo4ZKt/sjRKPZ4pcEEt
V0BWRhWjmWi/8tRUt2RYGAUjuCvFJaBYT7wylyTulayr8diPGBVj1RC8GZ9w2Uxw
yYVsVbgUQlKdR8pmy9O+dbdKpixyUIzL232w66mJSHoQvEmiNPQkDc0s8wYW9wgw
J8h8CQ6qDAOMhjtB+zl7UMu9i2RmM9pBG6qRvCQ3mEyfcvI3hvgNgJqVf+92N2VV
M8Kha20GijnVm1O4FwwBhCJOcaNSCHLxgD3u33EBJClGgK04K0CWkkhpxsx4ttp9
bWSotz9zpFezMcFSfZKUeGHytDOsRR3vTYkdCb31/En+oes2GvibABjpl90RDzAv
9Orjg7doyqcFg8chI1drS/l2B8HtnIgSq8TpkqHEZx58Sde4fmYeuvTmXOrL2cXX
tc2sfn5K2VEVIUgdQuvX/iLCzsUdfKjyjmTQR0T+YT1Rvh4a2RZMJ59xmJhV2xC0
8LXza4uSGedJbKJ9f+XR/vWItB5drOvp/CSnETqJlQexIVCAS4+pAnXJWlrwiXh7
LCol1z93kS5F0HHZCeWU2PtbiW4mSrX0wmIAEFNokD1Qi5DoQ9/b1E+HSz0h/3Q6
sJ8DRHrORc0Bg9sBTBslCucxY7xnp/K1WfXZI/lnJG8kyRaAZqihZXWz0Nzk0HlW
jxrSDecWnzaTtzOCZWcZxn5Jos6tOiAwL8Zq/6W6VJXy/dilVLMEy0K0xvjMgCPD
2/lJ4lq+HCIdSlT0moz89Sr1rFRYHl9XYzD8zTzSdJB0rxR53Ccj0rluvUS99anq
/8s91hoLOHLnmiqCAe25gA31vN8W8MLKq/T1oKcxeprc5vTBHxSokxGAED4VMoUh
zUMfTRCje+MQ2DdKYQiRPaa6uAv1tYK1c+35DpDX11KqAREUN+GwH6zuTwiadirb
K8Bf61dHKP4zRAvKyGdMTdjz7HfpvKCIFI3X2mNVOt0H8tsCjFruC/niw17u9wtE
nZuC4M4ZRn8PhFtcfS7zaHIlqLDWxNsNYMVd95D6qhnUhDbQSUA7X+toO1tGM9v3
Bk3Sf7pkISF6T2lHTA2jPEp3oIZ87YBBahafPdQWv7sH70dG5+Um+AD9RQ5QfyzZ
X/AyFVgHjOunaNO6rfyoLmB6In4JLfHngN7LcKwVWjHq0nFiHT8SGdHZrK9LFlRm
pgt2csXq9Wp5OPaKI9wLTu/FaHiEwZ2uUkfVN8EXalL0UOBym6OX1cTIi5fqG1w2
EC1gIIa1rTD8rlnTtv0ecw/9kGZ6reaRuVf6t5LtGMSwHMnPd13cW2JPPZ+WeVlW
jyKLcK0IFD6bfUWqtNyU2WgfopT6x2nl6Wk07OuaOqnrp7alI2/NPSTxLk8k7KbD
Jl550Gc2WriG4+pVxZqZDK/sQF3Q2BFQik0WWABG1rlIn44Ugc8m2wGGM1GdhHtk
vMW85uRaV3qTOSCIS4fT0NeRLHLzWhKNxSOtyTb1fg1+kK+3E6Fn/6HBQmU9xCAv
u/VFVjgJp/TiHnpdtOqUUrOUjGRhpJ+Frw6v26S2rb8MHPB87rfOnPzN5qvRrkdD
8tuOt/tBQgqG7gIG53DlrN1OBYhcHPUieLQQOLJY+r6dCvoP9+h43fzP1ZBDj79D
iVnAQ5H54CsDRInEWYBUPseg2dUtqP4PsMsYJHjrFAX8KVf1fN6wz752uE4dpV70
XeKZHSU7MXic73XjPx6gfd7glmH+iJzDk3nzGrHIuS52TTsPaon8ogPH0YH/adVW
YHO7obeIYBBXZmAUW8DmqK9ok5CmuWQ5U7N7Tg5dhbkoVTiYr/aMUA/+Ipc+BFDp
VtNvVxy5U8kZpjQbMF659aLGNvuyVlxjvchoFnXR6opwcFehr/6EmPG9R57/OU2M
TiwR9D0fn4qyK0nxpT4Ql62b7rYLOwPcYTk+EoPjPjbF/ZP7gRmwI0LmyShPG9Jk
c9YGN0x1t2C1COWtYo5P1YWKwaQE4wMndcpmQYnIdAhI4QXWhYzrOXyKx7VCmMbE
tsZoW2x3l+a97AGDVAoso5sdPMVYZDBUGCfQGdd7uAnFwkqmn+36nAI7VSWSlxKN
fIQg3bvIUN/bQ+mQud8e6uTzXbTU8TgVrUUkkMpo14BkYX42qlsHW175gIBsAEzM
mPx5+jh6g2NrDDCx7ubCz5wq2ASnWYYNzpMTiet21pk/Fn7g4sNJjmHTv0Q09N4K
oPV+c1FNhHbGtjBMGBFJcwRHbQi97yxkB6d9jzaGS5KfMHKxKtWb89831owcRayR
8I0NRzs4obpWmk6LMMRFVDVulprAlOILWfTI5cayoXYVVAaCVOkeEcJ3xcJYq6k1
DQ7RErx3+3mnmmx2SDajcoct8mvB/yq8dqp75lUe9aJJtVi9M9LyzwOnvPhpcOr7
uZ/wzMPjGPmSGriZZ1Q7pfA8wmXsUtZS9/Elo79kX5fwtd5BvqRBJ1qoj7/8OF0k
qa2DD7CrTAO3orR9EygEYvYlmlmA5VSUVrTKQod29fC1g/s8ZHwADfG1dTeiF7YM
uAPiOUNR9K946rbgUQvFYq3GlwRa4c/E0DHlVeJh84qwEwoDu2UTFTcOFKGM8d8f
9ARUGdyMs90FjI3O6DvPrPjwU5i23o+sm6n1kC1O2MColA60K4kqqtZgr/nBYCNL
ci6cfCduJbEiqPZImfSzX5Mv6JdWICYk8o2lNf6S5y8fLAIZLhiYx6HiJJ7IA/cz
orylppcYSOQZ5x+jQ4e59egsDn4/bFDp9ZHD8vPxxCcnKxvcPYBEfRiWiqaJR7Ob
6Ciq10oSK041JjMltbcNFvFv7kh/wM2S3cFiW8ht/h/YUkaEhMhg9pzs5pcBxZSR
3G4cs9vPez6hjycagSzNttO2wgYvMicYj5NMr3riCrhiarKFs10Vsbdq4jBx/RLl
xJFMYA/5mm0IqjyOAdGTbb3l/IFOgMN9fIKVfn4AQLmL/jYspilO1ORFZxaCU1ps
Rhd1kNLlq2Im/cPyqzFUe2gIwpNTiiaM5hkiOkeWUXepx7CNQDk4Z2vw6Tlrgwxk
5eY31xcvjAGHetJxlZoU1uVLWuun4UXPKpo3r7y26NdZDfCw/Kv27bP0VILrUn2T
gCG+vpTUzQcrv/HH3UprQrDuvLRgNs+uejiGRPhb9m4mZ7Iv6bX/8jCymQ/V1KlT
dqE7ULZ1c/quoetantUGMHUlcfK4ZpbdhGFsIrtGzwytDaxmznFonYnlai8c7IeJ
1a9aPtZ1VqzF8Ks5ZWQ4aeZn3vh4AB4+c5u85z+nI5nRXPZvgpT1/uEODmZwuuSg
dAUTkrYHlJ3VJdk7JVSUUHSsNCeb2FeflUBscZpZWnY3t2041gs3IU2sLjtzz0pz
/txO++mBXpC0Q1dS72byR3aEWpHJyHFq+iXmQL5BsTZaD3IC/1kQA49D0KvFjO4/
x5YWEjrZvrPLESbNvUrGQEuwOmo86ZSOfELVXnMD6+AABmCkciqfFXBKRVuvQzCY
4JKNsU1tHK3lgtXU9Jzx5GamsELQdV1StIHDgUpZV5YTToDII6Bi/Q2Bx8ttxjZC
aghJkFEfVagOoC+xF535kF11smcdNUjcbat3UQ9f0k04TJh60wYapt5vBSzx3qbW
qYYx+kvQfCuwl6WFlPUOZxP4wyawG48nwMKOd2PoGGOWDkemOblFQY01UIs4mYqw
lC2MVC8NktBbBBq0hgEairNTwy3SZJEhp/PzmAOPakyLhk4S0AOU0YK3mQWJzI+h
4Dp8xKl4fcbouJ5//GMchPI8R/WDUBXyFKd/NKt8zBOqW9Ocs5MaoBBhIhpwNBb3
b4MRN6w1YaXIhKYgRtkpGluDUO0nUvG3Kije7pEo5uRd4hjq56/aJrDeH0ijAZDI
rEvCc5Kd3sBzgDrVotMx2qYXO+FzFXIQZC3yKN2BjSIDnKXpCxVlP4KIuywOUblB
HX5j3DeoAaW5Vwy6Zsb6qMi7DiRFgvsWnXpeBfm/P4H+cu4piPiv+QcaEAGGGiK/
3KM3DgmNdzabg20dBCyCw2v7aYLfzhD3dNf9RpaYxVup248/Ip0omCKi6BmHyBi9
UwJLNVmZhAzJcY4/rrmSxGL6TsG9B74d3kd0flbgaBqUSeUzq5yMCu7awRjh4B18
Dflp9F6ro8kI9KaftO1FrwaWl/lnykQyKlIRiearrkNHU5MPYywmXoUl3gz82Jn2
gpArcLfLtE8Bml/vD0tuvEVYgb2Ws3jqeGZVBC6aMmEgslXGAVHWM62bWrjIuE/E
Iu/171pY6IBFvSYMLJzBiICRB1GOo3nV3D7cVWpPSDMfzjT2pOkyAdEG+ye2MMob
48EfkRxYDd2YCngCWebZ3NyCb6oVpY7veknU6iEZuqxDJJNeFahV6tjTddm1yVaD
6i5pnOqGP/lm4tEb7DgphCcUGhmO77ITHg3A0PiIa63MxyyULxy1ymRVnHLldbGF
VFNSCjTO0mxo6VfRDHlPqFi5tcMNfypyp25ay6pwKzXvwame5V+WCI0R6JC1JXdQ
yGMLYA5EZp4Sa38UseoAszdKNZMsNwcDbyGcIPe2LE30yLOleoAR0RwPL5jD8tNA
hPx4roWZq9zEQc/ML8KrIy/nYzzuoP5EydooCH8cdkYGcDNFp4lSEqb+Q0EFDLLQ
34kMjCVBXkMbcFRSAclw0r+J3JgmK302GJIGRbmhn35zjLLQMn7Z9NXC/fmnm5NC
KNqs4h4UDbNHBVNq9uhZZ4lEjTLIx3NMfvMZq8qIcNl9czLsE/CFeGMmUeOKJ2PG
lONxRfT6XodwhmGkaoOhY4b2kLeQm6eevxRBFzHIc83K0eJrAW1tFUpdh/9Yrjm2
9o0ryEGeNfQDOh+iq/jxcv858eBgMkWx+PBekaV2xvQx5j5NVjQxSby69AERpAZm
oSfJtJl+e2e9hjY+M0tHby7fRM/3r6GEDK7sGkBOMOAlsy2BhD1m1dqMsqTeZ42P
PytifU6NeaALpFrgZ6os9boN4gq+ldMieAOqDj8CJ6iCunpKfV1IBpy7EUA0ctXB
IwQ9kjQkjMn6DYlJ9T3szi69b1+UZVyfJ973iLYZKMCefDjmxJ1AOa5jwNxdE99S
qEow79S9riAz7eHpblZVSVameIJ0u+Al9FTpfO4Obw0nhNqifA1p1BA3qNTibKah
NteQVyvG0v8tjzUDvTBODW6c0oJnVhSExqz130wxTJyHIknSFo5h6NM4jvPVRhCn
ZKE5wUuY3GZ/KDiUbBmhbrjT2N3OgTFJ94bQnHlOk4QM0wNnPtqW+P2wVAGN5uFO
WUhY5ZlGi21ae+akD+gSG8KgZIcXC129E5jdr/HaOwfyR8b2Ri37sIewMdgA/KG8
ykvEZmTmWRtYmS9EeQOQoA7d4iGrf1W6S8tSf43IBKI9dz7tDkDMhDvPZ1TCcfwB
yjXZM9zmwQgANh47RzWIu8zsVDMTArnX1uzrmHTmJGhGYihs6pwNn5NfikBPD1km
XQ4dNI2W3eLHJLpohTF1T3xsYdfC54VHpGCUuFHkIQ7UBEUNQaNN9ovo+UNXNSrM
CxvowwQKqqvJ5+QuqRFFcrllozZ11uD4Txd6iRl/DNjlggbL5aZdjiQWiX34ljuN
0Kha7sX+JqVaoxY4gL4bCq42F1ZmGnrKuD4G5h+mSw1O1tFVxsMMi4nhZmNvzyq4
CAytDRLHwSnaOuCOm7Fc+TNoIZqhZkKUaoRJk8y9kmxI+ngFBYvCBYC5jNnMdWM4
33w8mo8yvfiDPP5va3q3KjDVelJXZ5OB1qm2oqducCTPJr6vxZ17UXsLM/9WIRDQ
8Jzjd/HqITmFGMkM6TDczIBVbhJzZXZV5C2TbIWOjwFB0579PVByXz93UUez1hdP
qPNLHOwLGkaaywBg2aIwWZuruf+V6k4hFV4LA4cWXPX0NdiA4rNOePxaZR7kDepw
gxZRQDBpiI7XZvV4+DQH1lkvAasK23u4+8xHgWqlDRxca4sDylo72wI6wpKxRbch
bF/yCmOSnNFPcWueZ/cemNvyj02rY6frFRJqmkh1Gu+iGq0HsFKz5MXjufF2BFaf
y4y0DYfRxyMG/o5se5m/xT3dRRlOkCC1jTd3kWtC+eZGeWETIYnT6vSqCGof0uWe
g+62ErOig623hiw/Uhc/0RBmSS+j24jrSukEP9FRAR1znXMryFGrTVXRRvN5kPNu
El6lbOghZwqam68srmCB8Hd42VZ4NulzTnHNuRAueP59HjAq4MOvc8XvW57qqTLn
GQyIVpu17ZahyG03EXuXu6tQY+Ci5x7XLStemSOMJgFip0GqmvGn7YEvrneY3mXZ
F5pzNTlG6/JNqBcsCKdERTeVgdr0Q858j+dgLqJdYugb0j6Vii6WAZXEj4/aYrWa
MyWNE4J3yoERl8oXtCVVBur9UnxLHRidAMx/evnWlInNqVcnyspRjmn8PlDT+XJt
tewaNP3POM8M1eov5IXn6ogThjc3WrXnB2DVF0z6G2M0Xf0sHqXy6W8Oi28Be4Sq
KBY4+MswwpaXhUrvqWHj1F1Qk4SLpaHyRRx3j50+ae1cOADqou/6nSoJtOSL696G
wZxv8MrT0gKjRzLdx5YZAyv8+N6xJ33dJJRJyZTGYQUruA+aWEJYRTLkg74kA9oL
ZX4Dp+hZpfsb9a4yvHObs1iiKCl3DR90RsmPcn3B2qKJfzVy8I470Ukwi04lCvF1
BE2lFDccDOkTOBquI5OkIWD+R5MhkiWE/xlOUro2rFAwr2kLWb7dPLfftS5zJG8M
xPOaGUXaY8pnbz1ozlEvOnCRNoQOv1yo3d7zQZX6afuFNyG93FAxHx3llL/Ti/d4
a91Sgj6/rQWcLB3AQ9qHL4UUk4maFsV1S1QJW6OyHTr70HIf6TBY/NuYiaWDYKMo
pKoa8O7LpVKChOPHH6b6jKMp8F7YNOhcs2erFAmAHeYbAJBjmSuUJNcSqbL5FrTh
p5QxbrA1KYgURlkII1fpQdtAXDAwC89uplFKeTPKvu50ddUJMI4HonMEIHZitJNH
4tqqnpInJiJhdSsesRnMDVXdFuBA2iAWHPudOdGVLqlYcgcCPw5216+xHngGSPuF
QU9mqqSYJwI3kyl5RTl8AQ0C38yJYf91O3/7XXwMdi2rq426lloMIhkI1X5Jg2NR
TO1ZnjGgrVFosQYJqAyE+LnTCTREX0qzECg5cMCzl0vV1fssM3/+39pROlXKGScO
FR9hLTUiRMA+Xf6hUuHws9RIjzn8AMGSFkEnQ4Uv/8HyWsr2xD0Soi6rNBdpaVm7
toSS5bYqxoIOTTWhePbhMxVxs7w6TUNLgLcsoROQZPdnGMXDSvJOTJZt/QX0F9LK
8NxlGsOH2C6xKITo0EWlECWVE57pqV0dnUXx0A7OA5YGiO6pkZAgiOm3e29jnV+E
3F7TK0tLyooO3P8rzyJsYCU1xbKDQChcjmEKUiFcP/vhkc43muYDEiX6L4joQS8K
Y3GHCfL/znXkwWIVADW4/FJ5dhmaD/4+JuODFjDDmnkqcArwO0L5CnuQmB5rOtZX
oguB8gCY6ZjhZVo0tfEZUAbHsWPCveYfq/EHHFNCJsQ3BBc0LJloKDJ7SH9ywac0
vyE7K+sxClncGIHBsSyb66J8E5uPcnbHBNSPYLPIaNBtqnfaDDS+7NTNEyVtw0iO
uM4D/7FNnQSREzjy2wHuWCAAuo2gzIYPKJdzgPphc8RjsOACISJH9Ktq9VsWAaJN
UB5hgg+n60Aq3jjB2lfT+MIoZiVoIa+y7vpmKSKBtLRoVLQffjJjRuNCMF5VqHOD
qoNm8OxgVPBtBnmfiNULQHygaxdxTzfZXZaRFCgyz6ZkhiyebkiqVmbBXrOTcIpH
FOx1UDEyyObm8A4R5T5D8RIzdWKyP59trf7h3p1thxmeTYyGgfsX6BtMbdVoRtjn
c0YAfmGkP1TzEkn5MFJrIr4LRNsTwX31Ofup9ZGW+GquisrEb54tTBE6w3x97/3N
RCa9YCDIpnyHrZnRcjOiIgmDFOHyfQODKN/a0VSxyJWx8pde7ylVuLAgYeIKigqf
HVKHVYY/fB6peTVMoL5VzX/VCYIvOpXscE+h0mZS6MzTgsglZ1S7FHWtLxin6wSz
ow3yIqDhES6EQrQsxeVnti47Wvu6vtWTLQVnwo1W+SlljYua+mM9kgP5snfiFYV4
qrZzu0Y2CCPauGRgVl0VimhupaLznawkdixR2FKFDsT0E37yyEihwILB95WKT+Zm
QotyHOeZImD71Xnag44cUwmxJmDaeBK1T4JWbKxBSyQa2lVDnDyycilUf6ubxakR
beDfucF6/d1zKlN10yBxnGEP4s9k4LGDhZkff9lHGOacEkFd6sUdJNicIEtRLXr3
59JKnUfSSYoQ7zsI0srdE8/1sT0a2rCCzxEaJalfsPh5Opk12E9SxIxgErv3ZkMC
J4KlBHCYmFk5HI7nFYlGjf+Yqx9hQprhGx9UFKAbQhmuP80z3ejpkKshQ/1vY4Vu
skbPrlyXgZM6eyb4qsc8aD2P9LacrBcLu57MsrGQSFeog2DFOOc9u+c68TwDDD60
IU0PaJAJWsI7B+mxQOfv+iDTX2lM0YE01/oCrAEqu4Je/Feigfno4vQDEDHKd7ho
FPDLE7wTaVqzUZpVFlSScTqRgLFakc9YS5fXTp65PCtXOV9i2yBZ5wPRfUoELe3/
YwjFQEYHi0WG9wb7NJbo4IPXSnvXPKtB9XUvDj00R9hc13mGeOfl2RuHAhwoUBlh
oXiPutrJ4aIO5+vHoKUUt+rZZMrGdWrCfqMsKTqz2/8Xwz3C5BWbfU4DCcD2VBhB
J06BsZRebDeN4o5Il6+tXZ1639iQvrSFxl3tpybHvWMTpH0LAl7H4dvvakmkFZqE
qYNmSqQMev0KG4thWfOSil5eXxT6Gxo5kctuj0XvUxrOQhs132hPseHwtDO8RjzW
Z/5r9uDNS+nEmG6CKX+FcVueWuxEMIqVashl4VM5WyNz4CePVTcFQ75xXhkal+Oh
zuXfZSq7tZebbtLAg61NZPM/e+V9ktFxeqroB2/SW8cuD9wek7dxRidZwNiPkDzt
D0sM5JaATy4OoQ+M3rp7HD3PKZZ7aaFKIggjO+FK5F5jbSIShfB/PQ9uZE31cb1X
8RTpl+aZcSc8AyE3mbhOh8ZFpruQ/Upy7+S7692aAehH58ZISOYGaA6fV6mJnwwS
HYZ9sIry+Ol+hhZQGydJew3QZ+93GOYYX5pGA/sXHuzQgN0GjpseltMBNJEi0YIg
BErApuJ4y10ckZ0dqeipnV/giqAMFjOgxH5UKoPnfJXLJWDZowfm5a4I9T2UV2o6
gifv/DrbzrDmSdKz4UzbMyDLbwgrDFR3afrPAvPfZrAS3Q8PzRJK+bm31xsiG8px
RDuCTMHKaHW+t1CzIh9M90CrIe5VGwqsNhIK+S1y6fj6iIdS4Sc6Sk60Xpbqxgw0
zdBvIL5lf1lug0kTSeFCnAYBIRe/QtpO8rHfJDlqA3/2DCQ7IqdK2l/rgqTZ2hJ4
sjTLw4zxkbDGFxyS/CoPYN+jyLLEQUe04vkPae6XzGbiQoCOK8cOsvCsrcXQiPEC
ME42KIZdT6P7CvfcfdyVX2R3HpNFylJbWTuyssHRw5nRQk2G8H1eTw34VrUxsqpo
GpjKtzTR89yLuAaWEYUAepJ2PyAIiuNcJnLmFXwiFTS1g+H8d/TWIOAT33aWzEu+
0xhwUIvWvKB4r0dbi4mawbpvhUJVKGOdd95zEzmDkg02K35DUVvEy7boKzynAkas
QOegldpD1pxiP2LvlkBA5rJNoZAShPP5uBKO1wAlUPQCleN1U9ELhE0LahRbwiX4
jMMT69wZsew5xIdMhOyc9Hxbkf9Et1dLXmJXq+bxECe3zXIoy0QRM8k4GScI5pCg
k3hL3T5ibXCpPa9335AiZOoVgu03eSW9lsnn+zE1tRh7OxZZy0sTzps8IWAKxBMJ
klEZwe8ATK3H+oEgLhMONNjB/JaUvoNGts/Ac1SBZXmwhwVuqQ9V+5CGJ3lHrwXl
f8WREsrlSLpnc+MfKFDRmu38ArQDZ+7AfzpMpztFtbHgIRwJ7ZpXoBYkzKWcRKNv
3poOJFCCLkwUDAmscArx3HEXG3dt6s04MOXaNM79hKBHhFcJ3EFS5I44GAmnuyEZ
rzkQeABtosDCUMFAJAaYFShUX5Cj3/A+E/on0PsAWi38PfwLFyWCoZrY+s66MlYu
g8jowaqLf1I1DbFuglLLZRTMW0O+cVlO6JkNPebp+rJVgTnccdPgDd6wQudUODla
+h3PImgpXxF/tRU0cKcSrfmGWz8zkM1Bq+m7S4+PdLgU95BAlmC42Iscr14ZM68n
USSJ/nPwcmeuri8nxg2Ksv6kBRBbofPBW/PRPDKs6FfJFpEuNd9xumEnzyDS8zgF
TVK7hz1xb5UUvqhv+6g7wAFJNxi8xNr0hdQGk6IfU8A5aYxCrzXkcINps8jvz+2w
FDDSuAQ44Wk79gPChBt1dFgBTxHGeD1A39hTDoI1f34H0iHlba5VxBFbBrkcu27N
j7n19ZGh2kG5vUHXRbJh/X5Z9vlmtC4JdUWYvshtz4Wz6t35g/rWYLmblkfkd8WE
HzqDTgc3f6z6NTf4DkOYrvMHRGjzaexKEok1XQNNiHt86TshaWgSjKELtyHxbOAk
ztaQRJG5amjgS2TgkgVj6xbWCgkCOEKDV+vuAgEcwjBGhSIQ3K2vJwGyaMvSa9Lf
xTGq6wYdAq4OQ/iZ4twvkl/GSJGC89wdd8GByjlJLMEwx3GRBvRW5/oH1tfm+mp9
jnq2mKqdA7u05Eg8bjl1NNo5ZC08ZvS8zo/om4EXe/U+BOb43JWpq48Z20qyKrdN
2qm9Q9i1xb42aC4q2C+Da5s/8wvVzfO4Jp1gIw1E1AuIOqzof2MrdCAUYK+uMmM/
A8F1110GKOyo2JC0VxWI/HOpSELGo18zeusyejNDXfdavFA/iivsLGF4/ZDiuctf
7uEf1NZaUg5RWKto2EZ39cyuHfhbVjvaomI4BO/2Af1vMVBPSv1q751CYhM+3geb
EPZeZf+xCEdw9OIXQcH6UQpnfhHjb5Nc3gF1pK/0s3dpw63gpgztEkOOI3IFWJPr
QldI6YgkFvOE+xWUD5SPFOvr5vLluNsCTVP7ecS70UgYRXMHYgP5q0MqgnLkOJxf
xOrFoyy0pasE1Wse5GQ+fa5FFF9+98upG90L7BV+2xXujcWRIiorVoRvp+nNw9vT
+uILMpVWmsl5iqkRReH2ci+jynzKzgLa67N5VqyuGPNGzoQ4Q2e3bdC7ksGywTDM
ZLXAWhKHDz15dF+AImWqCuMqUsZuDn9kqvFgLn/hcgYFQhzqM2gB8nHYGc0/GnI4
WcyiVPk4PMFLoSsm8i9hbP1qaAMJqpuiSHNNRIWwkvZPAmMPV457USJ1E8Qp9x4B
Ks7UZDJu5YUJui9K0e3G02t+KmQitFE85cXS27KzH4HWplVEKVROllZGUs3Z/fFs
BQb3wU/QIbZt/hIHnyMhlj9J/0/c5S9zOwXjGz+WYIhSiY8O0CEndFIEbb95S4rX
zyxRV0++N4OeXJVZU0i3iHKbyIadcOJQpy+DLHtt1MPKzhVHXhGitGlyb5GRd0jC
prtQ4oMOYd4R6a19/g85b6+CvBy5OVKoesDzb8Zg6z5GSEqcti6tLcYspVg08Dwp
d62de5A/AAOysSFIp1rKEzho78TW37p+Cxf3f24KvE1mGI5anqYM//UXr7fXe4/h
GV5/d5vVRThNkKDkrMFr7uKEXyy6ke3Zqs1/+RzmyBQR1g7I+XH7sQbSNgzQI2zS
HYHt+/X12UF8fSO9Si06SYomp4oqHlNgx6D42iFRFVjoRv/mM3xRnhHl4audz37X
bCClqa5Z0P1vSZxHGUe5QI5baH0qEGGDDUkszGfFaAcWQSkNqDV06VL1blGKJ0T+
CQrW3iN+2uwno8wd3VWkeBvd5gY6THMbLfqvgJJ4SWGGTAG2mcADmWxF9E6qmiX/
lq22/8XkZcg3iJrK6o/NEUKfDoLLqes4V5SbyHGNawvZ+IbDB0OS+TzyFc+fa5yh
pK2v6e3rCYnUqydCy8LMrCxJwXASPE7sWeIiSBP5QijX5cILDqNKJ0kgsFBRhgu1
TGq16U+AyoflzWM2t4Mf/laLlf/v7+7C9QmGrqnNDRiUJFYnRLXJSz4IjiV2Ck6u
RB0CW8GHaaGyOWY+gZSBmVNADGZ/tATseCYfkNJNpoNpPQhHBK1XIb07jYqd8CUm
J/mJfwLmEhA7DkaASP13S3XzJPQuWx2SGPGJrq0zifzmvxSzCmsB9zwAG2ua3eJm
viPffZCFypE4SRb0u39a4+86vhBNmmVhkQybFLW3X41C+rFIVFub0Js2ag8Wv1ZR
USOoqAAEywvd5WuuqK3jRK5TDnmolL9QEM+Ha3vEcUEXCYMG/1YR8DZVtEJ65g13
16EsmTkOiS7dudYplr3ysPlwOoFU1iF/hyK2EgB7PypX095kFg+ugEvE0DryZ8w2
jiOcvF0RVvaxJOoSANXXkjpXSQ8V168EfwefYoM4uu1zrYV2LdWWFgXFw1hWCJOH
qpq9r7XS/BNm73GMMCRnLCDmCU/JROa4A1E3O1IqPZkeymN7krZs8pp+JogmuecW
IC4sJYe6+tFROHvrBD6JeCB4Gm1Q4w5eHxgKPfZwQeBImxrjebRGt7tO/+Kw3Xio
bkuPobOAfs2qioa9FugFuma/8kBx+UMyvsVvv7vnSfWofhHra4sCT6Dwg1TT55aQ
WMJMjaMJMqN3aYaKHEtvguxcB/YW2Vr+0Iu7hDWbOU0mZhhiWk4QFKl4W67AiTAs
pybo0Ya4Vr3+KlYrfWzz1V0u0+noSeoSIF9ETD46+eZAGF60B5iWUoIUQ821yOP6
Fgo+dMxT3vL2ctI9VpZccXznISfpKq1Obhpn8Sv586e5IibNtdJ7ZhmsZ+MpTBkP
V5WJR/0eqJwvcY4TJoqOnXHBx/NKX6ZjuwdhcCGLJtSnvlk7+zUQwS+MB27Us9ou
NAs6+tB1lJ0AAtep+PB5TspRIgSfqssz+n7973Hy0/c6xHfdoYt+cQcPSosFTpCo
5W56HYGGOaKCRWmvyFDnRMm+lQDr99FM35w/gbkfH3aXXVH3fpCl6UCHgqHVBtx5
ixqtKK3e+fR0lctNri6qAIUIRiWfAuSCRM8kT1Cj3BhVxo7wPi59cfyo4ABEY6v1
KXajELikIQVnEIORMko2Z6wueR+eh4UBLSe0APbuxD8fGekngWny4esYswvqyw7O
sn9phlXncZk2lSRiq9mOK7wfbKqqw2AkT8+IR3KutcvJOztUO1bXZeAP9t/GeA5T
DBUTVjz0nwrvTBQNaHVmnl7lF7y8QEClhDT17OtQvPfYZ5JYHiukFO7PmphIqSOp
4wyXdnMF3acUw/NKoHNx74O2xm+1pBDhPPsBmzzW7cJ+Yqg8I5ps5BLVwtuFA5X3
Y03Vq9fR7xjj4JLz8sLxs7/x01RBbOtZE9AaD79oJ7bZKRs4eRKCqdW5NgtunCa4
NYLEqlWcg6hDOCn4g+A2Rd9Cqj4dKPaKiBIL2VSMRybuP1wl/ldPi2tKHURmMJRB
wUrDxMxHKrygStgP40HrjEJRCJ1SiOru770DlWCIgUiznHwKOandoxAn/NWCL8Ix
9EyDiYcsHHub+okULkC6MVT8ZHe8kBzFvlS5rhANP9lxH0n7t3+rE0QU2B5ByF7N
Y0KGXeIKHUVwsTfPrBkY4G6zVazriEwWo1F0NuQ6ppm8xEuqDD/A1ZHVPelirGdn
CZLcEgysTbq7lxIgQUDxbPZvqjRRuti1Fjx9n1yhTBWlCySQBx//8aqVxAGPysb/
3AQiz02LTF2/5BOau31rBoRRSAnhoOZJ5Vwzj695+WwxB6PXxHLZ6gS2b0hlTbBH
AqmPAtTiGmO+lokYeghInwXFFl4sRj9/MV26ajmozjZ/pcKp3uAbvnc8DpbK6lSL
4eXV9bbHYqZy5i1U0Ua1iy+aXEaURpssn2c1Sg3rIhTeOTvrPnOuqvL5eqRvtmoL
l8HwDzYNlNIGUrLaQFFeic2//aPeWOuEMlLQSajIkMf52Hzn6yChTDJ3bUhefj6L
jqHVzoZiCXQguZOHxmX4NH4GlUjzwBqX+PeqfiHe7DjR3K2d9mfLetgMRZtL7S/w
VgI5xUhVwWHlpXP7PrY9ZgmZxzuyg0n6D7wX694wO4VwnjK2CMiValSCX65qMr5x
pT7op7ONem9RUQtj49+VbVYHI5gclYw3sdZv1OaSnSwF5l40rfsY8QuwHp4YOLy9
zRG4H5Bk0j7/E35PTf4/EWSMotoxbTqeiGoidDKpC0myrlkP4JPdZEqIM3cvYdcg
Q+AmuIjaunplN6nAxa4h4i/PGbd9fepn/ctwp93bnzM7s7Q+OCZ7ZonlHM1khqo8
1Yr7x0EBbOg0TchJpzH/zH71YAAdCxYBDpHhx1G1BdZwJVGCI7x5MbYSIegBug7t
wRlynPiWeeW8OlNibtQZnhui2QTAOdGN9WalGsXUSv4qnqf70rKOiWJ8R/aNnu34
d4RwHpeQHJw5qs5UYYb676HWnZYQV5s4dVxZUGyPy/5sHAP3rXOgVcDkT5XUTlya
hbPHc0fRMoqEAMTPllvWdf17ehb87Mzxs4x4PKEs6+KVcrYR5Ide0UJx1pfloyPU
xLdJnwNcVpfVoKcbN5JKOzFxh0s7liw2fLpggcucr1GKno9ROkhhz/FQS26KAkwM
Z52gys5mU0b4uTq2STe37cB0VHlonxmDuU+8FLpYLFs7KUAS9GKcPT46XL/Jhw4o
+T1FsfIjSiDE0r3Hnb5T4cWUl2rnTHsBJgCG/i67R/YHcZO4aXzH1v/ZSEqeIa6L
F5iJu+l3jzQ5RR/EON+kVmTePhb5wGzpAWucwGFnFRt2fftW8hKtrMF80TTnTSii
IGlYN/bcSGmhuw3ad6sQQWctZ81/MLjuQto70Lbx3R3sHpOUtAuUlEKjy+9zEkZu
fNVsHxfsYIO3xc1zINUHvEzQPICpwePW07aYbJxR8SSHfuzFUz4tq8ftjYMlRUTF
6QMoiCn9ePvYMyFrquiRFpK9PcWa2q+vQMZZq6uFatpHpRTIWqixR5P7sWHop83T
hcyLlvY4AiuvrMywSYzfzxeEdlxpUuDeLUrWd4BNfdphIbjnsIiXIYHq+D76O2Wy
U4YimEtOiXa1MXaiVkudrR7pVehf4qNDTPjoo/mD5v6E0FivegG9k2VND+QQZeED
a1983xgVP95G2lhZ6NwAulKXPWseayJZ2ZKJWCoex67MqEouDPtLRrrMb5IDh+sW
W8V50h9TGkE9IunJVTNCTRB5Nl97qRgW9hOeOWk1pe5Cri6NvUyzGcG1BboG3/ie
NKJM7e0BS9KMHz3+mide5iIXK7/jm8MqHbkgSYrf3jRqqqjbO43wHTOiaH4ZxmnI
n23dz23geB3yX+hy4nSiZtoovadzbwKVa1BbS8JgyUxwDNiLnTrMc5KPAWRAbdk9
lyQymwhsdTOfNzYX2yv2V3h+jDpbCTDjTOpZg7W9XoYYNYtr1lIBf9YQjJsfW7Iz
QOWTlB5MKUNHIEuQ9av4QEZaiT5nuWP9nvytEAqnTkXtou1YxiWSPD9Z023C/Sue
bP1kwFBYdzqhzQNVwDXX4XdRiw+77LN5jqzQqXsPpIEW2rONyjAvPxoNMqlqyfuj
l5O7j2R5JiqEgG+ZRcryF+NdXdmn80qaVebQL/Xh27D/HAWQcy1e6BXacKed/EvN
DmJBWepIPieMWJ7QKzW7t+7RjzK5p1mGZfLDObPDu0gfktx8APVc1yt83Mxp+Fsb
xn56jsHEcaQmaRvUw4GyBKCsSiM+N2TPuQm1qZrWXJu0rFqt0Ilv/IvoYbnJbgB0
HuJ8aqziR2YsGcGBDL7NrCe1K6U3QFnPyGsp0xbQkCwtpn2tVv9qCrCApRpYJn22
akNF7L5sb5bgFnyM8h484s4rpV/d683kQT3Ja4hl9S8twoEzfLLYp6Oy07Sv43am
98fukUdJAlK4NbAtNS3ldclR16Wp7QXkDoj2Ao8x1eRk8md2LMwtoJ+JSgAzfye+
AV0tP48GDXWiJAVzibRHYakZ3krfkuGM77gcFDC2TQwDBaDDDeuSZ/MeGQqan4fc
cJnSU1KPDR5dR2k9/ioEBQg5Pq6paAqdZw0pZ/JzRr9hAeHhqOXKrH2OS0ThAVct
btqclWyWtOqeSnSOE/bGgasdmF2w9qMS7+KZursP8b4M36UYVnzdge/LE/eF7gWH
qJjAtqI3oe2RI0+RCXliaslTgvsRiwjv5DaGuK59tCtbnLiwUgOltGmZmSG4XTOB
hjDcDmQ3XC3ZMdwCqcd4hS1n3ZEg2JvLaPh5dYt9Tp9UTQOxV10EyZzXEpJIE00n
LiuXKjm5YHH/vdlVHJNpaHk32KvwXaB7+jpYecUkTNMrDJIhs6eSN5+pI8IrO7n3
ahbOZn/fySPB8nGdmWqN/2NDJcKfhjn4CWkrfoZedhQw60E3n8LcMVZ1LQCjV+eN
FvvO6nYqVthE9TcUFj3+rY4MjJQV8yuAxeTkvb2Eji39algov4RckW6mqS9q+pEj
pexbfSCa83GZ0Tidyz55RUB5wX8RX45LekV+kP6DrsfqIR9xuau258j4Ff/EEusk
+4rYn4edrgbcuhAjgMkYFa1UX3HWUzpB+DEI9ldliSrfSLi/B9AD6zxX28jCoecA
IYa0NooF+ZuXO1M7HxJZwiQSRLCbvo8ORzGPGyvi+otjO8XZS2fqDRaZZVmf0FA2
OeJLRKaNblw5+nIwNOP4i07usEhAjXTtjd9D3m08SCdw3Kg/IWeDfHFbaNMKYNJ9
UT2/CI+TSqdN3VibGdvS0GGRoxc0RCYw0oYp4zKNQeImBM5Jl/MiAQIpxSIUHr4D
n8YOrnA1sUlthTIKSr+xmm3RITi6+RfCUdk0U47MEGcSALQ8fg5+5oR/hqA49hnq
XtsMcCFOFXRXwC1QoR3kcQN2p0ytzk5sKz2a2sqK1DVjU+SF2X1Pq6SXmionRGeZ
xdR40DnjhVejXfgIKJCXX0b6JNZMKgW0zOg4xoAZVEfiD0O5jfoQwcKgElejFroL
4Ge2KRFdhigrUZl/mDYJ6169p0U1eR0Fi8YbgaRmkOvs511UXjNc6PTQlm3g6E7a
XOBnHn2aO/aTF7EHMHjmhPoElgjjMLIzd1NWJ2M4Ma2kDX8/omPTsEcd4WxL4wY2
uuBqOJH0ul4GxUJ8hSx8hgxrMQBaVsiF0c+p296LYwP0ya+Gc9Fxt6xzILvPYCah
Bpq/3KpvVL+OW6+xFv0fkiSYbNOOYpoRn8LdAetr2xk5IHjUVbzmEALbVYZbCQxR
7w5qBihDSp/turaut0Uu/Au+GqYyslzTFaRK6gzNmpKFiCb0Jo7AWSiVqPzGkW6D
EHnVj31HXNPsCcY+x6AbuFyjcJP7Aax9bASA6Zz5K9GOUv6tJiRvNggulVFebnE3
EuL836i61M6ns0UA2G6IxmJVHB+aquY1+7f14qJ1Fp1lPSI67JeyxH5yZ6aohWDJ
MkGxv7/AiSQnWsd7op34ilZPSdHNUNTxLbh73HLu3cPjbyG5ktTEJlcrp0livoLb
rV6zDmosf5JG9pBI0YRwYIQBDiBg3a3BrD69AqYeYWfJoPUP59RIwrFBKFTt6LDI
CJ/E5iYTUy27HVJRVLE529Jin7vKFYzprYlHkTJQZpu9hIOz4M/gv3/+aWkO+12P
dloryGkt1XkcSciE8lXv0aOsQDfyxjWVX4PHvHLOLLNQSmqRiuEEv5q1PJ8Wj4iK
Co9ZSCCMTzyp8CjFUjXn33hIxAtXriPFoKNQwc53IDRLLLrIEX++tqLDdpyS9OS/
/wUO2MUA+QvNkMewtmgnjVPx4PDwmPL8WpPQGw9EFereFvuaSHJad3VVXQpfkxjV
IvLccxyj/kLEJUj3v2b2G37nhenwj0gwChWMadoOANxQcWCU4kdQDbOpgVDIZpfj
JvVmSe6onWCg51YRBVvrw9SMIGRjD2/f5OFXk7dhj1cVDVE34RVFCn5MEFvG62ZS
JGL2G1fWwR+96GnRu4e/SbfxsdnQ17Bw6t92i+vulePJsvo8dbjDN/uK5mkJtyzN
u/NfORvucAAnJiQ3AEHnvkKOsJbyekXZ93vvOL0+u4fCkuwhlOf5qptcqGdz9ZMn
1/A11xc8HOp9seauPIbOH2S/zIqP7OyiFPyhv7OvgloharDQpnXT7lDePQwrDlWr
161/05VW0AiZ8fl9wa+cN1ed3UP9tnOJrUZO47SfDE4HWmz3Nlb/a3Z1HWw6KEZq
grrqlT3LCwp9WvIl+wpYMT9udUBVlBrZWYfj+VwGRzf28n6GXGPRWdq00bmoNZYj
aYPuYaJauW8AArfnZFFsrvqtqnfMgO8fSXkcHS4yBpVeoaPxGnCGhqIzfw04WrGM
jWvMNk2FLlnZ7R1mcr2f5Uy+MniKnL47dM9U8FUq7tAreo74dqsAtBUxj7xlCy0A
UGWbexZG4HWOgB3xg3B4H7NMxdXgsZawxwir3DIj9AOyXmtP+nRXqU/Wo6Pav8WQ
n5FOuXXrIFDe2b3sAN+TPeICHjnGTpi1TIzYuJXp8+TijA3evZh2+KKnDO3z4I/z
w9KiChPag4NlB59OVl7R6KlEQnYMHvtElytNrguigSjU+E592QaMV0jZFY2Ao/Rl
LKseEty2qtKEDCxs14898IurS0+bIACaxcp+nhezcxwzZMnWHzGEgoHY+NViTyxS
OFEG0Na/KverR5eeKLbJ17k+tcizxQJs3KI1GwgF9AfB8RrlcMXAc3w5dJIV7Fn5
aHju0X35H9f5lxxgeCN9y9+l2tX4pY0z/Tdmm8o/lf69x7XY5qAO+Li0ytmxiyWs
ORnoQ71JAxB6hUqtH+RMdWoij4r8aLKqEs/T0lA2seCQXnLC1Y8V4mCv5mkUoF/y
qo2ZaX6tdZ2xlqjjdmro31eXR4BRmy7RbxlWinedcFsxB92KwlLSyYv33zlUGAX9
UVkWDN9Hru+aKohq9bgZWN3/nGBP/plJTKSVxrlpeDVjoVDdDEdWC0kcrk5QM+KG
5+ancOa/qKb3i2W8UtVllaimBG/Bnllt2waesw6GGV7mrQ6vAcnHDynF6T2NGInv
gscpxb0Bhr3QUKVpPqfMp23cTkMsAQuMAql0XZOYZ0g6LMEcBlavNno/bN8dYk7x
4P/yHKxB7hx1S2LhJbb4bhYOuBYoSG2Ada9pM9H6qXpM0vDw/jO3jNuG/1WKo4SH
zDVI49XVs+ykGQSu8d0aiWTBtQHK9jZ9ok/7qdiCAg6j5wHBwdoNzyzygLaZD5xR
99BJ+WTEXRNdfo6s8f+rB4d2rk7rL6TT6dvn2XXhPufno2i59P7uZ4T9GF/0d0f3
BOscULQj665Sap37QZUWmmbNMwBuqkfmmp/05px6MwZoIcXL+RGwVsTbP/CPq/f2
eIeahqhQzGODbpUcQRXdt5xAj+8bV3AX6PVPs6oU3FGBHBGT+31m8Tf5jsC/43pr
tikW2k7otFAh+wavXaMn+LNM6LhQlbzBl//ceQ6WGkv8pRJpRJL+GWQESiYTRkbJ
IpBhZhCc39m4Gm2f4g0801uodoqQlxuevcTJJAF7KisPpVFlANn2H1V1W6og/sNs
5QuYRNX69sFGcm5JjF0Ia7rxiNd1t6WKMMwgrqLXsbWUmXO6GljexIQAUVR7osqs
eIMXKyMT1XYXPDrIuvwJC8fYt67mfe7Scw17tjF8hnMDms0rq72w/A3PhAPDjxTN
mlUsUYWH8/GR135AcH7OS3QbtzQI1IZt/uLV8ZxKrymoHr76iqfMJG7mF61uOAg2
7byCiZVVIVPX4VKnOft9T8l9gKWzL9Jly/gPV0drpzNOoEl7P72mNIKR+NnB7iC3
w4IAGA/8okdnQJarjIMwFc8xlpQIBbY/mq0VVV0kAc5OnpcnNXQNBT0878IjJnmv
SYhqOontiiKr5gioflE2no05awrumdma6bHj6/rg9JPQhcIh84AuLSLFCRhLEz89
D9xHzRy4Gb/bfR7/F+vCDfsLbk9D8iS1lGlJjLv7Tw8eZmK4rwjWhyFWHbgNDXIW
j9xM3L/rqa2zuht6m4IVsye10eLzJFCYtjlWqmWEFcOudd7+BogdXkF7pXeHR3NG
VY/PtkZ5ZTaQZbjCORv2zNR+YAxOOMHIH9ME1STZTu3ojBWX9LPwWR4DzGlEGk3r
oFv/DEolGcj+QGIDSJrxVbJb0v252kXbn/pWj3Pf2ojrVG80GSSNqJKvMgtTLUQs
+zKJNPOdef4GfAgkBO4ZHmEJKKCaOHqoVb5DzO16sIf5T7s7ocPk6/kNxVApT2X+
7RJupcYoROA+qaLFY/DJYcVf4SqbP/cAnUxyD18pkhrt+RiPBWmdGBDwj3QLhfOo
MxyoH1Y7Ec1nqzvtfiHiiFnzrr5mU7LK9UJNe6pZrgzXl6HlQu464/bYu+6tq+BB
iXLWpUYJOrMZ/AWpJ4dIUD4Fu3/iAaMODDmpXjUyyUzmDW13oZ+c0jiN8eL54t5a
AWts8Vz1Wq5sLVkLQxeUEpQFJtLxUOkL8BhHTABEFynOfS1M26JP5eKpAtqSMb/t
4/moWEy43nK6FjrB3UMWjO//3SE90WEPBF+k25M6LSah7VRkXSUis5I2Ys8s0ngI
JZWO+C4i0tQucKNYYy66/G53fzdO503zh6qgYswXIasO91hbIKm1YjkCUVTuN/Li
HvVFyz6kWwNTYN/0mAaYfwb8Rew/bUiZ/XpjWZ1L6FDM9ZF+7b7QtkaMOUAMJEVa
jiBdrcYNWuStkZmQgv09KO6fkN+lcXKm87CCOz4TZpA6yun0B+yZ3Z/mTZFnijrc
ga/3SLA8Ph/sUXfm8Y9YbKkTpMVkh2hclAXHZnHn5IwmkaB72HeIwdFjikn/7rUp
ApzlhkwtYhsXqh2f/MWfaFP5nddFznl3uq58GAtXe+ji4Z97/+F3ppRM7OnnKN5J
tsmVK1Jhe13QTzuERmt5vrTjJejI/MZ7v2ic36nXq0fQqZvnfxQUQyOPT/vRjh5l
7f9tW6nCt7V85VAH+/+kOi+emc4fcRmRSMMWbTBHu+qUOZIu+Zpi5foFQzYVSp+z
wUI8wo2lbD9yCz7Ek+Uo2xTTBLIvIR374R70/ySKO9ZX4RcQevh+eaOZYkPXLFPv
CK/GoF6UK3pEUFoQQAYnGS7OBRZN3As9OBmfe/60+czMdgsF2OcrkoqK2hkYRz+n
wK/91ks9m5XEm+oAX+BmxppsaBL42FbjLY32jYFopDbvA6Ka32FTDHAREDrArmq1
4WCFSfu1BoFajuPa0KA0BfixOdI4eEpNj3V8e9Vauychw87uac4NPP9Q5PXqH/i8
MBvikSOEuu+yz0twau5UB8hyOB4+sMXWcz3/QhScdW6MJI2QWeywkU7LNrtb/QSw
qNimHQDsQuZqG29SuSBM+EELE8/+I+3Em9846UxDL+wnmD+W5/UQ/x4HDhNOS/x3
t6PArcw/6NC32HjNzV2iTjgcSAnwSu992ggltKFSNMQFgqOXdgUbFjnkwYO/t0KM
pTGaZp9vklv2Cy96aPLbdd8RNpiIrhfaU6u1WgKJ+tNT2jFg9CQgpCJTve93NDiy
AFast3jgvNbaWeBNNcchO9RlQqB5XHC+t1aQn4e0TMC93O6K+wYfOfe4vNJme8s1
vjbLYH/iwaMHRXjNu5Vg4QS0Sg1qHE6Ef6W61xIhCLUM0Adqp4m53AugAU6YLteX
YhwJpwjFKu4Gg7w8wF/RCTvVF7awUPZdQ4iZUh+vIJyE2tEMmkFlMUkgsEb8xC5/
C4babTH7YF2zGRVX0xYC9S2bcvBd56HhazAp2wyQzEj1/sDVgVhFGloSdkUAeZR9
b4sTWnpsDQI8mU47QH6G3brWnz0cwZVknhlfnGc1NBtgJ1Qe1DoxRDDtleW5eoTd
AKhZwz1yz8qxCHUYPrT9OOP2JlZ0S8eGH3fH8Rjg2qg7qWtLNidwia/RKgJHqB+E
jSQxZYTIePEogvBZrRcSY+FkN6z3d9wOSst39khiqk2Y5U3DRAddrgSdgwSN6VDm
I3RLgpEiqDjgKLb7hmjzWhknplDKPpbXy92PXmcvZD9QmiY2/LQ20y9ofP+cR+xe
wKN7UoVuJDGvB5ceCCiXIzLsBSfn1/7gJmRCJ61GgfA8sphmbI/JjAhjZoVBWfM/
7OJB6+VUd6xaHSOsIGDZwqrX2Ni4z7xgTQrm4Hv3RmKAH7V0DX5wA5BYN+HYiW4l
ZdfPb8iA+UXatB8hRGMwkMVJicKqgz+YyOt6YcwljmDszQ0Qm5yNM6+UKJtkl7t0
rBrkFpZGRTQEcCe5zPDf31K0GmZD+xKv0LB0m8eN3Ro9Y+MRP81HMyJ3cPEsQqP3
3URJnbfaxw5LHdHpm3YOF3TLaZirltBjM8u481eUPcpNkssfFbs8OUC+FhmyPeqG
rXLcx1GGAn75RM6fJig7xZvK7o2W1auIbIryu3/z+XQCBlhEACaM7iOv+yVPMtVA
kx8GDm5kLyJvdX+XkRthi5mMmeUKZx/rWJrpd1jKiXk=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i1bmsb5On8Zq9187cUaVKkW8yC+ohmyPsbENbfCEwm8FMb0F+2ZRI1nMd8RySECH
lJn+fTYvhWZYbtge9YCUIxDzue2Hkv7FHnsXAjnQcSorzIa6wXvJ/xyu1mygS0kT
i7w1MJn+6XwDUGawG5QqwWGRjZEQgP7G6vKz+7mqaz0RGZKhfrTXbPN/hGAyrbl8
BFR6yGQLfVX0ydEXWaksL9Mketfp+fDwkRqwDkTmPoW4u7RyjQSfmMyvXxQfpK6N
mI9y++gvqnuGBp7PBV5sEvu8pBDr+b5pgF/u4q8qlZK2Rgq/2DbD608qgijHQXWX
9u0HKqgjtT1gZu+cPSm2mq3mfvtJN/ZfcEVXL8GLj5L3Eci20QVF54vV3XaVTokK
gmuJ5BWrrIGoXQz1W2HtZIuoshej0UCC6nVm7GnyPNlcZxg72KRO4lpPzE1khIkB
Mo2xwg3Fwy3hd5z8KT7I6Q8QurwZ6gi9izGXOAxlPh53hF9jErXfNSyZTngNHeRH
o6I7SnitesOi+Djlgxns8RyJ0uJgpgWmAvcdC/01Rwgj0OGxoaUeBT9yyhI7p+ad
/cZ6oahfaZ3dl8K3zw2qwQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O8rtBifX6TRSWtoUEp343yVCxzlBXQyV82f86fILoUMd4nHJ7TBLZSemQFiZvrO3
88kz9786JUSnCoZlD+v+WuUedZH3s/vu7qm4i5oCXxIHpY4GQcWbJMCWrWmiiOdE
cV/VcL71yF+y+A9z2cHJl/hZaFhE2hAahMP1iy8RaULuqWFAL5lrMTUZvgvBvUal
OgNVqf6yxZbBUqKmxWvgo7BsvTvSiacpMztMRt3Kzaba2JHq89qP7Fa67pCJACee
cINyWHKb+8VzMGNsLsBNynWxbO5SCuBjvDIx8CVnclEuxm9HQbo4RD9+keZQ8gZg
JYNB0cFilFlJMuY6qUFcz303NCSLGohs8ChJc3O2e3bUrqWQ4if2tjr3LSaAfzqh
tVyy6+2q2XuMRjyLwOiNayV/DoMdrKINVtoOPbOH5WcTvC+tW7dpBUAQx74KJtsz
T/7lysDBFfAmsQvpklUe4Juo1GwpJ5HuJnFlXu0k5cb1bXM3QBudA4upjufn3OaE
7dyqNTmMcwOxWdr3VyxkQGWNk8+1HDYu1dDq5QFr48G0l0bItIJOM0VtN2e2+1WO
j/fkVEIgEb4B2/2rK0KSmk7vylhWyaw/lSuyL4FwGILuiuQeYpI2BkVKX4cQzOFb
GecKCszt0ir6fuABHhAvicVVJ87wawmbappr6vyaQlhXi709GU25CWZOh1WiQjvh
52Ca3IqV7kLFpMJHKBf+ADINCvTi2MLiL36cxzYnS8Vu4W9/sK4Pd2yTBY3dIvlY
sn7/jptJyHME4TvQz7+rU9sqPVKZFk3MsZoXM/Z94nJE6IP3APnWigSyqttJ5Ex7
5xuzGD/Sh+e40/vNVZwV/5vRJa5GV8aP1gwm+3pAaN5YLnyjVLl8Whw7E4raqVKV
rqCuPoDZqwmUjSnJE3UmZIjRnQG19JMXxj6OVtH6YPY2u4LOGBvCr9/O5mppwMq8
Qu2XRDb9cc19PQ0zYM8Q5qDhnN9cys0Wwz5xUSj3qvmT711W3eCvkZFkqlHvGImM
T30ZpiQEyz9rurFGqhv4ljO0IUMJy80fZcfGKJpB9b456ZKbjJsiSE/vjzbK82Jo
NaRJO/d46Ay2BHf5icyx/lMBaBzI/96frPqV6ca0S2DRFyOw1VsUS6EWA20b+NaM
4nfrXSsbt84gsk6DeCl87FgaQrmz913HEwLKE4mGuvoSRKe+9YOWtkuGTfzIquGo
Y2wdYKreCaw5TI5yDc73G6otp2LA0bn+7rtttnDLLlfs3+HSmptpRPZ1L1p0TrpO
EFOJyMsS2tpFvZ8r3YfLnIIhgGjeYVjLIbmQVlX9uiChTWo1h66sxJ2wcfK0qq+g
eUnqmALxMZDynwPHQxCbRTSAcmBRmjOT/i3ORW9g77sQb5SXsDebh7a0wjSf0/XT
/t4MeEplOp2cht8AWtbZpsRasJkDllAbEAs1p6BTdrG8wSMnOFDoHkxi6cyXrEdq
uU02rOIYWueZYiWm30NRLaDgMoRkg1WyKO4qdJQqER+BdjuPrL5GIBWPAxbYFIoI
13numLZnDjYgFw+zMMLjAzFrP6wgE5iecJxIPQoJEK2n1kYfAWoeewH8xPNwE3Cs
gqgvv8nbUOL7XifxMw7TFFINFuypNyETEV6XVrzc8jjZg7C66q3L26/48vwFBWlw
hxoFfHGZv/fo5jNTx6u82Miy+Kc9IRAOKuGuodR8n7Um9jR6/bQlcVhrbykG2XZR
MvnF4gtO+wz5Htd7uaw5t5uQOO4Mu5B18fPW9yW9YocZP7ENaAHZHXL9rNoHaIXF
LBqEe0c7/uhAPBdE17JKqydaKgj4cDixlP4nmA9QScypYt2a3Oo+AlpqhEtwQAAE
Ja/RX4DqGxmBw/fJ/6WuyFHqk3PVl7VoX9kXQYbMgOo74j7y6SkdX+nEB+tDuFAx
3JCx6Gli61SlpJ+e1Sb4SMDOihbQtGdwk/l6KK6lGXdYQA3XsjebJYnjF31PhpTC
0Fl2RcWKvSnhj4tg/fBLfjOEP4T7um+CxU0LPw3+YshfiPctn2QigbM9QhWlS1rE
sO/mtyp80kuJhVY4SppcMGeagNlS3yt44QeE+B/f3Iusy64JvLbDKzabjtZvQ7wP
4X0qhFrzYlV1cxB/+8BJk9MExqam3v44KYcMClWaL0ffUKQVVo+h4VWchFEE4QRM
PURBcD2Dx6+HBKo0Uz3Me7IsDublBOPJrO87VaatGU8frh9BAKLQf/dWTctLJa6c
dtQtpUaRoox026vQsDi1LB9DAXKgm9WhIJdKLzUMNIdVKifKaKlPd6AhyDvi5q0z
Dddje+Y3Uw6HQXqkTB90m/KJY0nvJetbT/q2pHy03vqQ2zYrnT4dJz8OG/VFMMwA
rNzy2F2umhjc16kjNbsmxdS/25UlmEniv5cxfn+Lk8yXtcISSKmTvMfQ8hgE4uQH
wpvO9fhF9mKLv5RP2gxJvKBRP0haILuludPUkyrC5f7WwSY8VwUhKE02aE/kCy0t
ndxGA7ozmYqxqX/BQ7isMA9y8aRNGnCnHypUpfduR90+v5wk1/sMo2jRwalwWpcc
e0wtFrrn0uZx477Guy7wDsJEiwL8qqxwF/CY9aN1fXT/3YzDjc2WBasaF3uyg8P/
koTitnaQgqltCEpnnq3n7hjVgJrtP6V0QzfbB5hggt+Im0MJUXBnID0rv9muyvs/
nkj1Uc1JkansSTvZVEyRV9X4eO/3HOcP1O29o+40oraMgmxPvHGSAZAfRcL0imHs
oJqGJjqUCKgqxVH0wCEVGUJi+HoZcncfqi19QFaV+GiolQTAMxocwXfBIHRIr3Pd
bu2O8jsa/rimSj5fosv33fOYLNB9XbJxKIDTx9V6Hb64InY2gWZNDT3Yr3ubX142
/HFhKZngD3AGYIw0qYo7yHnPETKZS55Q1kACn3ORS8i90vdDUhIZDuBwnekJUJkM
KFt+1b2xUbLNsN0Wo2gCPUYOZzbfCDMvDbnevUUh3BjTR7i1hdNPHOiqvNXx2Yjv
O/6Pvx9udVHUOQN41yde6Wsy0ZeIRow1qBPrnDRu7PurdfHVv3cftWKT/IX0ORlN
Tf3HRl6qfs8/bhhg5ejDHVRoacrWpGOQwuT6Za5lLXAnGHXtuzhSPHGvj+64i5lm
r1Vw50J+Wv52+UeaqhTS+QSmWPrtfiizKwvJbJEve1kjRZP+uZ7AVYPIX2Z05W4L
5aN4XtPbJWsuafzJCVWA7DAzPK9l5u2/jwZEVEugDr0gUPL5nIxOJ6G2Ey/iWN0U
bMFXAKhVCWvbt50/YbBoBJgC3seTiQTsOY4mhsGL0dqDddT+XC/YgHdbnvdq/bA+
toJd/sAFVYU6DK+wxp+2q8iBfvVVrkFfgjOnqBACkIvHi8aoBq/7QPD0R2C5xWwS
xjUKIZGh1fHMl2lxBijeKHGcPHA8z0NzAVYnOiwzs/halBtuIlDKXIL/3iTFPIeO
YCvwb6tY464UnzYa3iTcW2G9Hqyd7ZYUsvxmglZ9Y/FyRFl6yPOK7JDcmu4r7HrU
JLVaRvLWUuibgZFwCFKCqlKHabVYGGwgcLFCTIWoVZFDAJCMh/6VyzmWWBAajY5f
Rizk1CCGUoVLLqbmOYXjGKC+RYxoL+9lPHi48qRULjyhQ+0PgI3gDEN3dO2kNFHw
+PhQaW9BreiZTeNPEtg9lkjA6TxRjnGYeNLFy0+NazRbhNzJu1WV0DTId/tUFW8x
0gqwW7S5q3KBLG3xEyNXYJ5kdZTcbEm3aP3tY+3S1lO8pfzJTjmmworztt/e2dB5
q5LZLuRkrO5Th5+0JNMfknUKs9yAXgjUnXuQ4lAeOoUMCW/AKz9yRhwqEPpLDOx4
dYmEnaA30FtY0Tl5LUBLPZrGaLpYeh9UbInrVkYhZVpZJMCHYqnoSOM2QMpBVY30
+TYmWja4jG3KmH5gS0jumseIIunsHG3Xx58/KswZLibff6buITHQSd8+sCXlM0eM
5k8Qb+CQJQPsbAf3nLgGMGbdjvoGCGvC/exvheSs/QNJTW/vHbVVG5GzYFT/VQRd
97PWmTzl9Ko1Lz6LnwAbYmhfKoU3/YnCkkfO8lZoVqFgAM2D4AqY9/eC+IfD1HR4
LenRv1V85ppMHY6EnJQVqbLWbSOi0J8GH+trB+oozKPf/SYKMYPqYXv7fFHylVFQ
OEvy02tb0D81EXRCJk8TruNWk9lGG+TQrdkLzVeEopf1VkE+HPTN8I8ky/jDU/5U
N0OYySVTysbGQUZqnoZNAIN2w7xuPDuc1K+fvogIYq9E8OgqdVb1za9kjdM+NJtY
4Pz6ZkM0m3W7B6J3OLDt8u7yjW0jgmUmXVu9X1Vpy1AsntroeKwh04xU7SZ1xeFR
3FHwjdr1B4wjXv5o2PPsBlPMJ/0YK74yz86c/C+2YLjNc8CmK5SqHGsAl5BG5jtF
9ZgBrMzRudtKMF+Bo4aHuzeybo3jB7WSxo+W+6qoG9AWLYgaRdQa9QdbCJPy/ssv
PwKv3iMIPZYAfs7K4ej/yvyyN+nXCSweSjkVt11svkmePAIT6msLSdXJu5Nu+p2d
XY8di5kbc36PrxZMbMXBegUV3RNamaiVrzp2bAFZm1AQpzaNbNbNn3K1rZ38oTJP
IeZ1BlO5KBLiwQYgjSVes2mRmwGuJihtijzMmy6KmTNMT5CaUhi8xAwspKe/KfsI
Vm6JxTDJ1uKmR2ythaQrBv29JcRvIZbkqt7GeNHEyLLtdqR+zqjKQDzr+WOsJUq0
STOcqeB9HD5fkNs0Y2imDL7qYk80F8XWLIVTaVj1MDLvpesNnJziCbsnMy3ptzXf
bQSoAKVF3RkzfMJw1jB+RsurhcNd9TCexrA11aCNRMITFNAgGgp3+Qi3HlwlHgT+
a5FyJL8zwj66kaBhsJN17JZq602LSunhKRbUaF9nkpdDXNjGYkiaYZ/xUcd1cFWr
8P1rSkV3S72NL6jy7BSxd7SKtIEfg8DBjJK2668UeDAatScppGsea/K1Y43/LVeM
Ewhs6nS5S0WZTMksO/SA/XS+qqAvpTQ6uatnraeN5VWpLuEaY8jRMDsDPK7Bmy75
Gxs2yJs2lgG5kXzKjSh1152iOHLTfM1pCkvbdLoKP2VCJD8yBCGf0B5mg5nj8liw
thd1vTijKVpKhMFvxLjvjrjQd3vbZxeFWWieRSvSyGK+wLBtNgIuGQgQwxfjtVp2
QF5JV7L4Gu9Gh/aAfdbiUjOQ2im09AAlYl4Nr/yoU7qL+u6/MsxV9oCYeJsgj2GR
11MqPHBBYtSCpgqQop8elHAnlxMdQlqdhCVOrCd+KfeuhlpIkMVa4XW7tQFjIiS1
KoTP1Vqvnk1tSaq0m8QbFxaz4TLSUBoXrY/fSi2FDH2ukIrXacNCLIpF6N2gbwQE
BXp72D9CmhxnFX4BTp3OGfJcVY/tnIVThS+4lHC1LZ55vLg90+8VeKBikoZjc6P4
xmyyEXkmtfH33kOc5r1SnJ/JO1+6kZ6MWqOlB7cAGnlCXvP/wbFf3tYlkRm80E4U
N9qtxzXDvNE3B9rKaEvELBGX/EQVMqT8n6BShAbmNaNohM5F3+0bT325qajU35Ng
zjydehFA7684Y8vfqP0bk3sIV+wCg0Jf9XZMdLrXbUsmY4CYwprMYMOhzNipfCoq
3pCfSqo7IgnPOBfkP3AWr8/eUdwzEtp29BlrsdZqhrdcEsxiB7vnvaGuP2NvE81o
0uszzQwT4lhxGs9qnSR/3iq35q5oFb91E1PJTChOpR83ekJnYzAI4vl9e/8K0IYq
XkxTx2+sEPBuA/b1apNzStbugltlTpNjc4ImeXlKGVUR0h5n/1xYRNeY33Mc5xvT
T8OC50iO+MXJ4D0D0TuEJLX4JVkG3V1Z1p8g+ZFpA6+qwINcG7yQpKfsHyIDNWO0
gSwCO9fyGu291L47YmCH41BKozqHDKhXMPNm0gixKUxa5Afoh7UmB8NiXSh23LNP
+dNlS7xUZ7hJcZphSF+ON8m8b3boSGDURkrcauaGwZnZZQpLpWL4UlVoFU8KQD2Q
020vOAt0El3s8XjjFr+k9UFuWYKVg73BnfjXEPZYe1jBsb9ra14TUX8S4+wJDZ/M
KH1HRQuBbZw6IcCPWha9AuCYTBotkNuGezL974qd0sISqA3AkKRm4LItbp9A7bqY
1NDC/VAZX1cFjAs5ogbyEGtEodm7Irgi1LQW+LKPZZOjTUlSjmovv7snjyZSFU+Y
d38VteLcCzgFJGGN2o3YYJl/TICZ80Z+9jL33xWRL18wao9CgVXyoNyjzihN5Ird
UeLO9Sn7xHG/DjoMuOXBeUOKx35JpM75dM+u+rLA1bSVnykmhifbPJUV/2OVce2Q
ZuiZ8yNQgSYuqeVTuwNASeVDKe8vZe6b6BXlAnmY8DPg0ril4QxsMBObtPyWrb6O
wZdb+5tBGEnkj1ZkHywtoCuY9cO8QZ7yt22rQPR/FsyxXcoa0m/BpIFLiAhD/YrS
KbzRkLWK5xTiq48DttfsUIsw38Ftn8av2+wVwEsD08oSQvL1FddErWOY7NEafBFy
O21gmht5WMDr8Mx/Gx2Z5PRWWYKBTyWUGPWTaHAZ4Gkm0uFvELJiDf9b/6QZ3gsu
Rapo8MmKnmRZ2uYfJguJJ3mJ7nfPojLH533ibRZG/Ml2mtChGgudNBLqRmlpCRl2
ZxsIESNGhvwYtgrhPWPikObzvouROYtWWh8vDzw/8UPPkFib9rgiI7NCQ/2vmndF
5E0OMwCai0rnItBrUFIUs45jEEXVafkTGYJdoPvoKXYAC1U8Un9ONVN5/cflaCJ+
9rXoEyW1Q39uG1S8sNc563jnuxrrNF7S7ZLkHZ1LhE7T623aHvTTOpeUKKZ2D72C
bC0z/MxkdhlQSMvuhSLiDjjWu9dELcwYBw7qDme/Ar9r0PbcWPX+K8fvVhAACE4x
mTFaBrrNbjBAr9NzLqrkSEhYlvFGPHj60KWl9QqRp3AbF8mL76VdfhTRB3rb4q7J
wRR6sNwb3JA8Dyy1S4uhsuYp+OStes6/02vnYbb1BNa7vRA6uvEBEGMRms2eb1Ee
fdnzm3hgkSATG3bOIZQwF+QkRw+lvIkzI8nY4FhTPxZR8lp//CvjA6fq6l3yG+uM
UqizRQrpcHcgIRG1IfKTCK2zGm0bS29O7AIBBExYOqvbFmg0ybupYotnC3JACErv
u1MSP92qCs4DNw9EKE1Dlr5+huzUBUWMCe/OmeQ9ARLMQur3yg3nhsHuymmakqzH
t778MLBrS+R59njZy+nGXiUQeIQ/Ys9bL6sBsGIp7fG4IgaQGvbjrL9vqxYG2srj
OvshhBl9DEI+0o4X3T4eui0g8HX5dBTKaki9tJz7LuK10iiWryqDEEHtr5H6C596
+EX8h/bimq/Bugk+cb7iUqQVFyCmxzRbypearbcCRfqg9ywFTxi/By5TmDc/iD2w
2VEzVqfmb0OTNchXPOoZ8ThXB1eV5nacKwZm30k6jllHUE8b03xfVpZcYndwNqbz
DzyOoNZl3UcCgy+3g6l2NDgK8fj6GcBHknZ4mgHRF9NSiTwDXARSDIXvRnQCRhZM
NKrOqNPJ5ZxIu/d688PW7lJ0nmL5SUpGNMqZj1krhd9hMSbDDb9bHdVzIZBTQj/l
kHogKyzZwRIq0nBOnDm6TPaMMo1yRTjqYjvCTrPGIIZMhz8ECsVbX+cBsdogAHSc
r/xbEuFZy3VtrtDiFcTcbRAKHu1M24b1Dc9xBlW9P/YpvGsMSLVPJrJeLalAmGt7
rG/2inwxG5ZT75FhPkPdP1uvDQ4TS+c6Il2btN65u6YgkF7YrG2g82So5a4C93HE
hTFY/Axp12HKyB2P/tB7hB8I0Oj0n5SABiuq3eDNsBzPfq+Anoxd1zIjMk7JS4H8
lBRXeHrTGewjhnWGZjKWPlgvU7HKo/HZwbqVKvhSEsHk3OEk9PBcwET+8Fu4KmKh
6LhYnEXZOJ/Agsu7oOVaxypbGAppF/RkEuaUJREv61FrM57+o61l7XqkcF8Bd19Y
6ofv5q3tnYWdoh6p+jaKMldzmwJtZzRTXx210PLPXOm30Og+jOC3+tXcLG0YBvdk
3h3OVt5NDwReguoZSSpA7sLGs3N1FiPMyADShAi909lhR2ozdHP5IouCUREAXzEE
0OXcfg2riZeK0YGLOHybUn3f4eLwCj9lNZggdOuBCuNzS9agn8r7BiSfknciTe3Y
ulmsCrPc1Kb3ZkqFGY5q5Mt+ulZBm4cVgmQjZB2+bsxmYaUWSJPZD6jElL2r/oOf
wJuBO+jHyVutRcp87RAjAP5/VV0zPGJFaJgPDZocnFLWoUodA5sylF2h+TbIr2vS
8pdFLitpCadwzmSHp6nJZ9WHV7d9/1whUL5WBzN01QPyepEHSrno7gb4pXChcjmQ
PDSbty1pFDsSj4uRdtZC4wfc0NIiTxpO+mcUe8XqCjOBgc8LbdAA9/wu+KiWPfGA
DhZYn1eeWZYirUVJXCsplJ7MYBI+Qwl5ZiXO8UBwUrcOUD3X4lrRybjLGxNgR01x
IbKePmmBMP+oqH90NBPTQGop+kMBO14LQgzug8ksnGS7iiYKCwvd7bTU2mniMD0W
NEtdT0HJ6u8DGGnrSFB10PymTeu97xx1K3/Hbj5WySRK0aQRZoreJ4lb2YPMzZ3U
cfYWtgIOAdIUH/uRFuqUIJooFT3bPAafYhb2c2Fp4HSlcP2fn9gupdV2fk0dlrTP
cFZO9hnaLK9fn+fRNAPEO5MWThWyg0HaYMIFuIkv1yl338vJdYIOtEdV4EG+0BNE
0fnagh9D4/2LqfeHSDfaqetpKrcCFbaObD1yF34+Wwj+KGX+u/1xtm7gq6qqbi/d
IBx6wgmPRNDURewHxdLOeoFtDrjRzsSCXM4hPd3Nk9iDZnJVjV4NPTzt4k32Jh/r
tO246JI1+cQPGpvb9pQagY/qS78k/Y3G8NY8CbEZr+586x2uwEAbSSTl2Egu1UI1
2N7L/xl/eyIYxWwV8tZTsZprBG/yKGMScsFtc99oELVvSNhGEFgEC43BOvGDqlbx
o/d3DpxrSrBvWCUziwEkMq9cRBcWXfeJXiBRPyMzC7qFGGsXlpzqP4XwIbZza4ox
34hejIuYZAa6H6po5gLgZBjqiNAc0i8K3oX8EzU0keVnQ2DbLmBsrjGox0aIiqbT
tuxfKNUZ4zPBAlo3A7VvYJ6b15AY8z49BOEUr9iCGAXFD5xC6iQMYnlTPVkDDFPG
R0ZTBGauj6Lwnll/wym4UqZ4sOt2E+5pIckLA4yoFTQ9RrcQhaWttAS/7QCY1v5m
1ZwhGJYR4cK6WAlpPLNQp8QbW16raaUImjI2rVHZ3tkKnba9LJBMpMj8vQGDnrCW
uPeHXfpLGSCR/jLyWmFJWs2zbvDu4tOPFmUYdgClCm+U7MFglIJpY/4wMVzJbFhA
/ae32FD9kGM5BE4KI/Ha7Ik454fJunZFfw3RTBJnrHjDGUrndUQrbxJxr1Dr2n5E
3AbizFqIBXjFlqLvpsPlJe9mu00gWZmR3dv8dFrMtRzr+pcuklBIyU+lWUfKQFzP
CcHmaJdQOxYxe6oTTgXS+KhIumB/2BTIO2j16Sr623ZGzHR98ZIYSFThu5jWH7IG
h3a03ieYpbfbRaU3OXe1lI4QnPD3HNJVf8qCaIdW4iBLczJ/TLl6Kd6zWK7AQBNV
a0e22nKhNUTvjUHQJ/0v6b7WaeqMeM4TTNg8dwJ6BJcV3jgFjk2OQFMWLh+6WWK0
GzOnh7BdtMTn7JeO4PqH39/Ap3zzzN0w799S4TX6YVlwoPG0XO9RDk9yZP3A31GQ
p1r/uG0mSYQtSwIl1BtvZpCkcnQ7VsU2KC30jtg+U9vELtDcfCezOSMjkQIY7UuH
kn56OVv+pX1cSE52icUo4MP5fWb/v6EowJn5qAixaeLoIKWL6OqdrqTdN3O1FKLX
EakRuDPQDzWeETvtL27DF8upfMgf3yWbTWnb9XQNAXKzz+pRNYGByFZ01tMFU2H1
KwHsOn8pSha1nwS1uYrYgPc+H246+O9sZhEYUFqomi/wz0N2TDL6r7uGavhvTy7X
9O2NDV+ElHaNRs0xC5uf3mWbbrLZ3Or7jEmQcp0+oEpB+N1KjWA4VStRT42rybZu
kZpby1FGbIfx1kagduhK3FPm3GLSRieg/qds94v6eMCQUxREjEZKHcyHQWzYnRVY
/PUT7oajjf3GgdddUQPVFEVmV8HugA5oB9rcp3ykQMlWbdYdfBSxyiu5EX8Y0ngl
CD0liD/+9EJBK2PTde8PR7JyKCpXlu1AtOuLLUw0JU/4387UrPMrICfsLXHAwIF4
thy+384sMfe4wo6zTjAMf4fwPdo4Gvr7t35Ktz4ogRwpFNs3duuQGEZ4mH6uk3Zs
PigVmwJXhfCY2zoncYN/mFpnMh4bzvka4hgcTfcTRvXhfCF2deh5+BFexRtoS9Zg
jPeORWUj5w9JiwaO6m4g7G7DRJj3E+is1mMUDv6A/FsJ9kIWKbiRX5N1HISFtijO
1Mopm3fpm3y/Lp2th8NiKwCFYAf3LNErVHS+CafH2HaqQbowDNCFOKzZOcgn6gat
qV1BRVe+sK/ihvHlWg0DxZKyRPa/qegFAnzu7k9CUSOiw1HdGXOlPfEZ2hm9b1dl
Qc9YiV01ajJpi08LyiB7lHBCAFGfNiqjXzXMV4UaH944nZh0VpvNt5AbAQc85GXz
Dhl6sVXzCKHnsNSx+dHI6PNs7tXp6+3+xz92ISzv3FMV1pubQro/1fCUHEnfg1lD
JonZ42lV146zqSijmOi1p34EbyCQxHrDCdMVhOtzNN+5KBUHIkfl1+i8f/sbSPUg
UrANll1zCY6OBZXueFtxmXeV+Pcg0DYIfaFaAdptp4dDy47Q9oLA3xndoaivzTr7
RQsDgCvtsrrOt01t1MyhOviW75UxeYXLkpha1c3jez7uuBR6eEvlFy7QCpZzaVUk
fBjNhwqp0REKpIHEZlPwqJyOs/AJqIR+TpsjZXdfjDHIbtMRyEqLjAxZcBl6Xwft
vNacETffzfbAPUIQuH5pEX/rlAmEqSZdzVkPCxxYkSOa6zfSguc5jDYsY/d68QsQ
07aRT6ug1UWxX0p5Ln/cASjL+pJnZKeS6UQTgrZJ+ZmJEQscPcbPOYdjWYoneNgr
Hg53C07W9tJKBP0sh47AtDsvrgXykmUN/VQxG35YOKjnEkQbo3XW87bz+k8ymcUR
jiX747MFxNmZgXgXK/02vSvTrqw5Ym4YIi3AsHSRUqWnOzcepLFL30BA7YClauBd
5xFu3iZFhw2Zd7fU7XEQly+K3isiXPsbue7j4zZQ8gBB5Xa09PubgT63TGMvp+k7
9+MqP4qgb4IduQIi3qkBAs75PX5HPtPS9hZSHkNEjnXWs+lRZo3OdCzcizMNzJDY
Rc+TZX+mwJQJdgAayHymEC2OhKh8xr0UJHs+Swmg7oGJ3sMcsWNup8/cSREG5KrY
KOEh6r6KQfl3sFT41TIDIVQOK2SOnPPLYN4+8/73E2MNLUgH3R8rEg/xk63QVL6g
D8vKNw8XjYAyaDH9iw88BkrVqEdg5nv22rH9brqFeW32GyxLrVn9ht0QrMGmRmnZ
C9O4TwIHZeVM0uimQXVjRzQ8tr3Vryl2ilNhlHhGvypjfZwjp/KxU1eB6frl7E7k
nNPjPcOohLHqWizIokmSwvqZcZYkVqw2qqmN1rKqf0irbmHsVgWrU2cXVxFPhdHm
e3ElK+YVTSG10A+0POh/hS4TMYZa2j7HgWEEnbM82mTvAGLwo3G9q0VOlnfeuZ9E
LEBdCnbrNgo8VAeAMPF51jn0VIzmsyaKC3ZsQT5Y2dYg6T3j7zM9f+BSbWE80RCg
pGcBLKph0Upz8yM0Zw1C4uijxfsdqWquwInj2CbHuiqeJ/75rtyTMwa0DbjBf7jk
1+BlYQvBkGJP+3GcQ12tLA4bigkt6W3FpVJZAHc1rL868S/ZY15DOsA0V8wGcfFf
6grdJlqn0feT9uDSIBp4eyO/DWzxQtchrxsqjWBL06NlJKQFMz7EElS1TycLFDpG
nyVu2N1hyqqi/iDBl6Y7ohNutQgex7G4fJEX7CNhqX9TJKKiD8ZoSKLrvsI3EAK3
yUAeXgXZsYY5J3cAlo4bjKtioBS8LCqRsRvVMajcgb4dlpMZ1RFvpNvSauqLduaD
Iq08YX8k2mUYRCDFTPO8b2EmNgvuoQzFzLiN5nibYxGGshg2xyfjE/Jqg8aDfKDy
EVPiD1oWxsVKAzG7OwyiYsGTUEAtjGxuGDec7a5w9T8hQrg+wO+dPPPX6PvfPtTi
mgJfFpxpFs62J3Gptdwop1lY+IhhNOt0nq7wWw0fkniEu5qGxOxz5YdUw+C6zvPr
rQ1hsZyq2QaPlf6VGl86uMCkdwriaMmmfQPi/OBXxwfX2qoUriCPBqtCG8zjg9yb
AO2qoBaQS5iIr/vp0CcFGD1zJTBjjjZbFf4LVUxwfjPci2BsSV9EG4nbaMeXXAYH
qGLIFvXl9MjIbZS+BDL5b8BDlSOYVHqt4ZCBrgn7exf6a/vBrZD9l3n2BQzV9WUa
0iKytSv4tOP6kq5cDCmFiEWOSKtJF1U/Xg6Q+80sgxi7ITeSpx+hZkpjg5iojPok
RCZo1dUjxuY+L6Ee/0rOrpUUBIvVvBiICBVPlnYuhMJ/luLhFOxvlTGYVHwQ5sk9
QkXqi6xCPRc7/+QwoWrteBaxlfnDtoNKWM4KyCEKaNT0unhYYrnc2VgIrBrdBasj
C3xpxyTZwO1Ta+G0OeY5jCFn7PC6Cn9yRs5I5+7QDMUC9IAcwlq5eEhFH/76xz04
sooM13XGjzkjTDIcD9ubp756vKqsef2UdjE39MFIfC/rS04F8G/L2ZKtQTCPA4N6
VeqM7KqGpPaClfstHivsV+H20qtC+0h9zvwBjWMQqFIgSc2HdziWyZ8Nw8IiaXBk
LcfykwTy0UNXY0OJlhqQ+Qfb4nAcy8KnjTBZJ91cwYa1Hlzrow7C8Ak7gi5qImF/
jENRMJdWMJB3XqfuVbtfritJHfFt9exhahta6pa97KAJ9dS+jW08lq8xv8RYXUou
5lt+yQw0J0I5fJ/Ra11fjSKcF5U+RGIMfKwjEW10J2Hy+grNME3YRktUu9WE0GJ4
Xpf+x88EEImWahoh/wnEVTrqK5cDxMHiWWalt3qTHVWIF7JUoB1K66JxarG+II1J
axJspMePDLA8Iw4Qh/FhPb32h/he69ZKIkWJrne14DLAj8sDoxYlN++TsLUH3sg3
NxANELmx37JKgu3Xn3rc+tsHco53asBoivwRaYI7UFb1yTucfMQtDGUwyInCPjnG
G/gI8NjDja4xnORmN1eOzbFMBBSGbhy0OOOUGplkaII3NWCzMrHmhHLbjF8XAsxp
49ECL6SS5PzCljr2dgwoOjuOl/a6trdnhPYH0fTzA9hn/5+XvNUZKvt99qbr/Ybt
q36q5CYNBsMAJ+W4R8v+zANitiAP8kKnMr2xKlcDmf30+ts7f9idrJdtbRmYmZ8b
CuD4Q2Kx9CYxLz6ChTmv8zV3/5uhwckIm/Vvezf5jaeyljk/k7bg/I5QzbFRksDG
cyJEO5jBPxK5pWSApfhCnvvWeZIG7TIKoLlmmoJ/Blqia6xNXqLX4qocymS8CSQt
7Zrh8QjL8jL4gDn9eyJLUbmlapdflwuUJKSVPGVWzGdIQiEe6kVLRrvs++cFGnwn
GjdAcCOFvscBEgqgi3h56zfAixmzu0pdl9spLJGBVsxw3pMeRjQLrEZLAPHSMzTq
6jPTUIWEMmJWhJXw2lizoF54c96A0DxDp3TBHyuhhjP5bmh3bigceh3RFIOQhSy9
Irrx/e3DlqbgI4/6B+H39uO8OPckbGyruRNPEPYwwpXigRNg67xdIkx0dkJjDYLa
Ga8bt0EK5iLygnuY7ahRTyjGT3xYAmX/VFSS1IbsKfe8bk2cgbQH9hYeRTlNgptx
FAJTmLC3nlUpgpxJoQmik8kagkcmBxDW/1bWhDjTUvDCQ19+Q9P4YmIMBq9AX0I6
7A+HBoyLjKh4hXdg5FS9c6SJOO00OisfDg7o0TDN9el7Kjx0gGn4PacTVGfXsUeI
B2y70nrzxmCqE3ptwuWn+wxCYQFseoRP2fKO9xBOv4Xbp4ct/AO9YUa5WmACAsTe
VOWKVdUJVYku7W5uIFccXwt7b58SToBV4Yn0nZux48XvLuw5z3NP7A1o7H5mZh86
OkSYSSrz3zZJDWZqbhoyAOxErwPBuIv+n44Xi4EXkvHZvuemZmwYRyjOnCIAAi3t
mG8V6cjlfag1/5X1Qeh4oCJu9fOVhzocio4EyNcr/D+AKTHU2leH7BwzSlaAYTEt
3MpncINc0NecJ5UBqeE8CIYf/kmWaR33dEp4Srt+mB63ILSzXA+1MQSI6A8BY5Jz
Ynm+qyHdUgeJ91Y1MLE8WhAUK1BdcEnH8f1zd7X8vVbUy0CqhOxtUCRUalU8OSrP
7mKZKYpDYQUJJjssEH7B/DyGUVcQj0hlYh8UgLTi4E7FnxwmiEH7Itq7aApf2b0r
PFFWb77DqJ7cIFZsZPiI4MvkHJK9TLGDpIEVHmKT6OletpR3xK3EkKtPw4bG+Hqy
Jojb994cakEolvJAA6WiiXdXUekWtqM+jTR3iYnngrZP7Q4kkqtDNIQGdqn8WAn5
slijj9Y/M4XRfNYKXM0bfPyC2v+B6zkMkjr46hFTorNnoRvssrnewkjdi9YifKQj
6sGMF8sBqmL7+Mx1PcKYRIiKqHpEDwfvZdxakwN9lYx0onuiODGMaXFRxqEXycPZ
Fw7kEyb1bFBD+zPBq5yDyarERvavrQdeqzAPIE+jDtZqUxdn9VGa9P9h90WPK8xC
iksLbQRo8aNQnMju5JJGEzBl4xViWksEYgjgIq2m/Ligs5fNZa5el2FSAQe+nXk3
9eMytsgI+ZGPgsD77DHaKyeU+gBZ771Z50VfgnaMMzN8D/PYPjmhat8v4M2eCT04
68hbeQHwDS/mBG8oLw1Emfu2pl/KroOz3kHhT7hFZWDrYMSZt4ENZwfLPiRRacrt
sDpWJ4XSVQ9JZR3KX+EOgkq8OJqouneYHV6JV4n0i1eMRrIDQi/kkMlZmfAa+JfA
TB5kPrqe4cAtZoWqEj3Sz4M5qWjBPvC4qWFejDeAyBdgMEjNq+F7Avk3M0bb0MLw
SaM94ndV/SjYbI44PrD+a88z8tmdTDQfMy0g1v9XZwkBbb2vkG33nTQJFXQjLDtz
nwMSvSx6gExmq0GjBXvF9eJF6rCYLyebkEiOLFqLHo8ixDWhEo1ynhipgwPOtoOI
h13sW9PLpni6n3g1i8mtLo65beAHDbAkAAnLcu8pZcHGYBXmhkemyOdR3GOdgSUt
4O4lvkxmYrwdc3xBsuy2S4lm6JuZIMgGKfKJ918UDtbDz7+GVb7PnP/TepOZBiec
cQ1qb/7kIHWyCUSKAVsos9oH/q1aYIFFaUKjWxb5r6/oJV48WPlLA1dNqFruaPrt
VyvP7xkWzGQ3u4fCShr48ueC6guQLtX32M7FBL06Bq0lb68t5NxXa9IuVhlcvXFM
NTK5PkAVHG2Fe051jOf9p8gLSZvCWxjoLCYtGoIrVaW45v8KLdXW0UzmCOUEeH6y
TF06oQKv77+yKlV9BqJZ3NQKGdbjSijDvtZkBwg+erVZuzX9QSaNgTJPVL0eNfuq
5AITRvZ/joWvI3kFyQncD+dLYxVImCtgxJy/uzf/FbXadP3VtmIO8X4i7sGyT+fS
XY9ebR1lY69Ctep7pAyF7tDeAq8wu1jCAkNKDu75SStVPWTyrXCGQPnvHomtsarA
wh+W43fkc88ual7NjS+ltWPku3wRx8UntJd2LA2j54FXetUsTYfvw827UljKFeKW
jKLVtoZ+k3/ITQCIT84EQNCdtEmUA6BJyah2h6AaLJjPUxNmJtODtn+fvrJBC5zW
5Gno4yDgLVxcCshb1qTfyln7Zq6y+VgLsS295Z7imU5M9V26vP3WA21lR0EywUhi
vRIVRgANV/DkT/+FpXS6GtLUbIJNhtfBIvbBEdQE7FW5Wi1KRq1FCVdoYqpGWHna
K9Tfb1hfyQLPN5O9GNBa8NcjVcTuh+12PPyxe+l/0w3w+hohZ5kQxnaVdszHHwlX
AGYdAhb3imd3ixLT13lxd82eumg+VxunoIhS6aJ9VSIN5T1+q4j8TiBvTj1Er7Ld
iFmTGCnMTXJqnhcpXlx2kHbK2onj3MRToDQBYYtxTF1/izu8ExrjtuoMZAxUeNWT
GNq8j1wOThMPGb9B9MR806JOlD735VGCOXXo9BBhTpJC+u/COd3phAPArZcNdGZg
eFpRGAGsxNHhGnbC3FbbTUqd+gsfsAfqq4uoff0UHOza5UuP2ZkwunN++L2YvyAe
pcGmaE8ePdM3xlZMZmK3zlSQCU5f5rDJnOjvP8F/65Cr6LzaoXXE02ETWfLOwvJx
OEiWXME33uQGN0YWPHwsvVMbpnEGfO/RPbgeDXjE0EIGZ9q0GGXRjndOMu1y2072
RDQBMKtc9R3dvXVND90kFvV338hngqf1D/GXXMjsyjPPKIhRWKY+VfClSr+VBpan
QCzSdjrGuqmPjkSVSaf+5IdahlPWC6Xjx8pcH5Nkz42O3lDvwnxCTjKm8YNfeSy7
SDObfgfQATr8AxLK+iuquxn9tQ3s7CMls7J2+GahGsuoPXD/1zA9oxxviUqdPVDM
Inq/aNDHgHjS5WkmnTRXk/b1e07J16/1fFXEs/64LPz2Jq9k6RNcMP4TFzL4vfyT
hWJBAySP0sNTXL6kO2XikTGcdPOBH4/+KoUOkKspebv2ViEnwQJ+LWBL5k11A7qy
i5fi4bybeJWAjNeF7WhoAiMn1u9ZvlzR/SbahRt9iKLVv6yRCvi3jHikT0ba1Tso
yv1THHBnd+k3loD+dWX5ea9+LfyyRWePvboOrR2FAHcKFMYblbzpw2VrYnOTV+9z
E1FAeSpG7p8WbUC2q5VZcwCjYJLFkHF0NC2PLWYsXbmVp81NkEjmL6I3deKLZMDk
8CW5DJkonDYFNTMty5VP9Kd4AaxsfuhNXaBpLaHc6mBFR6O9R8yLbJzyidWf2eaY
ZDFebhaI+/jE8clKXYVy9e69s6RIK6y+9aFwIL139a3rTbIVoKwZ2uib3ikMrw+R
Cj0ZOHsO5xaXVFAnLz9YR9M+4t/pV2Z2U1ozUDlGpAFxusmKs6aAQxa5AQjKa1RJ
WDsuOh2KM3P0Jh3wEUuzRST1sPyI0ZOxcNKDTsYAsXG5s1v09nfzgM+h8f4sXTSA
iX2R9f8PfxMvkHYuITzQ4aY/BSmhyztG7LPj0owIvgeMpS0otqrXYDIpqc+HLr/U
l3Sxy8ggpFBAhxIzHqLr3DS98n5kQz4NKg+ifvgBmic1/hc/SbKiOToqHQnXtgLd
FGgO8DbuxW+XX0u/ReGs2JwMLZNX8/1Bwz8jS3vIQZaya/oDFSaZ+mdf5cAloNWo
+d+4VUMWcYVKhFJWk9nwjP3+vPQNTvprNsb5/9Ca+P4xFMNkOxWNfHBfA8Aqu+st
4/D4BRXH5uy9xNkhLu5ZznF5ZyA63Ut/EtSU0FX6w1cKR2ZEgJaOjau5/EEFjAzZ
INTWWaullqoaJbpJPdjNJ4pXlhoG1QyX5csKZ4LhjYaNbZYD4Fgz6Xg6I4pkV2/5
kuf11AvMAnVpGBWcARfNOU4M6yWiFB1vXODFOS0/6LaAyIvr7Mnp7m8Tu0xB0vOa
CRBrVHfiwuWo/av5xzkAyWZlMMRpiWwJU47bJ5A85dviNPL24EIvE4y3BGh2zTiy
Rv772LwX6Ab5s/pqTZruQNkwXxjB5tTu6oh604X03ljIMggy1ptgwLitF3//K11h
g77TIKOkOKzqiS92ix1CPnGZptRn+r1rp8Jdur6eGng6Xxhiw5ByreUBloBGAzu9
Keg0pzdkLxuNXxgD1rPa1/ORzH3ze/NCkYwmDXNE+YiUybspS93Obv9k7O9TGESH
Mao4sxnzxbTU3LOfK8e/aDrTH/e8OFSlBXNBYNqdJ5moLvXT+X89/djelXeYxmCY
hKvUku7ObziHfrdwcjceiLBy7JhvfEA39bQpVsyX1brm7c5qDo04R4m5FAZddap/
XT3dHYOsvsOFtYJLizptJp45Jc2yRwTLV8AcqYD2HknjHUlM/O01rV8FqX47RYGo
kFQbgW994PhLhu8FaKVLq3CrwwOynv9ecKwRlm73fvR4594aGz9YlByVpzs08v8+
qViqlDpZE2b+iwjf5jFOIQZFf4u5iRTb1/p5iWnLtkx52TSPAeZmlDmfuS+smGld
IXMlRG/B7VpLKkp63+669XHDFMXelZ2GKToBMC/Bq+s33hkTY6844CBQ189S7/Ut
qvZhM0/wbZGf89TN2UOtZxUN/sb/Gak3Hdk0P2l/haABG/uRDzQXTWPspeAyoUIB
6c6stP/GterkT7ARMm96Y8SJCo/R21gwHah5Ca0Bae1YS47wq/07NHMxy45z6CYA
O43mTy6RwVm8pS3Qi0hSGjs3Ln7eEUxshaf3c/Eeu5fXazzHZ0/3GirLvlCrdLSc
fOxjc5s5c9VI9Da36n3c8rzReU8B2QNIBa/gtxe3h9Egh+MRj82jXP+3Y+nwyddz
QtxDwpezQqfSHvQEOZq6KO2hDEGHTwDP4TYj6K0pVyyKbFRcvs99UC4gOvIGLeSA
gLr0rQvdqhxn2zaFiFKh2MNl3qarw4/pEJRmKGI+dgS85jATo3gwj/iMH4LvmZSS
KK8h0KdqJ8yYQq6FhBr5aLFo1fN3f7O9Ke0S9g/us6SlSFunufHOyWdSk75f5Jvl
rjGLFfgeD/XkYiNE5lA3lJJgqSQ05k1kfCDcLRNLoHob5Kr+1hRey/7dLXWmg6QS
znSc78QA+1Mdrcp2/VU3j2pLDjk6ezzdKkVpNwPHtzlhrylcpRWRk1D8cIJcx2zM
VD9+qu//IGzYwv6Ey2hV4iCNwOoxWFq8G6EF8E4jxrl/7pekirxtoyW9HdaoApAU
j7k/W1v36YCJmcvh6/EpgwQu/Bzelgj+WAYHhlGMj4aK6/xhBH5xtDa85bP78HCJ
5IENW7bJ73E4gTML3HbPlSk3jfRxyLUWQ9Y7T4aaPjR7JE1O0QfMCa/BSWV+0Oyj
fqUP1RGmcPeSfjRGXhklfJjAyUV57qouACVvvtY2r61Dx/9mz2a/LrwMhDzvVzaC
AWRXn/gPC7tjKzxSoa2HrxEgyhN4E2RSh8aIsU+OuXrrt9/hoswy+/+esYK57RYF
+dv0mFG6bjwqk4dbsupLICm2Wdub7W2eVDICycfdQ7d5lKFRCzRgrx5iO8PPbInX
JGYWITkh4fwZ9yxUD3GmFzYO3QPLITDmLjDeJDEg4qzw3t0HDfc+zJnSbFjb6p5L
Pw6jg+LU6piYTnrCxnU82HRvWqdS/JT953YUwq3AOBg9CON0E6eOExen5N6wsUDP
5n3h+DMk2bS1BT9a4NuD3Me6zemMbo8qgDk9e3AUCu9qEyvB4waGlMYWXxuTAjf+
pjG/eg9lKDwOSBa/Y7LtaqsonKV1gsmPFGGfawEolLZfqwHP19MXMqv3VXNrT+cW
/HXI4d6c/sqNw9p082/0xNqq7wbSKkdwrsbYvEBhqfJ9Y4iHrFR5K9C91L+iXLGf
+GJ5owe7I66IKgy+HK81UnT+YYAQ1Ho9FDY9MYoyzgm/0TwKuKr/7Pn2LZqYkaIH
ATB05BmD6um/O1Duj1DG6Xa2v1Kg2slYa3u1kBob5DUKXJNwDUcO1DjjixkuBxtc
J3YHGDuKW5cwKVUEa2YuGjBsW3lF/zmKZeTQBtC6m13r7cogWAL1ul5e0s4nNfQa
RqouRYQdUkRV1FNQiz/L1w==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRb2bg4GYY85uFyF8BAKcssVxBc71DmYCaM0gimDzSZPARYSF+Wr8mF3Kt0R5TqJ
hIoHRgsHbAlh5HPHlYehjEy995SAbOy3CXy/BSs9AMkdVUr44gMaRmC1EBWzPL64
S/asShyyoVYqTf3iDn/2HVDEKAQ6vVLRDu2DcxjZLEHqzHCXjTTZJhi6zJFVI8Cm
EKma1/jGQ8Oi41uIiXwI6U9WNQ1Qea2Nrv5IHdyfomjyqz4sQNP5NCotO1BCs18b
ufTRUM6rsJ1yevvvjt0NupNC3Mj5IUDLJafvQrMsX5jem5ErcMy1o1e/huHgrXxK
Rz86G7laO6FH8W1NQ4BOg5q95E4rhFUgkI4pa78IN7+oiqQ9chkLMuiqP/JEirv9
wQnAHpdEqsiru+fuQu05DBCB3rDhDXLDLbEu4V/GF6U7ZgVwByCSTSssx+Ggo9l+
wk3FOSI6A12nO0Cm/qG8P1o93k5riVdyQEffgajGmbT58Jjpmiw8RqhiCQsxg9k2
m2nxshtOJz6KIAiCAzYV5rP1NWHy4wAJfzWnZU4/YDZWNGKBs9Ge9kgECja9zDN/
BPDyqA54/SnL9zRvY9sx8a99HwdjIAbBETMMIoxWKLax93lBuHNjbe8Bgzd+sEYe
MsSvzB5JXRrf/Vg8aaj/e7ja6mG32xaOW6sEiTK3Tr/cidXs9RTHyU213Ru8UAiu
nOULGT7swh5fuMipzLoofl9mMz3x+8zlPjOn8Zu2kKZ1gVKQCg9NarXv0z0m/CAR
jDjEoQx0PUzrxTIR1revNUsKQp/TXRhjUFEK+fpaCGtIXX+NlwCS6kOa/5pOccRx
PWpBINqRVlmkCMrk39YIyev2nyfNtXAJ30V5NUsg+xIgIYAca6KhG9gyCKspD2Br
spEFkECn/NHvXblAbCoifiCWPt+4h819ChXaPUY9WajdqASOCLyf12Noy7EqthFz
rTPz2hdWvLm6gPg9wtcZeXztBDxnZJAZI7WcR/QCHErAoq7kd0BWmvZ/ntUmO2hj
ojpiXCigiMMQBl5vBQjgYrgWDPd4HMIl2vHf5ug5n2BT9vmJ1VivGNQ5+TPlGWW6
pFbYm/Tpl2SdMt3ZtUy00s0zG7O6lig52iAN4C+gtg186mptOriv5KezY5IGmu+Z
Y2YlSKvnlHft/GHt5LXAiDMny9eUqTY6IkBhNEYx4REFvMhhdJRdMFJJgW70Ztuq
35Y6I9GyRkFtvDkqJdBEmm4q7r+4g/ziKMHhfELVJv0=
`protect END_PROTECTED

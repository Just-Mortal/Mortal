`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6LCgA2LYEma+9Mm5AL+Y2G2AaEsjQ8BsIOnwo9gYdtH2uxV9xyg2lQdARs3Y8Qy
BhQdDZ6Z46fHZ2kNkSuhaBLhczdvXnhcOOg6qe/sBDYrwk0cQ/OxDbLpO3sbqKiY
Xlf4GIVBU79UQoBxJxS0AfPFOCxKtePjv8kfRB/kvXnLPQK859dJHzEFJY78hGal
V3R/QPPoYhGwNhyQOzJQaokWi49jh37/mYLoL3tRB+UerYHrd4E+p0pHn6ywyQ9E
SeRRkNQ9cRrIhYHU6vX2GT0RqHfDdYEgCEW9cNB0b3fYAUnCbSUsGx0eTBynjGF0
3jmYmX5FXZgU14ye9W9E7DBVGplUPCzWWDumeFHDJDcZBuSzHWnMaxO5NxDllLWn
/AUT9A1T+NyfP6vFBQtoh8Axf6NHJXFvdm/sh82nt9ACm2QtfqvTQMDz41tb05PL
k6Pz0yYtTANWBnG+Nb1TPqwqdUR0d6axVTP+kZ7OreMgPl99eE2x1DAEahHDfKvb
7KKc2H584BNsdOG27MXWLqn6IUy7GXZSAgHCIcu2Sj1mjQU+5XPmf+JUkvfPVFjL
8H8181YJ+NePqE7px++L+caGflWgWx/n1rfiYirn1vBE5nRM/h+zUAVcI4gsQS/l
oh1Kbg/DnmRdhmOEfBWcInEixr660LS5KGZf62ivzyzMYphVq+QwoTqrGVhcErhX
TPDiNSt1ZmWO319/xzBjoKzilPMcfLN3jpom0QufxOub7AitXubTjq/6t5EvPgz5
tToJrtl/74FwysJzWDHNpAIO4tywkPAP1XnempoYxNLbvG4z8WOhsgFKCav466rh
T1odomRJ+s/IgUyOvAYxBLDfNdrVu9A7nj1Q6CyacYTjcY2JtJlWqi+pnJXZoLYr
geAboH2bLEp8atFzGYPom9K4LR+XUcjofRA3Kho1yXXzSoDao+RfDKCZZ1hv19RI
ROOwS9VfLOrvHMXvtFb1vszbFqtuGjHgwZa/6xiO+mOWnRXomWyF6SyTrBMRGzMR
QcqnBc0g5pcB+mHlwQKWYkOOYfx+iYKHScxq2oEgw40/7Zxhg7OHfMDuLfG/46ql
5guK7T9sQTgS4UM8sEEHQUt2gVxO9jIAUzqYa2pO0kQSuPrtxoyOTUKbQR/IvZBu
M6n6N+CRTDMW3JPBXhb6E8HoGBluLfpFzVf7TKQM4SlwmuwqaW3om5QSmtNW4+0P
SIWWdRMhNBEDG7KGsHtxE9O5HCZW60RVnce4o0BY6xJRwLVyXV0JMP3GaY5B6T0t
LsYkFZLOTaRphNpD/PUJpb9snBlYLDuQ9aAErwi5MqxDJ1JDVhyHJmotkK99ghBs
t8UlHOPkGwCkjkTvtnOK30STOMT6tjOMfpEJQy6pMUzrsGtmRvwvdhEH1iLIqa4Y
U8F6vV0jCCxIlQpECU+9X8HBD2aT+pOjoAKI3a0VKDwdKw9N4VsY2fAZpcCY+b6F
`protect END_PROTECTED

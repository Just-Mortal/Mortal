`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2qgn+G7jlzrmMUYC9ykQ8UC8QfNROsxlq6YWT3GbjbBKpGE7nWCSAFV0wRadYuF
/RIdm5xiFOBKKXRCwmKJWhX7W2hzNb1iszYqn+hW+nGLAxjAc9vubRrBnkg2iiRu
yGsQvR+uDrGlR9j2evJQaPVHHXcYyNU92s3MrYzAZvF3QY93WYVWRmB/4IrkkpZ5
3IXXrNioVq6/pkG5lEMyZ9S65VggT3aj3ZVNO1QpL30kAKpHGNfzQ0Nvadvzn/FD
nXLZyi3DaGFJtg/MBz/aKNYFRTDEiQlWikkSdTPTKRFDB9D35PSygrmY1TC3sOXh
s0/0R9spTKJ8JUwmmRK77Pgwa9kmCIPNw61reJ+JChGO/bn7KE0sbqcs6lhi7wop
vcGX3+8FfKId7xmd9e99S7IPUbwPVy2RcY+X3Ivcx4/glniFKpTWpBn/8rGHhEBB
DKgUqvIfAn7EpI1M+JQCatFlnK4IvFUYFdYF7Q4FuEzAZ7jne7G/zuUEiYvAAbOr
8qViSxohQtP4tIuR96+PCfXYC2LUUzFsA5GZDAUmDvSvEH1Ue9FnWWJEYPv/FQpU
KNTIFhZjMHLjigj+oLqDzmfZ7hWW80G/PPj487s09G03E8sdiIJCCmSbl9AB2AqI
JbYeGIJjey8ytJ8MiXRE6rb3Uf7OS98gFqUByd5TeUvvJ12M3J//33GF5NyQ8m+p
rqnvxx83KJrfdj7opKbqkU56zYVDgdsDWQS0cv7sSPsYn4V1ZHwW4k1s3ILjE5W2
dVgYtqugNSwHlh5enLelOdKTJcA/RWtL4FTiFEAfTG8s8M/SVe6ZNsN6kvWqJH9O
uLXLJinlhhXBEhRPKOF2fjHE3OczTf6uZGM8PLnHCav9VCF10pn6//Doap+9lCz4
px+JCey+ijSkKAKoIXrD4dkevp5kIcRWyXfwRP1RoSJ4d+Q+CNYJ6PqkVRfPd9nU
edXySrHG5Lh6fPkp8RS1MWABvUSyQuu0/K2f/fKyMyT4pTNXsHR5Y2L5jFyQKtE5
WmpFqOMWFJHYxQ6W9AUZx/3GbfzDMwhtBPwd+Uw0KQB0mO15XVt4QfPYmWAqZtNH
ZDVgYpbC//Y46Ane/8nEm++HTEB4aTkDa2XRYP38+Rh0GAPqseod/rJ89QpquOaT
rUZuSrKsqnUZxeBSMoDZrlkBcG1/Kl9dRjHam0wv/o4RGUe9Jh96qu5Xra26907E
dZ6gQGtH+18t55K+zP9mhVHuIfYu/9E+wlLZV4rzR9gHUoOEIDsK6SNe2m33v1ax
Gd+FPXSQ0r9STNXdhAhMagT6zBCDBJEP2OSOtbUo+ldZcXRHj2pQuC4Ly9li/8y7
13sa0rkArLclwFnh1KrdaVAPj/cYNhzQhtewA3y7vUhwScWhOaExTUjCQN9uy39g
KMEBmIWvxKUQhhQ4KWJ7gH23aAorv1jOm/d9eyEXzKM6M/kknfVUtOz9NfAx4HMy
OOP3j/3LYC2dZMYyDtODCTDoNxJOrjcJinuLmoDqBX3PHSPCXwcptd9RqMcAHURF
xYHAz4C88D62e9X0MajXb7XLoGLU5HclCjYFsRUQxWqlBbLz6sytlpLpGx6hIaYP
4VMtdUTWeBSQndsIbnr4osCKMGA0azr3y5x9Mu69jbqzfgFvkGAKTi6CfHKmm+r3
uLcr0mBIs01rI2ENfJ1P1O7NATxBVqE6kOcbH+ZhL8FeS1Y6qxuZAbYF0sBJxPnd
tud1PaQrBHA3+IPrjucrQ8+IQncS2t8YSafOoA7aP2BdONQUf9b4GQSnrmGaLt0P
N4QdSrxH6sWCe1rtIqSk+vBQz1klByzmQaDRvraCiawzC/iEvCDtqNUbU1bOXAIe
/PSAR1Tc4yCwJhfJd+PiMVd0Ioh7rUlCpcs8Wd5Ii9RYRE4SDJYJJqc2e4+E+hfo
SKnsK4Nu5vLXzEeEMTTQ+ko7eofCs5tyaRsGrAPKKaZhQ+sVwKc4QHd4Fas7SBAn
5JzhFmGhyLsF0przGYL2rgGAsK6rR/6gokptKzXHagjKPr3ICS06GV8rpWg2A1jZ
7IsQpEOl3GCzH9+RLzNFoTokrpkOc7rKsiZgrT+WosqEW3k6LdPgWBwZWrcGSebO
CU79EC0ApIo1ioUL+PUT9tWNhawkw1oVdPvBKS+BB7F1FOM32oJfDOO13VfO4Oe8
So5KLZ7RJ4OlK1hUZbGtiP5unL1OQ+iR+46g24aSTpl1pFL1aZ1v8RAUg+e/57uW
pNoXN5jzJAOtFZLgL2KZFmm5muOXDNvGioPmdPxnANbf2qXmWupNNl6i2I/lV5gK
nFXoclRJG5sVQZCRDPe7xpLBfFe9PvEK1P146dw+/BpM/tZWtbRnvkb3i7+7E/Rr
JK/gr9sjYtVZK6lI90KCNn9/HSko140oiSLQVBboFB+7dDjpy4a9+poAoR3D4Ic3
WZbr3MrUGcSB9zKHceDRJqKTPuHx5lMZV9zMil6b4tukDIBi1/ab8OwBr0ugYz+x
qcppIW0UlU1lO73GA+pl/y1QTHM5BoBo4Ru/fSxaYA+aZc9omZv5kUJ3LMao/T1G
ZQbD2l2SCb8E89GDHXrERZiVeb7OMmjhDxc1a9cjkWdEKmfqTRxh4IPWwJ1GqQI4
HoRZYQuk0PvTbS/sHi1aMZhuNFXHGWi9yK6BubqGTZObJQfTvA/5z0GWA5mfKSxm
XfgiCdtKUDdz9EvGBjiQRu4f+3udAtqV4CzHSut4KsqNB17ugexS7q+oG1upPJgt
VE3dZ2bY2SsdR77oGeH2IQiT/qNGPyg1hLwwVOuUrdgQzAh+eh6k53IlNyE3Zqwd
5pF5mRAd4KxRiz2Ccw+QJWU19O7BZh3diSTtbdnlNHDOD8LsPwahGi764rSa/TWv
MgrWNRQvHj9vXNn0852v/1DiPu73z53Rg6L+CoX2rffU1wpY2bK0dqEEppnxuh5X
UwaewEDgOeaynYkQ6qznWgVRUyUz8yE0aB93b95yUDY++gvnNvuD9t1kzpOdFh9O
JK+2/+qOA6Yhv3rZ4bSzwe0sO5FyFDY6c0UPC8XbnpOVA4RlQETlGhX8NHrpGlxv
lCskwD0vilYN5tgPx+rFpnKcXjmxaUS0f1CW+wuLoxLcjWINERi2K2BAtD2gLUYO
9fpYt4TxQOC/4CmfLMgk0Hm3m7c9yzuxcMqa2tHUDNa72PSP2uK+Kr5ti2ceIwkO
odqxUr9C5Z5ntZ//+7FZiXudQRe2yks0f1s7spJUsiTnwgsTeyGr/FC2A70Ake8c
7+cO2bmFyLoHcVVpn0dKJQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEGXazTP+V7dOxlNcHwp27980iqGsk/+gHRF4L9Zy/BgrnXOmyOxrk6R600bcWPI
Xfn7sRZmiY3fJLTeuBnW0zOuPiyi8DDnzXU0GDkAmvi/pwCDDJaaq/Ak2peDl3NU
YiEy7DDvzg2LOh7jIZGiKt2xg+VoBhAX3mQ7FTosmHmUShw0i2cook3Vqr4290vO
fwbvC/khCCwkvAoo29fkb2v5ULvA61pLo/1VFEF/tLhrW5iRyTm6C1RQFghMm/0J
bbJHvQScbd9hwivLKtAdN1O5R2e8cwjPzr18bYYSH0Frev2A6dA884c34T9t6ivw
OLRAhyR0at3+u9cwsAFtYbcT9+GJNOiUL85ygrKKHdw+UihOn8XTti8syW+Vj+EX
5A1nSdMOMh4NgIcr6fPEfFixKBmckNWisNA+/Zow1sVUkf3mkCzOIy6pncKhAP7I
mvITi0+4PDbtqP5j78tPaxBpvvHixMD9fQv9Aoya1QRORd6Fx82082uPrbKnhWtg
272xBLyGupMsCKc4nv9Ev+usZWcmKrIFbEXFzeQMxUFDmOdi2XtErimYTZoK/ANx
TpXQ+sWhVxohQr75LxOm9AQyNK4GLiB92AQL58oa8Xt8p5gq0X4SOtVecwCnxIEJ
K4bYWyD9LRJVdwDA/2Jr/JKMayji3JQ758iAc58gd2U25Bz1DQ68SaPadi7MCYXb
W4BDjxE45uha4YCo1zTvWi9OlCuOrYSNbBVqUjx9DMSXb6mdIlmz56MyzM9BN+Kk
EBhk0PoiCGn0YEbK2k9C2/sf+GEbiwRR4zOdoQ9eBFgMc6BOgs4IULHfh4K9/046
k21g63TjrPAkJ8B4/dbFxVpBxgKx1Bo9HHFw6lYJ/06fog0sl3zHmqZt15TF3o89
7cbh6bjg8e703F0J6q3Jx+6j3P9weBH2jqOdE6SPt5L12iO0X/RdIdBXxPED/S+S
FLusv/QykEXMPZKga65CkQuKhdkNlXc/rYhELbNKCWZBb+I/c2UNOuza65W9jRgO
JnN1FZreBhLzkY30X9de6HGEyW5YCFDUKVlZvR55xs0wcWO2syRA2URojefibdLP
b6aFuGadeskQLwSb0HKL9c1ztfh49WdrSCD45PsSFhMLYQohGEvKtxrdrX0BfXbd
JFVjW8lvmcIDM590EMEJ2eAUyjsgG/Q9CG8jFRw8/XMQyFT1AfVKBI4t88/iCcdT
DQ7+OpCDg/eCapoLyiH2CbOaPbF7n5svNevWcdbJ1bgwFzt0BQenHVs9m9Ko004X
34vl1mRgb5dmvEa43S0AKByImgkVSD6VuEKa+jbqMdPGgztngXdhnzlAMYp00bX4
dSCvWvUyc5mZXYF5p9D7AOPMLfiv07+yP9nvl6LJGv865CKURfK4nYcsfn1vjhW9
Rz6mHkLj9/QcaHgUwpDAmJcuZk15JX2/Fct3CfehBM0gEZEjFt7HPFkjybj4pXOO
o9AOsAV/lnLFml+o1SrDYcS/eJXOZyN2tE9sGxc4DCDstmgof2C597/yTVoO13xk
WnSAWFJx72Pimmguzki8G2a0MVnuPqqoaRunZsqFDTPPqoDoq9Pb7dEmwlouZglI
hW8VomrH/GbrKp4R0LGr3ejMWKY+/vB+HkW49LVG4NQ5o65TLkz9zFIRrSW8HTVf
C0quR2+y2NbPCepi7f0DUw9VuJ/fsAHTikHP0CdcpjTi+yN7nAN/xljEDXaedE0x
06hxDQF0Z5hdSMNoNnMBeP2HvqjdKcWV7LIoj86UIshvJRe6QvyJGrS6mNvcbyfV
rGrAKI4yd76s7iWMPH5My6GLqbTtdPWLOzIDzpzBcQKAr1ihrAXtgCqbPsphkhj5
5dAP0BFVpkmE+XmgEpPa4LjIH5e/eoZJjsx/rctCGqsIsxE8WJxVs9AvzNh9CEOT
5SYc1d87ns9MtIjiWpJgzoLfdHBKqM2tJjUH6ZvXfzH5NigczryPcr90iPJ7DGtp
7kFOQvZkiorpTu26NOsMhxKNTtjo9J7YfQPAtqBQRsAWkfrUchcZlDGKm/aLqDIr
Vqh6g4jkTDrSej/tgPBUb6bViZJ+4rrv64WCFXREwqHRroCUz5iMXxYVqzb+VyPR
0h60gQaRD8RU0dWKWMcazMLXYyouxjNvYwqV2bxRIPdiXQ1cxFTDSRXSc27/xmSy
UbIU0f1injeN/0F0Kq5JqZmjJG/zl6Cnb+uReaBDomj7luwMv6dHh+gKSjZmVwaX
XMu9svsYeuZTb7Ew6YMMC/E903wAgy0E7CJUcPbnjj6zYoUvHc8X9BiI2smF+2MN
Z9BpvJJ9n/ggQRstAW+XQxh0dk5qw/qbrj28oI/nCCj3nVCoc9mLszSAsJzDb4Vc
E5oeMHuQZUb7KbyxoQS9gxmW9W9o07GjoK+phAWll3SO/bS6SBaz5SNx4BhH8Jsg
7EgxzGn0jac6n8JBwOZglJ23/+mNTRTjfp5PAdti+qO2siTzhiiM9hYKn84Ty5TW
pOI308IzcIzs3qVvNXPz5Xzx4OeUhMn69swyD7xYjNLbLSXXf0J8NNLgiCck0Npy
sQSXDcy04+WNCaxk2p25z4AvNbNUPfNlYw4V2PFPmX60rmum2PqDJEiT0fR7uP6x
05GrDxo1ZtmJheygVs1SLoB4CmSkKMGExV9+3O/8hFdLL0bVSLQ318UqQhC2gDwf
FeMCjvKgOL4vfc6l6/E0cvkBidmD1VneUqAsQ3tv6DobWAzkK9gwbbCZbVcAzVTJ
WaN9y1rD6zEh3gOzEvkvd/SJUHCnUqHtJyntd9mZBgJuKUgKnOVygEMaoVNx9355
oZHLU3S1sca9ZRK4wlYNbyPqQx+adSNjRMQUtk5H1AQZfAsuEXKC7rYFdwSv6G8w
i9e+AcdCW9Ey3VlAay49bFc6RCkfjvZyDEr5GrlfUUfNP4mX2sx8LfLSl+4SX0Km
NYWZS9X4TW2bNWiKTBzqy5mDKmQk8ug1rflJcPrjKOC7Jqzpzs7eElXG/2NQhfBo
krfWiAR0aAIuAfJl/QZuO0k3cxHEDjdLHrDddDUyGqz8NW/hRQlSvKpnXCwkbfXh
taErzsUBMA/4jPgJPBmC8TWemY2kDNJh2hXuhsd2718MDduSF1m5VeXuiNOCL9WG
fOpS3LHA16AXjdbTXaPWi10YUdeHUVq6XsV4w70VFSL49lcmFTGPk/VMCQZvHSAE
7Xug/0QuQc8DdIFBGwUG5rUGxl4p85+heAjEcYo4h0+fu14ob10tLgnJQl0I8Py1
+31vQs5ikIcTvGZPmNBcufc2cyuiyG2/TGhKw5Bb7SddGeSjJtjFlKn5cGmVBPV0
iUYUMjcLxbVtXcSl0I6FydgHPKS2qv+/cPSyUyw1QYXtYG+kM3hoE4lwAccztcM+
v9FQMbbr3Ede3lSfjpDKKnvg33PPC2VLVUo8EBjcoylZA26xGsPR0doRrnQVl9J3
rnJ5+aYeWIXwt2CZKWH7JWy3A2wbt6IEod7b4LLxFRT7Rlv2xLoeS0o/45cOM7zg
JJKEgrsvSdqvLoZsvfi6EX4dXuW9xDxekHRujjzEMlbYDGrmJntodqR5GQKXcDL9
+daLKoI9vyb1W8VKK7TdA1rcKBgNRx+I/jn2TdLoxAFrmGNZKJ/O8F9U+O47YCTx
vFC09bTtDEw5MXVXXwYWp9unPRHsfrhWdtxUpdDdaIaPkNUd63jX5CJMTQ1Hs8wp
6vTV/BdLYc8d/rBIl6sIAVXtR2/piWXHLhpxniXRe+7539Rpbh89nkWc+DtAGnEp
3un7rW8KIScXCz/GPAcJAFzlPwJRF2jQlV36BgvdH7E9hpZqmJEYgZruB0JUX5fJ
PPcIr4g15H+6dawbgJV7iK2ukGWTYIvCJNoaZoIgFx9DhPfFYRuSXvJf95z00Kxy
GW4eYwydIdroDmrjUItzcV+y/9u12AWyTrD7uUQdppBuX6HK+BC/wvEmmHH1thFQ
krm9DmvwnWsGrPW6JzMAi3pFBYrjZk+TBDY+M9pXgCaUiqpYI7Jq7UaRj12hCnzm
ID3I6o5Z0IZw2HpRYgAsflq5OTND39HckKf68DTgKVuZz4USH2wfCi5D/XS6VbUS
IVOCCg3uJeG+Vg+an6IONJ50xBuntkIRd8fmDtaCybWBzDzrvm2oj/Ts7/lJDA0r
PYef/iJV2hKeBvrOGTKxEl2qLnVpWjO78bEPzbjiEcV8MZvKRsogyPVvJCvdt2HK
IVGu1fvzdwveilQJehK996yCMLfHFF9tJl18w9J7Fssb/PDVQCfzl6wQQgeYWjay
wWmLkkmpKfRHVyyBcV2WB+zBReC526hLq5X0ng3RSu8ysVQ/L5MVb5awev5zmAp2
xOAipbdUu6ugdTHHhbQjyYsTHnZzoLZX7hImSYfjRgOAo6QL1SNBLB5o6fRS3mpZ
+a5HAfbePKDn770FqW097/pMno0oMndZV/1T5/OFY/2eVE2N8qEclYLCyaBKuBTQ
`protect END_PROTECTED

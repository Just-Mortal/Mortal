`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HoFhvikFeB5qhQ39/zHjDED4Cut3PncfkbaRRv+TU1kG8sgIvANsy6em5r12RYJA
WHRiSbkNHngmeM9J/iHibDPHmxsutsY8siUf4ANCPOIAWi50A8IAtK7KkhJa7Xp6
DTsuJAfrJuHHmd24RxCyS1DHhOtVOCkHY986k+jS+j/tDg6bzSmkWmwCPstrMzle
q3qw84VTs/TMirVmZI0+Ktuk1x2eZYcmU6UQCd4V2O0W/XIkrpTXxYZ00ObQ2UTm
1CN0ijU7rSp/smEYcry33zbVeiUYjTmyacSoiyyaaeX2kPwK559aFOLZ9p/tV49u
zvVf5NSee23A0olp2U9f1bWTOlkUp5WASN992EtTuGgutd2VY619NLmg21MNU+Zr
QVkgQIBW+kBSv3CBuDLHA2IVkNOltKW3ayGrvVzWOQ4kvErx3dGrwJIPVpiMMsEd
xbzaL+xdsfRnRhY6MhFvjw==
`protect END_PROTECTED

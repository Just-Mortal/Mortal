`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c+vC3l/f6YxEB/hZ4ZEtvAZbeMRCidmPkmN/egX2eGqNQokoDcZjGq0jppp0q/nV
uV+5hllHVRero6vWPkdsQZrfxpM74RDdA08LLTQtAkaDz4pAL2ZsB45G1wjxzBXJ
GQlxA/H3eRh9eHgyACXOevKnyI937oAqi5rHDQu9/r3Mz4oi0asrgxuLUtNU6IQh
ZYbt09n+DVch/i4oS5MoyB51tfMI6lHfIOKDNNIoe1nMGDqF7bT6P8LrJ3y4OFrx
H+CPhl93eD47uYJaB6EeQN7GE3Urnw/nAY7CFKIdFO5mp0wppcEFROnTEJi08sEz
957wpS8BSDD6Y4RiBzAzNjsBTIbju0ymukPnQ0s2o4S0jYh3GNNfdjRnS1VAEddL
kf/mFKcIdzFMtzQZwd4xQ9BvYgEedW7ol1n/QAgV7LJpN+LFzWWFZz4Ae+G07J5v
n2+u19Mlw5uBHipilsr71pvv71uJ+vaXAynThukshVGh2Tm/GkMW5MqTqKlsTcz0
l8ShXaXTMwquvC71YBw2d3byeCmSB6NvbjczB1nC8g5AtYSF+z4Coz5ATRKn0KK3
bXJkMRg+c7AM9kIfW5HVHWRfS0H8re/DqY/mQ9Jgf8Tyn9zybZW/YDk7DIIQWBi5
qT65AlXD8BD9AceVb7yNuDzl3s+B2JXFSE3tkCzj+GI+Y8ZsGqgydkyxOgPm0NWC
p1R58rlZnbLyOunbMOS8kjFexjXCbNFmW36uHOJUHfYtcCKHT5zipt6ECqzUeubZ
MNS7jHTu9dB6Uj0DBE+KDsuIkPo2QmhoJn0PhvMLjIEJOz9xusoZfRyIFNwUZ73a
RZmAxUqBmQSkYhqBeiwUxagb5Ix83xWWtlatJTlU9+TbuwOgQB50XmTdVzZz6/Zw
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ntVbH1FrGpsFqpu5SrRLRxKc8tlgVHDxQWEM4K9I39UD8v1zrLEpNVOkpSOSWWG3
QemRDJZnpABAQNtAvsTxFmNBdz5IcRAh7EAaxeLmlbm+oKGZ84GUe9zLknbyWxX5
6SQf8s70rVEFyzzgKzEYI56HsFpEv+eeL493YT6LrnN441kkSi+Xv9/xyusMbX5S
Lyccf2eSogCvLB392jh8r3L1ZatRoQIu3GbRDd+BiAHRUVQiLMKoO7yDGi6XXh5I
uKb4thagM15iaP1yUv/uKLqnPhUnpZV8t1+QOeH0+SEItLIqFmSk5KYbm/3cD2Sr
SzwMttTuScVenZACCtxOtQitBtnkB8t5s0PclYIvC8OD1gtdiMuN/QBhckFt/Azq
vRvyQr+2wyd//FT5SLcEJK9jqyIjfIu+JmSGvAzEyJOC0JZljzTHSy3IqtLFAhiX
kZ6l3Uj4ZwsZr/HnG5ELmkj+KALUaYjtGzSe35MKSTDDMWC+SBPRPrrli8efA/Fb
vJdAU3QL7AoGHCxGOdPydH2mSi9aAnLa2yj/egNtNbwwHC5U9Y9C9g0OikccO3Xr
VAcHYbSl4xH+dCrnWmyV2eRQEo7CARI3HW601qt45I0eTEMUbmOaKR766vqvwI8B
+imNrPBygteq6w3WDUxV0o76xhi/mCcF0fsp88FdyQgUzqzfRIP/iRp2qqaWeP8+
kkInJbhuJrlersmKTUQgOBL30yp0AfkIeSeI93o8k0IQYFgKJ+ikJ5NalVGPtvW0
hciaiuqRZ0jspqH0uNrUHdkzFIeOkKntJpad8RTUXDXBTqsdP3CmwCGO2ikHoBF2
NOZJDCOpQGFZ9YgxX8b/XfRTaCqvuiFr32vhpmL3MZjjYWe3/iFJ65KdWMniZR4i
To7aRTTmvgC+c7a/vZkVppkJ2ChG38GFdaWf8L0QjPx0Yj7giYjvIHEZBRe/G8Yx
8emlIN0GkMpYHBl5kTy1/IkG4Yv0GTxxyP8XO+1984gW2ItRbCk/AH6k0cJB1+VS
jgPb4gBQyN9LPX2/OAeJ29N/jV11+doVFqseCUoGi1G8CbelC2QlPCgDMLzRiq1I
/1t1TGUFnLUTkGAY7Szqc2c0cJdpCWUC7FQwxoq/qRoWaRm3Jw9hEJzvSFlTFtU6
VhCla71RsBEH3C45NK5HZsZMWzmtD+006ohFyDfCxPanHZhpHncG4uGtWl0AZ6rW
ye1P9Vg5fRMcHbcFUc1NuxWuKpkheYWpEWaCIOw7hWJJDz6TpM6qSf8dSgQHsmfI
y/z5S1Ptdtb/F/C4KACzLCWlFkncp8A40tO0Kw/gpbM23dd7/SMG8Z6rfsLjyimh
VMjMISy9l4xOF6W381V3Dh1+rlwjzLW95t4aXeidJD4lTwWn1gJjXmyTdH1eKbmO
RE4Y2JfbVQU0pdoRhauRzYY9EhViGBrTz/TCP8LhVrj8EJX/YWGlYnqmAMuKM0yg
dlID81Zo/Yipy8bPv1CDCDP9RyypqfQ7Z+3HwVjYgiDlteHuD7yvzX1beTJAk3Fk
inQsac4HYyauyUpiVl9ElHb3LLRss0i88HSNYGRAHAtrPaL+6ouPHnc63i4TfsLJ
8flE6az8MmXwlTaxu/mnEQVdqNXqKJR/QbiT7U/+4LWtebbjSaCiw0LIJvktBUNA
fRdX6lzPWZ3fUQDxMhF/r/zMPELyJFr7hhu2LciXAtF6NjELvycxRhUt05G3no0M
llhwWNwiZxZYXDCRb236uk6BQpfdch7EERYyX5EH6wRlZgfhQDQBxok5SCbbG9Jn
PUVjejwz4gFY63w+GratE6q/QwDtgQ9OXXeopyhPvE33Yxa4jeXeeDEdcanF2oRu
/kXx9GaxOlgEnzsuyjbN1VDgyGWPyzU0VEf2JElVhXRKhziH6M3ROPY1hxQcmSjD
JN0BfAUYIwCmraopPP0XkhT6CTbEYYBvPlkEVmsfoePLT68wxq/1OjaglPbxc3Ae
hSVHE+7Bkquekp/pZZVcjCioFgh4BZIDHp68P0MGWXFXFrmQ8p5w5Le6de7kFB5l
kP+pawHrDmk40NLZ1XRqwgBM/zxE94yZYnc7lqDKAiyTwtugqFI4m267+NlbIIWz
OPu7yIO9+sGPBv1AAqM0Xfk/+AXXwpEevKK8TJV1KgICF5T4SLViJHa9i3AuYeZw
F+/Zjc67tBYPWS5XneRZplKYm5Mbh0pZDE7ECM8NPdcVuG8gBaLvBNBwQotgaU8h
ux45tMLtC7SO/i24AwxfHE1A0Ygvg33EAH3HAlnIx8UJUl+y/DaLFL+wP+SGFgJW
YQrkf0b74GiVLk0DFzvkI85RpviLav6ummOBZadN2619vCoZM0BzsN2ljBoPsChp
QFZQmWnCnJNgWb8Nhz09I4qSQosHEeonMKD7F25YFEb221uKVVSISIDzsvD2qAQF
GVaUM7mfWMUZzSDzMz12MIWNTOairfOQYfHyjt2KzTdgt7LEomYdV9cGaZGml5xZ
vCtmLAeApULuCM8kRIUdyU9Vj37dfAynQCquyE8kGmk=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9pXDtHOzAftQs6CQasugVa0o+YBTljD/LITKVnBUh4MClgaCjbaa+39N3lkcogwf
jPtw5BKKV9k8vdLaMhpwZmkOUfla0Vh8zrMHFDJXh7rZeAhP6ROLxV+Uz38LF09A
oWWEMySJ96xVMuGOkMjvnkpRfgzVAbaLkv1QbyBQ+EGQaesj2Rv8oD21GSKMla2w
xVmXYBfnAw0jSOxJN1k6gb9tTS+gd2OP9ubKBmiqal69gbNEZgKZ46f6ug4mDjmL
L8dpdml7H6hTEKc/bBfXOWun6zAiXVlGRV9ymUCQbiXN4xaSdPftp26JuAHw7P6r
YoZJgfJJEO1hiXjpQuecMLYFth6LaKwIdr7aubDRw27h6XkQftyO47/luLfnyl0C
fILRMFB/bAaxRsTOscQqwEbdC8ff1jqcy67FKJ+66TzLF4AxtvXm8b3r0zoRg1ed
jRFkfq+KMsNitSzMjyAVjvuMtewoci9XhvuUvaFRARTbmtkUzUt6IIXYaNgn5ZB/
I4boYmiIvAWJgQOztk9gFNLpMnjbYBb9er9vPTxf0rrmsKJVzOJJy51Gusp/uhcu
8745Zw7DPmLQchpG116ouPPuEOMYKLGdui9ObONPgQX3mVz9HMDfF3ijZXfULfAs
N9z0BowZwM2sVk5Bxb4dj3+gBlWim03tC3JE8wB9TCb/a0xEJ/Mx/dGoDsK9bu/a
YX+j19PNO3oKehxO0vDrUl3eQylBxWOWXv4rvVUlCjkeIBGLv8dgx8u+kSkJq4uC
DxN5mOKFRgtEvBUJyt2mx53ekcmDNJaHJHD6Bbxy4YTimuoPjnF1kB3TBgTGkyu8
PySPuri+vUtgz8QIe1s8oNV4D862PRCpDuXps8i+Olf8Wdfig0wi5S6nt53h8GKj
eh3FUBYQYPBDxsupKHAjmns7HzTvpWg8cNfxuiWL8B/hxgyhm5BUcNDqoiZENaVl
vAf0EWtzpjti74JwCTiaH5QvMYhXAWrJpNeE8WymcKfU7nbJzh+p0zgTOq22zrM2
pNUnSSsTEcXt4SEYUshzXEzWDpjNuezjBOcauollSoE2HOGkS5iVsmJ9Htn11Huk
W5K6OJs6i6B0O9kdtistZaSJJX161c/JQRJDqCiH+Y3GLn8mGUYm94j1cnj3z0qx
EzcMZu77cvJtboDuwJLz+JM5ulo4Qoz+XjI6XSDy5UFMKq9AhhPm1QzAtxuh7X45
WsobdxRnGsiBGYwPwOLUZi5DCYwrZN+fXl+WSSnezfkv/yU6/A12mV+7C/K6tNiH
6e4m1oo6e7Rk6nIoHk+PBYenazQrkTJtcVRrfvQ/QmNhd/RlbIP0CEDU5eG9LqGo
SReWGEMiuIs7AN1STnSTaWVhtiRAQNW8zMpYQe2BCmya56jRAViz5Ezkbo3BOXoV
/FxcBBNgSbQQ5w1MY74ED5/a51v7ioQP7YwHtDy5L9yBWUUDsiwSCKkVsKnwIU8v
rJUWNXZM7n92aXa/AHjIcpJApRf9wvnPpsKg5eprx2ZYRho31wbHvREOhn22MffL
gWsszVN7lxWA1jhWz7dhHZA260LWS9nYVdpYJlmm7FKYhmgV61i5WC0J/z+DcECT
5emIl5hGiA2xbVG3g7HphQWHOFwkeyyGGfWdTXqNndnHT8Zj2d0WKoN4gNbNgRlR
kHHJ+pIBD5OVI+n/BBJIe2JTMZuHcTjZEwf/2xIWHLMP9fBBAAMfd4mBqFJxgfSR
0iTVwx3atThuCxPSqDX0N0qgA57kijxkH9RwtOCqVJHYMMmL3dHRcxPVfZDiBAZm
HToSx+gUPbXs69fNJfdDpSFVYUp4QwxXekvyafzK23j1Ni65pM1IgHo0IFWqe72i
PI/lJ6Eea3zvQf1lMH8KntnNFuM65nOP60DFL3d6zHFKPEfvxYZhmowVtjtQ2WCg
HgB50z8FMOFwTullnkgv4w==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7tXUrpyco5cAWupe1kXdcaIKpo97MG7hYHQebQWm6ZqcylEpbTTYYO+NE8A7EWmO
Xa6gOpx01cedcDeoqY99xw81CpEV09Q0K4XGvwJAPGE/i+/BDPXzuuN2QlFK0vQ9
fSyriycoiMtdfIqUEMyfek2+taX2K7/LqLJt3C3tz9rws1fyc3ySUkEnEiODKCBW
8z0ga3+YpOr9hRyHRYnD/jAb5K8wieeAjBTcG3Uc/pajTs7qs3mLtXQlds7skQHi
rblvkz8iil05R0lT78YEzNfhSXWciUTtpqpD2k0Oi2WIi31AJGGW48eVplus2VXU
PhNnjrx4WDeiBkjljuOv0eIV3xSnVMEArY76nJstwLPLYex/5Toz00xIoQugLmWH
W/oDJBD7M6a0ofeeB5oFzQjHao5GBWuiQGnUVFUMnBJmCE+/AGJceqcgxcjkuYv5
Q0LeYIwrtxo+tdlfd43kszZMulmuf48r4NjYTfdcsbGzkIUUPRhOeWSNIhpm02D2
A4dd3+rrjFaHuI9NkWhmY9311RvrsXm4b/BI9pUgqvetveWMG312s741mUvfNwH8
TiBXT5Abxme99D8wjnkGV01nX+uqFZ/eMO67aGrZq1P28BUn9TidqWqIPEcg0Z3R
a+cVbiJpVTiO2pqWCpQ3Z7vHszhO6pFOBxKLKD+EHDV5vVmDsiQf0ZRXM1enFVSF
/DBX8kCovSaYSwG3jxki5FgAZaPDjgTVVvtYr/8ov5FsHwui4wKKiK37fFdYHpIB
8zV0VF8mN0+2wnVOIdRxlJOCgQfpooZElgO72fxBmfiMep7NzEGpbEOvktZu5Mf5
vtlt5kef1GBMOQ4qsxZnrFUuD50EGWRWReyB0NdcyrYHNl7oLAY2NKnWMl12t8Xw
w8hBD78DnQPOy84q1l3B/OFQXZLBYDiiYpGTvEYExwqXHb67EgXdPbLna4FEaA4e
O9zCTP6ci0crvFTC7Mgo2pzr4Rcvsga2/N6vQyTRi0djsooX3txL/gPc26/ztKO4
7JPjMs4eVFSp5J69qOb45Id/NbgPOBO7krWNEYFVh+O8K3bHQ6+FGNosj+8k01sm
xn4LX8J6IpsPxIIUUop7dyzS+N5797pXauXNhJ/Pu3QxRA9EFP2kgMOpmT/hWwJK
iYwcfOHmNuG4k7p6Phhk2zWNjnP07esKjjfmiao4smskJlZx3D97u1rbXSUcBWgC
JKgVR0+dRGauLEyndHKc3puXywT/zDhu/butF0VnmjMiNlHZEb2CPhUBkfboKrWM
0hw7wfu8rv46g398iILc1EXjkljyeovNWKv2BV7ojR0PbR51hYEWJoR0yXWMJtFB
ELiKmbB0rLO5qJ6eJIP/mQ7RomGskfpMrAcGISX5g7dabWZul3iwE4D0WiikI+rA
kEu04ICrY7KVqfE7eZMdbbQ7d9BQ171thXCGY5W43MjUIjZIBj6eNqpvTR7rUFmJ
oujthEaFc2w1gWNPieLG33HY2kgz9fMji13QOIWSMt33v+72wjAYT/lGeoNN48Kf
YY8WuaRutsugHntU8Jul61EIeBbeXfp/nVL9J7YjTrn/gysVNJXLSLsGun1GznEK
fW+XGcURpLK/lRUfyx7krUODEyi9lqS4UOxI+ZXHZBNzBKMrj27ZCdSUe7VQo43z
4jHHoTIqLe9dt297Vj9oGFstvkJfvu2fWJnIGI7QWCr2qf7P6ncNI+Z2IUfJiLnJ
g5iMbgtGwLPXh9WmL4EYkipCNba6Qtp1MlbPop5w4wNqdtVU2BxIAUpbqRWcWpGN
P9oHp+690oIEgkE1PiAa9xOQgTgXqA3YPXA4Z8GPLCLL0ILS1w8Ci5Ab0t9D+gSK
oCOiJhDVYboy1XvKPGGg1Y/dWKziYMKbM1S/8xN6zZU=
`protect END_PROTECTED

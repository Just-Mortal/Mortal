`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSYqbzRDZlybU9z/m2dGkfpjhm5OAMY8TgnBhGgLhZVWDbZ/lMybc8wH2Nkig1eF
dm0rkGzcU1kHxdIbdh7Ngvd/+sz7/nPBtivhljO3CMaApOI2fBStc8ObxAxguHT1
V2e1DaaW43v9JnZCKLrR/qsS+L/8mScmXoYVs4965U2QAl+PxJlwhfJUwRMrtka4
jKAfJrmtO61RmgBXBe/7nN4cxh4JjRermDxoNh833/xHTLQs72RildrOMIsW6jlv
wvZTDXPS27ypArxuOxHUfp9wgKmcgy+GEKusFSorY8U0dWam6wZIcTgHNkKTRjsL
EyhKrbVMBUZ/2Pkb45g014J2RzuCJlbXQKT73EprivK9kjWPlyao+YyX81W0zbeT
eyU9tiVvwPyzRbjnv3rmlF2nLhgmf/2WBnqVHUWrtXg0rqXP5vahWy2I3t6GHvi8
Y+DnDdxA+nFLIy5euNCSrnFcDlFluICpraelv9YVc8xTgQdjdj9UD9HY05JAnOam
CtSglkviwW9MPeTnOmKA8f7XvJVd3noiI0h6ngoqOetFPTZkqgFKbI3t1whyRw5H
Xn6gYXmyfuRMiIEEtSNniitSm/h17lK3ydxjfTNxsjJlOESaV02xFDifIc5sj2hG
EyDIQ/2A3W7W6mZJxyUykxNMM0U+bjsS2+BQfFEhjOeDpkOXBNsoSwYuf4p0/zj4
7568QNfwbxEL1IWPWD+WnHVsx//38pzxmEJzRNPaIwNcHaQGjO4hDZHdWjO9lDux
4vS0CZkj1Ij3ajL6OaKh0582y9Gb6vtIVwMTXv38hIQ6zbHpaILKLAAjCoqntzwj
oBqdToLVE4v6l07nEqSMT67cUcFwWBJD1rBTfDs2F1RsUB7C87T59RG7kDXMG7B8
WnjYRiQ9em1SDt5j0Xf+1w+1SqxRy0/2LDMlX8hmbcVK164NerPKyt0D5Z+CCmDk
BF1uYob2cdvLsKakIfzstQ5XS52NHpwjbS/71WLsugImtnWex+HOnvX82/N6ds3G
bYbEWUGxiSWWB/Xh3NTVEMBp/RP4wE5QLwRERQx7SxGBx4nNZPxXeAuHYcxZ8JU7
m1q6HDLULSSXYfmLhbgXrwleza+ZE4LwNWMceF8IXHW1u+V2wU4W8/XrrFRDnPCO
6o68e1ClgitvNVhHlkVkknJ4Vb6MYHD2BvmEYWHpAcNBw8CJZH6govHE3svyi9Oi
hfbmANksxusxlKpDIpvOPX6PoK3FhHbKNtV3BeW1Cs4W/+YKOzl4WBjk1l5wYqLF
+IyPa6x8zMVv4DmvzzuDx0HbeQ4HxLnfIy301Vhr3U1rDn/zqero1hWBfdOahqUa
5I+gahFSuYCcy3cCx4U3QlglGCRi6hSIRmKlVRRkw2Kjiuo0B+nqeA6LQuPObYg/
vrp06pR0sKD8Wn5xuX4pltUx5uyptEq9OsegTX/N7bS9E73a8Cqzsq7j06x4bEbZ
QpC4MhHDxL/FKbf0d8PyUMspBkiwBpWImczozShW6XSJmxBS1STjm12FATclvBW2
gQLkSYxum1fxc41fZBF4Nd/fEoznOQTXllVFZrH+LE9wNX0S/RNpnt7lHKTM2CW3
hsWNbSstTj4bAJkxeOg6nTKPxwlo2fJt0W7nsTkEAOBrQBKg5wTAF+Bbcq9aDNdi
iA6yh1aAMXfMyrhKBiptm0EJU6kkBhFCG1ufXvkWZxegeA0lrUxw8GHkq3GV3FUX
O78FzY9PSfFluaLRu3SwmXfGhWzJGMBLFt0YliguvuIyxZKnLCQfQfEVF/g6f3jV
i6sikVux0y+3EUA0mBTM8w==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hy8oq/375vKIPME1Phr9W/pkBWF+N9QAUwheV4/N5kw+oAft6Rj7i8aXHlxZRG0O
LluwR78H89lPISAy4pElorZCPOKPXH2wYU0kGWfwcPIihr98hvGczfsVF+Juz0jk
uaqvVIgQPB85O9/0MaOWMNr0uYYCUP7CA6eQe7HIk1QECqYyK/GyqbONWR3A0Ls2
/XAj67S9AIFgliT5brNNx9D3HB6MiW3NdWsPI85A45CPprV893eA7XW8xYv89Pa5
qkCfT/3ZWAZSdpyRufzthpVHlmNmqIia1RLEQZz1UQqw4BehL+fK1yrBA/usq+R/
albVFHEwxVJg6ME+2EfowbuguAlq/TFAQVwrh0F7m1Lpna8GraEvu1uGE05pWfJ0
iEFleqX3nvKTEWwD7UXtBGr8JroJK7XA41ZvTnZQnForCsE/NhlyCrwSiCSYKGmX
TK70TxBcUvLNmrHtSIEH2wfp5eydl7JdnxoGOgkYHMhwEvqjl1kwB38Xu+/xRsur
b2wbf9tFYUFUI/uZ6oRZyddGVxo6t3pWi6gLFJ6wdFVzpCPvV8cOo61oowSKyIcX
9OCTW9WnoEuWAI4FfTe48Y8xvoUBb213t+T974Ik9NstqxK8YLVZGKWP3Nj8Zsfk
UFMLfu+Dq4UdwPiQAb6dNiH5M6/aKkj8MKVvhHv863fF9jn8PPbUGU3zXT0S0dqb
SH6GBKT06uVxWBz85j5RAQMlt6AOIivd2uPuTrlV10QePF0wzfU8DX36ZlFBBt8E
NMywg2KiwN+Xs3JIzdu78xePokAuEml7+JwoVZE0juxDVCoPrEdW5Z7mOjacURXo
PSIP0FY6jQPtYV2m40hcqE+BONzEzlO6Du0ipWjLnN35S31DDWqM6sraDlUGYSdF
flLZQ/dD4DQFfHYNysghiBAXwiUHSN1OEAsVspkf5QNlxzl/s8vBp0ByNLN5i4TW
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Br5ZcpE6b8nyQvhV6l/gDZC9srcZM4sDShikyXSCcg0/7PJaZNd4bJJcio32IyBB
4hM4nsS7niquYTuoxZqHBOR+4Tlu+JnBCWYid5LQeeNONpeBvJEAWdYha5vS0cAD
d3TG725G1gYQqHiQGPOptaxrLKvIUXJFaDkMvYwSxq+Qiu6oz7p7xC1xa0PpOrWj
aWughRAA5C+OC2D1SxHRS4lWJSxFlXM7BRmgwoSg24YGxoF5jEnyjQTfTP441/Ts
s4AfqtSYFTgTaOtFpcU4LeecL94W1PGobsKJa3bOf0xA1CoHaFcV13ag2nu8WGbU
8at5Yrn3rhTKqmNdYCuR9mJYhoTy+EansLmdQ/X5lsBA28jTbyctb1myTR7D90AB
X2Ko9OinDEIssts72cfOkSHlQEu9QnGDJIn7waJoUkip0HdAXiuiSKqN2Dmk7qyT
mH/WkHo64wTvka8I155MPKE6E43b/OQpnuqULDH7FbsT4TXzmQ3Y+WyR4/zVXkQ+
t3SXkSeZYq4tD9tlk3spl5NBAssej7XpoFG+SyToSyE4CiCU8NiJLvAoFCG5ghii
2GqUbLIJdDdgsca+Z35a+gdzWhgcdU+s//8ZbnTVGAkjd3V57G0t9S0HkjwMckK3
6aVf40gH0ZitizaZBDUmuOzpaju6Jl5CSKkJs4rkp0yESBEbp4dvto7gxfBvatDc
uhV3cGkz96o0fB7BArHQddpZ8ku2UvURAejIHLFH+TndzcYvJpk8hIxVDvd5et91
Fzgm9Q+JDG/6PtVfSQVPDFk2htLX3vk3Rjz+pSmawaDGwXsdlLbbtsgzbzpqpcNR
rIkNR0IVZPbT1ubZFsyEaUGiXYy6fTxoKY5XMbzwBrtU+V0O6FkSKv5gsPv15667
e7VmIL9YtKeNT0UwHNNP6X686xjFnQzrtrciy4TqQL0aTpKeLJiTquZflWbV0jgS
CK/ITORuadPKc86e3ysi6Cz83OGYrswE/x8AmUeURl/AOIZxLbkWX5b3BlWQnRx9
/wY76rYX0D/oUQ9jG8UVwpzEqEhwxXGz0GKddbm/ZcM=
`protect END_PROTECTED

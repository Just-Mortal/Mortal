`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LZd38Bmo0NxfIVQolIvn6aNZRiBDmT+kiYmaNH14SKgyNvoLOk08cJT7G5TkInma
yM1b9XCGEkjw6L0ey5Hl2oGZETrxdy3/KlnOx2o2ZGSd2nl86c4bBXBZbf1sIMu1
iY9gb5Zm9Q9t7aNbKXSn11wk/LS825PXlVRjDy13crTRg6qpxdy8bdSNU+MnEQP2
30f7JJPCNuxxD1LxrRzOByHBj0M0EmAOquGvsI+GAoh1o8GNU9cJUM0/4jQS397G
yQSwjKmKRhLyr28K+vX+53Vs//BFWv77UDks7alVzPpK/eDCwtTv0uMMW5rctCwx
eTNAZNgukd4llNYN3ZIhtAgBSkw9rQBYVoMXmsosSM1IvtWvw9FDislF4ExuYVd6
3rn+fLLDUsNfVrNUXJO/FEZl7H38SdUk72ChJiOVK49PVPf4RurO1Ce8Gf9apLwT
IGP3L0ZD4xv6X1tDr2SiquOSmSmaz5OUZjmMTTH2Qvg4AGiZLLrdWVn4yoXCCbGK
GOpHYdBl/V2t7pegLAIIAayh8FiGzSeT5/07N8JN8bxYAN1A+hJw8vJqjIWMknBo
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KDM3gexxNrWHVQ6G7KmhXy46KWM6TIEiQAVi0Fm/4iATWWNVtz0ys3KnY+yfJn1O
SYTa5KIUx9Vx74sBlvn88k/DFS33GIdiLCNQaZYWtRjfotflZKDVhgXnRxMplqf1
hIQFBwatRH7I2Ht7mVkgGo8+nPdW/bLFYsdxNPaB4qdrlT8+v+jx33XgzcV+Yjw1
ozZAQHXo+nsexzNH64H7/Q==
`protect END_PROTECTED

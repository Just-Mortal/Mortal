`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lSRFwOpBS4IUBGFxH1yFl5q5ZJNDoQrmFgwfXx97eSOL7zOJL+gIcdMTq0hdG67+
UeKLtPoqj4zvW18kmKz4hhlnQE9FDPZq3q06bLqcXa/rPdn0f3eW5EiQxbL+yi7F
xQFLnmdnMV42eNU2A7hKlAwxl5YYXuBZ+3XrLck6O+K4lGCFRTYXLuCmQcPmUKfG
kr91h55QfWpvgttSjhIvtpJo4UZQJ5RRd47s41RVxkpL6AM1WnmDDB6H7086tr0p
qknjvTYcP7qIRCzpGPH/JddpsltoB9KIf6iXwoaGDglBA4oLwf59OUjDQwappbO8
Mg8UKfW2Ywd2U+LwrW2rAvnm8rDKLs9HSvwIkunGS54BiTK/XxNlbgKexerfVUw1
sDdbYsB2Qbm1k0F6JgwBQDplk+oxrcpU722ERRF/NZI0K4MH5twUlb9uVW7/O/cJ
BNJC4AO9H+r9la/PqVWRwhy6Eg8qyvBoOStzSSfzLXuJZ4xTZz+srycV3A+flNPN
QJyqt5xv4242nzUeQPVGp3+wajpCzQDN0rCpNLCY1gL/QrehU1/cZatRFlGpHdyY
JMtIEARJDTl0UXzlEfzF58Gefmiv4FjxzYfXQltTaYRDZBkXftUVb+SmZZEWnBTR
rQpKQCdDaQBPSoQc/IiNpjB6k2q+KQMjboLUdsMk+3w9XThSz5SGZ8kTjmJ5Z8Nb
C6s4u+hiT2CXqKtYgghL0BJJOnrFzU/jVXn/bAckWZbj75lwWNfXVcslSo6OLMKv
y3frEyZrn+09+PJqTzieh2zH4jFLZe+1g8J1IKzhKBi9E8o/Wl11HwrotSuGicdc
vz99vDCkELFt4XGzQHyhxF6ivxwPJ0Jz86EC6LJtNyaTE9fQ/Rcmd/uBxp5PqHnn
SEfu9YC0XE4VIdD8Ah1Xk7p8pmUI+IjyfUEGu1DVPXqqSN4sBJBBAOsnynp5Hws1
GXk4uj5qqLojASCs/DOuAkQfWgUmcn3l+aPcD28jgsfsvowIBKFAa14lPYSxzWac
M7u75WfjH8JR7l8u8dH2RCHu09UDmiG9gYxKBc72sYbd/5bHMmLQH/4sjd9s/2h5
mPoJm1pZyKxmCiHD4rfdD0azUeWyEp7g54B3YsMt/+9w+1YgZ9qymeIOlJgQtFA0
2cpRzJnrVYikFOKn8b5uzVE0h1CBB2/GyLyUVT4XoXs397TUzf1uE1s7kGI2+Ne4
Liv9F+nzEbuCLC3KhA6OSQ==
`protect END_PROTECTED

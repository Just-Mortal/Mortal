`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IfzBFS+kQs17/ZaYG0vBywSNNucC/s34RBEYirxgiy4vrclke+2HM3wXRyfI/f2e
tFwEv5WvN4Yd+96sqWP9k8pFT7CCpwDSkdcVfjEN4RSd4PLTkC+2/QjTYKsX6C1a
rEHWCWD278uqE0QlfZYGKM6Cr/MF1hrjzJZ0wAj07hXJLaWdkEBK8Z96b+hr5jIS
GtNlmeRcNEys8T776TMNMrLgCHtzhZmWFSTnZlhhOUJAO30LZPaHkEgRZqWCXPIB
yCQJh/2SrMzrH54Ld4QvdiKZPnqiM4Ct+lArMcz8OnOKN22CQCjYwz+dL3S8zSIe
aUUAN/1T/S0X748SUMV+p/CxunMfIub5l6TpJo3ElUequdRfJaoz39/Kn9gjaof9
BxwMYS9rvbgYR6CxcVFjKdoLvM8WCBXPdsz4XmpLj830Yj3bQDAP2ChLwSBmWzd2
3xwtr2yvXPRTEak9r/KO0XhuX7opWxk5xf1+YGTZbSIrayN5+wrV2HM7UudwR/So
dDdvevadyiqkSC0CNpMR2GsW9YXslSbXpIxrEAVexseTaTljTvzYUgpoSpEy6QYF
gf8xvvAilFA6VqSMv8jXGy4gcXVo2aTvsYZJL+zh6TUiyLDD2RNwkpxvpRe6op9l
551qIVr2+/sXiT3G5H06BTq97ScCLjrWjx84Jd8zQ0CkkOzrt2NSGCi6FH5Fo9Bf
C8XSbmYEIyBpnlVgmaK6U4cGYP069yXI3/kTisOVvpELwKYxC5yb3VYv/L/gXJ+j
voY24NTXD80ru32ORnVB2iWptJ52kKuAYbjUOB97zZR4OoHwkG4z4M+xjN+ABZMs
buDyrIMYCmlRM16wndg8Y2uRMVeUYebmA6jaA8vcd6LtYrcPw8+Qxx5ts0yrOrJq
t6LV3xmzoDugPKiJJVDogAbHKmdyn1YrQhZiOn6pU4/93WUBkQ8ztkWv5vBi7E4P
kX+/PSK41pAxfJR3Ex+DZ4J0qTOico+R8Wl6QWlbo/tS1Ds7ZnjjF1KM9xARlRm/
GBBt/X/PQCXyXnZYMBXO0r4Sm13VO7HhzsQ3Bca6u7r9K9XDVrxXwp8EbX40ietX
LlWEgHdriQotNWoEfP3I5JLEeFquqN8MeKhajuP2wCeNpLWxYoKDe+2QmAovi4Q/
4rh1s1HdESK7nxjq2+ZhZe4oVT1CX7uXQD+J8tB79GwDlO+cOKvCbkJYTFj4ePO1
7z3sLSQbWZejLKdfFlnTRQvyR+j91mrgZf1NBn3/Cl7Bmw4/FyP5sd9j5Z4iXxlU
+l6YhfkyuT18AWtKqMMU+sVOah7f/6DKCuMg7/9KGyFoNJI5nK9OQHyDydU4Lb7/
7jAOk1Tl73oSYGMz4ssROsUjLZWC3Fex72MKXcBXejLUp5ovJp+F1i3rQc2PbQFa
X2/2u8eo+Q+LeQsWIWjmwYh3t7xe/9f7Wij+lJxxJ1YiznzS6YekLysGkdfGA81X
soL3NKL/py5F2pJXkTVzbE3whpi0GtGPSjdp1hfmluJvEDCHZ2UK65cmCLjb7ZA0
0K03lE2+9Zu0Alzz6xwF1rgB8prwWHZKbHZO6Vun7qAB0P0xQbEn6DP48CejoFNP
nZKfYKrVQZAOWCzxA+zMhXfrzp9B0J7ydQERzN7dRA39sbMgldkTWO51sdJYo0zC
AS0y11xqNudVYJzZq8+2EfmHTlUn4QbvwYLg+Wo3kpg2GhzOxsQY1ntsgjm2VMYg
08IVICqKQprN0kwE8eepB5/EgaHxfuQHaUQAJ3ARoRjIGKBo3dbXa3U73B9a0zhm
wVoVd+ovpY8pz+ptktnyfDVpgBAL4XWgOevdv6IfdcUw7nI77sgxo9h5ED4TxhMa
UHNSMYzRXDBvYYtD4hcR1DNXGouFVDnfTh0oqCkRIvqavMoM2lLlbVTtk/RJL1tO
LyTwuRiAuDZ5M1UVJTZoYPEAvyHYwg5xVSf7i/sezBR9x28yjPQrzdCQFsYy/zeU
FxqV/t0z3gNHzhA+8mSNX97kIDyJHt1I7mfsoNWImru2/mYn3SFIsnUu6bQSiwbM
WQFGdKr//iBBm7WmQ1ocpHPz8ngzE4V26DhtiV4hPj44yiCy9EWFEmpUBcnTPQ7x
y7pboFltqFPK4Tcrw7P0n9hbZBrlixXv4vEqYrt74XSUpY3zR04oehdY/C4o60qJ
0Gm2wOVc7sLJzZuYIbULy8Hb8FY5kv8vHCaBsKinxzSrPsjVAeEtDUNu3+iY6zOk
8ln6SRUl2tGmGqagZAyL6YwK8huPBgXELNmff8bpuO03/EO2ub//4/SNlDHTk1gr
XWN4yaVZndcgr78fVfRF+7za9zEYMZz7azIvmxnpG4AgniNqPpZROfKzujCXuP9H
hG+lWeD+4ixSLIfs4qkAfJ2fOsNxLnZUkLLQahmqa40A6b0pbIh1DXTE+GKtGF5i
3vN51W25XAJKeWpc+Zmrs/49GUFJHM7acgt9BsO8CZXaItnuEt1K3jpCipRWiIfn
FxDcfraMchZledwhDc8X0TYMbpr4cXJL/EcI2tt25HdXPuGr2287Vs/10pcIGCb9
f3D5SdZB4qVbs/lc78eapXxp6zKFiTV7FkC5BbYrGkitoN2YEy1Dz1ggpfSu5V16
fKG2EoEFpa2n0kPlEZ5ZFx1fjQRhLcmKAWu9BuvmY9cdZlIbR5/or2rHceF0Mx/W
5qwjB2bqIkUWUO/DCRlmRGhtA8+EHsokOaAAwWQFkuTQOLwHwBNFU3waCwxQxltV
kRFE6nzN/TLcXu6x+F5CtxIrBLCNXgLpcessToIBRRJqB/x8aPV9rvMg7qwHcKXS
gcavtvf3gDb9zleos7OY6kF/O7KWdZ80eXQhHMBPZZ7ZIt5cidOS4YUWSkzhJi1e
bntUkHSpC56jcTvO0+AF1OP2RVaA0hwX2cMGyJrsJVPgFvsOe/gl9SAW9SJ1GyU7
5oli02o5jeOUM09ZDxqQ+rA2K/MFucNoiWB1GEjRwSYKeT74eHSceNK+U0sf9G8h
hRcNt5es6G/GnMqGvpduIMChFZQ7qAzWELwifK4Y1bum5gpaj8JPWW2rwxTFMXg1
ZVS4rBcgaTQ4gtI2wn3Vti8JXw0aBVOkPkZ3MDcFY0uABdxygOEbM/FdB3lyJ2Uy
/M8kGsWI/70tRnF5npWWn+DKI+9CW00Hq4wkwIN0Qe2VQeDu0GcQYVnVcquhSx+I
0FMoxK37vbPU87O81f5uGTm7MDF8JGHPzqiGAag5Dgfm9jtAOIqP0G1conhOMCjM
+fZq+93/aUvIbt2O4+c3xAaGHsarlRMAGlRL3mp61NfFo8XAbMV8xHMkIl1yBxjI
GP56g67PbCl+qntTtwAB+z8hOhbT0T1wujRgQ5hMp9rZgK46Fcm/grD4igmNWweB
5bOfHVZ17iCe/gumta3El4YBxJKmTm293lFtUXrY0lw1RuQ1Cb7V9zxoWC0DKldg
`protect END_PROTECTED

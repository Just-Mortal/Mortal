`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LXG4aMyUFVhPUBmkGi+Gzi7cdStf9tIwswaXuXBECI/FmZOGW7UWmt75YauD7KTW
dA9rZLE7SD19Y/J/XgmI0R0cjHsff7Ghd1LOVawYFCFdKoh5cN1UqHd7OIDp11j0
+4ElDIQ38RlDZNauf+r7wINJKL/XQdDW7gJ6eQvjacmjhfy2rNJaK6vJ/QRhJJtg
quLdM+d2FPNp+5ajFOYS84efiIl9UdkKNJeLeThKoznknEb5RAIbUrscCMtBcMGI
4/TBHdUJ/243qSXY8Xt0a0LUsUaoewjri/HGgV1pkakN4U3k7Ok5/tpusU6Zfe5F
ZsYWWx+9xaH18GMtmpDGP1KN97yWJrdIurmO9V8d0BHsXil/OpSS9MQxdtTqWOxV
/H6iEGqjXMsfuYkOPx7R61W9pUdVZkJbRdGaMsYMY9NCQB8r+zypHNRSfet/HpLf
Khx/YnzDlLW5pnRd7SQ6a/YILcW7NLqbG8O+4o9pTLyq0Q1u/6Ah5IVP4D6pGCrI
AhmseyAJw+8zUQJeE9qGdOg+BcGjjoVAyR2RCDlzE0lg/hvWs4bum90fzwFzHdGD
X+NHOgCg2HJAPzrxxlQQN7Jr070r6uEztbSqSzoJf1X6xok1537g7mZwuasqjPFW
gWS/LaJA+D4f5pMUd4abKHewh3Uov9UTjFAo5O+HDCgYwDAKOkWf1fcrpUDsDr4Y
R1oI7C18bfbOAbV1GqfNZ1HF9T8y651+F9AcN4ffZk3ELtciTz/5sKXv4vuRmbPL
bF4LnBNTeHDxFu9fkatC0QrCqSBoRBzEzDvtmGNhyMD85wSseXpekIXXNP6Tzycm
QeTkk06IwxyuOITst1qSQLzF+YMCWM9yE06JC+VxqifLRwYHCF9VdBj5VwpfyYw9
K2evPnrWYhsIpCWuwZL4EYW3E6zrFP5UQQob7K36lRg5980dfC+R0foYp0hJy+Y/
1NVvDYEPyZFZCi16VptpiRg6yM33c+WTBNi7z74NuFYYQKvGGorGZp52H7iSkQYR
5kR23UPkCDbEBsic6VaNiieVXiLl8D32tipnT0Cu/Jm/Mqu2Dlqp5+MkFcBbnclv
wVPEjh5jUmVFpHpu4p93wBI6MCTnt5yN6xj0asqjcetRFkn7kWDHhVkWKj3TPIdM
3jm1aKKKBSaUCGHQ3kck6W8NM53WQ/LCxkqvgJsp48rjgEa8jutJw273U/QD4A5o
x6HafkWyfLNC/DYDxFoo+n0y57l3ecIhT5U5fc4dSVMMnT51yOXCYnzvY8fdjOU8
Z2UoH+4DWTxlxw6ANAkT70yFrdt7spvaogYmcf6gT6EKS/Aaonqy0t6llwe2Lwga
a0L7se/UNqr81o7ifkaBVJPxXdKeZlBBhZ3regYiANVILdPW5auZidk6mXhuhJsw
PJoXmLQMBYji1RP+owQKlt0Ie99XVkfPNZoZ9OB0U09BQCoW5KZYfF/ePpGydtKW
v2EKDxzVNfV7RBFmuMcFXt5U5ewHBlCxzrLrniC0SNFHEvWgvLbeMnn2wUxaLaso
5ymSBfnj1iMgxPX4MssBL00tofCuJ7B7vzhqqr4Ou3fPvmA3el8FgSI7WjsSh8Gp
3aICtJe8tDIagXXcEPiAxpA+utMZJdt3OE5tzWmXyQ45Tkd4GGb1hGq4wNInFBWw
UrmpMto1rdTz01WwvnzzpIoyre/cnbY0+E0Emjlqvb1aUKuyVkAdvsMOxGpQgwG1
+OJf/xPjXlAJ3vczYcLlN4DMS8ekdMXH3oP54faE/s3PDgVU4PLMOQ3lTWBnTV5W
Jbpd08DdgHZVTb0CRP8FQWra3QmcMaP4J7qPiZDDzQZgwjMvilwjo7W3ruYT62fK
jOrkw3lNjKAAB733LT2URHop5iYfy9GdWqXcSr/BGkeuo03TIiQGmgttKczw7X+N
nlsVSFZpjhrShqcwr3RvITriLGAsAtl2OoFfZoKId1us8m+Ajv45OcvkJINpGF4H
ZB1w5VNxBtYjirkPY1dRUUdci+kp8mgo5JpHRSAdd/ayCsbeBXGhbyMRUVbqLGcr
PSMwAJIuwCwhzQsQhbKzcEVj2KjKsDuDtdDzUqRuziwQAP0pAg7bDUhD/eN9LBZA
zHvHkYKpQiusxop0edYxWWlDpCA2V8bsTHwQD1mqd1v7YaYm+0PmupR2ObSiBrZn
XKp+RySDiESOESCecvHCPI3tLvAPVk7tlpj/1RihhF+R/iDunZGGc9o1ryPyva+C
soKKs+Nl0XkyF+IyVnzc9NxO8Yus9KWV882TT40Rz6Uli2VNHm0JSVBleZNI5xhU
FIdv9pUp5BdMKAbBu/aO+vvzV9CsNpLlxV1X8VTuVZ9OTp6SvuCAFA7BDh1j+aKL
IUaKg3d+I3aP1GC/UuZP6t5zBa/f7FCxyc58IkY5wRHzOETSe73MgPXa5i6RyDAB
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1JTT4svKmm3cOTCXBJ/KOnkQbQdkTHC5sRCWVWjylnARCPIjmLcwgBoB0dZSKym
P9XXXUhXggutZPsFENxVaNn5Ump1X6z0Dxnpq5i2osyQNdLvbw6eNleo7viXM0xe
ylVRmPqwIZgDcqWyv2QgpmjcW5OFK/cu/GY6c97Uf1GUlpF+HLIWx53r0sN0k/rn
HAJl149DbRvK23PHtsCkGNyE7OK9fghHKbKj79NIeQkM4iuN4iNq6hLzriiYrtyo
C4iSXXgTKgE7mo8GXA+o2mgE80weEc4OMr49izORQoyC8cs+lx8EYB67qPhmhl5i
w1FJimhbJ1WNMcc6/Azo0ODpPNsBt4JSZiCAMUqy25VRCMCcRQdzzNYID4b1jK1z
LIVED+179hpROEAFv06qqhgfh+QxKwWHjU7jNeF8lTsyzqj+y18MWfvwyeudbM9Z
E6M2HrSHFCNC35HDKdxTpPqmcv577SQ4WjYoJ7yzHbmHbgnwfGE3YPhn3fZ+jR2h
ppg/4yN0wPHZRnLQE7rQzTrK2gpWt3VIzszY9JmNYpBoKaW2SUnQbPmm3hsNze/9
ICDUVDrEZFPreJjxS9q2ZDH+mwE6uwvCJws8gbvTU24KGZX0bU8wpq4nysaTS7+A
tARAuy/JhcvP29GZ/tGqdmRRRiu9guHYx184IiNMPAmUPWyCroYrR3nTuVPab5Ab
FO/yHzDgNUIWjn7NrTe2lHVR6ut/h970zkV7wx7RCEL0kuCJ8rQbNBdh6OxEve4G
3AD9gbKOpIozEWGobucwE+13K1FD0CzqmsJd1QRQHktmlSHqdAo6Y2ySG6SUpDnI
Ea9icwD5YsLz+DIuZh04zvIDQ+dpL3oe1MCZDdk8YeEEBP+/hCrzdGMF7+C6Wixm
wGChzkeXedU4A+PvcEQbvt+NRC12WVqXLhpkw47xVFRhFWLvfrMQOiewGp8Z+EaF
p2vhLkB2H/+LyFa/+lLgfIJrtCZhLf7xuy7l6tF6yfXiUqkCK2TFEg53MUAMLCMb
xt2AqkXmBegaKq/JOFncmq+buraTL5g3y/wbVtDdcl1WzpNgUxQVTtQvZ+jspMUi
F8AteAfTVoCYFmeehvoebWOvLEMOLkHkIsf10RBLrZ5Cv1Fi6+b4mjm5uCqZ/+as
MEJ6VJrHAy2zaOLPHtDeBifAoewzUnFwU8EztqxbYqG520+tmvaA5cSX+og19pxR
ipMFoF8D/BR6RD6jxfrHuhJOAirYbHlyryPPp5zRLzDmmsMmVj52EGkk3JjpJd1w
d+tMDO6Bb97AZehJh+VKWqkdEZE8xMf3/HRbnnUB8F9RrZf/dm7sgvGc1cM8v77n
lhOsKUmcK5HZ0l7+F2EKcncH6Yp/94+99BH2/h++g4BVzbWIB2+ncb9ajUy/rDTh
0AGlYiSPzJn6B70yD3xLiXqrgHYpqVHpDmLYsZBI3GrMBWAcsAure7AyzadUmG+z
gaaWFFME1vszWn8fvqZS2bB8Se16XI2BE620IGHNRd5Ye1xhtMRe47RdyYoeV0pZ
9ywfI6ijAZ8tRXHUllIBC/71g7pFyiDDwGUcOjk1gBK/MlXFFC2sRwT7vUioMFV3
YAJWLy9a8sla2hHBSL7C1tmb4Akgfbos1q+/+p1hdq4oEUlPvIR62d0aHTXj/wl0
n6iYDdFW2fbdF2eZWyjCw0pGEpZxA8xQ/tq4JkixaBtC+Zmi+py3RrT5r6dICDao
2FtdT6vc5TMAP4fXxmqTT3Gck36MwbTumRclBmi3XGYmNV04E7GNzI6L5sZ9lx89
hsCRC1tu80XpVJxoaTRYpbKjwpgJUrRIdmFbrU5aMwrOJw3J9SwRAmS6E5odfxWH
0O6Pbt5fbUA6RSmU+a/qjQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/JiF+kcr3RxR35jFnhUk+ZGNzNLM6ep/asFjdVKtUrtV8aj83ChWwhXmDdH2IsG
tzLOYae+iG2aeFxf6rqJTcJM9t84jYCkSjIBo9oTWtCga+y5B/abS8YU05NeQ0qb
eaEEmkOmFDoYQy1ccY3eHMGpeniT1AhTqGx9dhI6fzBy3FwBfMJJKXjR2u0Z3kXY
kskliqWZRvcDmZiQ8cBJzRepJR2OJ1Cx2WOEkQ4vlpYEFDlVEKZ2JYuaBP5RMj6E
e4IUCUZ+Iy91T3dtNLbg1QgC+oNpiS7QeH7A6Cso4ZoMf9xOuK9pMd3VQl30WskX
TX2HQYK7zYEqzmWyVklVhMsWT1UTXDlD4fbJWq0g3ao838nynyc2uwZdl3lLmYKK
mkrG9pgf5VbDFi5t/W7sRSJlFH8Z+kpiR4Lrc0M6SVvORPdNvUW0RGbamUmPfZSI
0hNGKFzc+ooNr3mRHmZDg6lzPf8EVJp7gsjmGFRDYmN69/naVXA7afd79d33P25m
xexpKajEPQCOfHN3xaesxFL6y30KnwcSIozlcO5yrZ4NUpmespvyUEk/IQ93eaSV
EFKkUh2mhf4kPa2WMhtNJA==
`protect END_PROTECTED

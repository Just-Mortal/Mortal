`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ySn/k9CfgqrVlvO7WmvTnjGHb4ULWwFUU4vf3I+7r4SByUaHkL0rMjY6hRtJuzGJ
qZeCvAKRQDsDxngKJcUND2L9ixtfZ9mV/DMM2oUUnZsjHaAzBnf0ANCzFg35RemA
IzgTASlZyto7BpHqwWFS+6JnHzdZuRnLaBYFzQVzGdaaaccWcwguu0Lsu/6HU2pk
LSAsZt7GET/F+Uw6rEiKrhk6nFp5AqcwrIlFXyuqmxd5qAzIOXyrvAe3PAqzHJFq
gVpF931sXuW6CkBA+WDu0OVizWmbE+fyntE3xZxnAv0MyfHji1hEzLp13X5Yh0FB
WHy6LELAVFreKW/lIgBg16yQrAY1aseZQci2Vn7GWhTKPn4naCQqj7KNXhxPpJnV
NHSP/MbxON6hRZhybp2+SJRlvyl7Bel2zlU8CmyNdY94OZbGivSrPVTGUpHbwiBx
kDW0hNEZuszGNL4TH2VO8rYUBfZluXqy8unELyPuINmYAB/nZKik6Il4UujfRqWE
/9kHLevp/iKjjJzauNO6dFmLTS7nRo8FInY24q+raYKI8OjKB/60P7OYajsR0THy
vSKqgRIboZTzY53SxFScE5y888XPjKt1bART9TSddcA4pOTe+lshf3ZNC3sakuGb
kM2Zo2H6SgudEb4VS/BEV1plqQ3d2LGhsMUutjKhGWDFjLQtp+Tg3kxhqFPf/JRM
oaafrdFkFo83TJvYYf2gmettUbAoAXdFNBPyr6KmNdZRek+NzW1mThovYm9VBDMh
MFz+M8nI1BRTk+4Or+JE0aRREJHiyjgnaSQuAhTnCfM0oN0OKGWxFgFr194+htxQ
opJk2clbJiEIMpLFhMgxeNIwpxjBdSIBuur2xCfZ5UEWct2uCmcnm8WIBOPUZwb/
6Z2QvrnSOIXS+CDN3gU7aJtkqF+EesPmGv1wVG/k8DKtAsr4nFxxRTIuTbK/iU4Y
Cw/RqnAiqCEysz4Lkw/clnJnPH3Ejaw8NqeEMJ2pTl6HewqwVPy1Zc+8hb4bvgXF
uVts5d8ncoW0HjVjxJp6WeqMNn/ZQ/a3OjgEH9HhiZOGRc+hnojnOzg2Xgdf3Dgi
+SjzoBpnvChldsSYREkKTDJDKqnBX3Ez/gmTe6bGkk1Kph0DpywuM3JQZ5AzRniw
xfX5TjPt+SgyfVtpCqob37uALvzYf60XGY5Q4BbYLvh9mXPkSHKiM31w7JbTzuP/
4QksKfLf/8K/9svwO0uCXxWbUdM72dalTSo8AFd+zk9rd/pQNWFFaLhNca7Wohdo
rtN0voGyY0+lIOqFKsaH5IKY13owC4B9157uqlHuDpgXhmF9RUhHZPxwa4k5RmyB
QiAGLZRXtXjgBNXNpp1ReeniDW/8+LRF2Obq7rCi9VV9QJsxpRjqtVy7rss9fnDr
jky+ZOrPQ2h+wCVlPXdwJfpFfP3HiSuaQ7OXD4NWcBtEVP1F1IYShR5qTTmCJe+D
IFO13pZBbl34YBUdSEgTc+yaUEgJrzG6DHoRbTEpRUFDp1BYOwNFzfCdtMZb6zEV
CAn6/XNpjV/o6YSfo4C0WZxWTKtjwwOsalsKzFU4icVGuQ0Kczxie4b59Pm+8Qtg
pS1pfRwxP4Qq+t9S/Vwhj0xInGPQLzGmAqj2z2F93nFNA0Fq3iobtyMGDPhUB5++
KgM8qVlF6RUqEIffZMF4dY9ygkSIMRO0uheoSAU32C3FmtCvU9WoDoNU+rMIEAW4
iKtICiNjmenNt725VDEaS3uJ7wcadBBkkvKN5+JSZPfBeQBwm+cSXW+NksDIZ6ZN
po1kL3j5x5U22ZjcdTlW4aC1Ao0BLyy+bsJwZU4+gWxkfEC33ks8OiFjz3e/Fgym
0fdB6eexyaFcpthHzpKrtxLLwmGq8770l+7c2Khd6aD+0akTNbGBgIwrWeRDDV7Y
WeOSFagYA9XgvlU8uYkUpquoc7dEIVcodQKpnYUJ2T704YUUdOZZvbU9f+K27WxI
HikiMvlMM5U0w2mwulUnt2p1ZFb7ePeha90SnSLr96mKR7fHtCk5GFiXNfS2bBrK
k8CU/BfkdI7vQiqCZOQIPYtQ+3ngO7Vq8mwmPgGQyrP/ixhX2Q/wyIQy097pyMUZ
6dIwTD6w5xy0t2ylieain/ozHBclzBWai9wcjY/RoWWQeCC5ikAcojyk/mCPsiuG
RWv+Ppkp9DPaZzUyBUn6YCTwwNts/4Dl5iDg6THipsbQ5UJrsVTwPWyfT0jOL9y8
yqQ6aib6CXbCWS5UInEltWfcgZi5NZKRkqcXP5m5SrtLw4TS3DWrCG7FcHAfvC0y
Z5czFtIHYDuIvVzUW/pj9ozu4dRqDhzEhHwD6WKrAsezdfuAuVuMJ0TB138Bk+bf
SX41qC7hMkfu2GlSrrn0Vm8mRY3r0VUeJIF8E/cNbYSJbObTWfVjdKS3iUjQJlIj
99gcoKCso3lQtggS9nxu9RhaGtp5U9TEcPHyb/jOu1+6Xn1UyscR0WwHmc2xYN3A
mS5BxlhvRBBcCttLtypVV5UduNTGcPrtKJ1T1a3g3sB1gm5TCUZJzxP5OJ1fm2di
Q7lbgmbGMx+J96keEoRlbaJbC/Aw2lOvCdb/cW9/IghxbH34cXzWPkLyUD0dkXes
65mnbNODgVgfGppHdPIKN6ZpbEC6J8Eh6jhZPs3A9iiUPwJ0S+f2W2+ryFhLFUs+
WFHIOPXrXU/Ltk4A1t6EsD+B+QfJPdP8D2vv9vxPZ1f1NPW9rG7ROt0/FQa9Esbt
IMbCLmSQn4JJY/zqLNwRIb9o/rogN9yTiVoIcObFsC3FDTfRcaztM2Khmvp6g4CG
SfER4i2WwgaAuaut6kO1RzO+Y1mWdobHotOwxA3odp8Rxh2W30qZz/MRsmiXc7U1
Hw9VA28/yfqMmEU8LbcqJAQK1yyKjd4pnmujFDkVwHbZOE1DLoJzqj2bVyO3RVvs
eqhb+ezFyL2/sWlHU2oW78DeGXR2PdDrCQ4KsU+ee5YqI480Qoaq756sA0t1ymtP
NVmQ+jcpffXh6uFOZuRN2fI4H0Jfgq11uvijji47hPhLkmc/xGMAjg3urPiImc5g
/NTrv+49FpdivvlRAFd0jhc1cVIhC8t4kCmjTEx9zOovWLzcUopwmQBeh0ppg+pa
RzWVoh7HKEqI14N4OVIIqEX+UyOqm11pjAzvIt+45pahb5xEGS0IompcZrj/EZwD
JX420wLxClvY1SdH9xdqqnzY40wKYGRD46igNw8s/uifWTxovO/6nGRLFOjFABpN
l0U3QMIT5Dq6paYl+kv+fOtdykzyeQ+0yRzcd0yl686xdNEUrcoDk7ZvfzCUQcZc
5hczn6LjtB1tFgQDfaNAKTqNe9Jn4c4NaVoPcTsHFD7Y+lhqDqIbAsmH8Gra+RGH
8+pqss0MjlyN7LjzNesg3IqtfWkH7R+ihZuHA3wuMQvMwy4emRwbpgR2c0C2cg0e
rBL4U4BjFvTgNcjOISgiSs4s1txhxtA5HN0urXgT7KHWxHvmiAqPbqse6Fkkhm9H
mKKtsbO/0mHOG46eWWb4hz8VYczE6h9I8bPvGCwo4I4QADuKZMvCQqBEif0QayJn
/wF5gXiFhER0MTQbLuphYeeObL+OCaZ79VH/FY6OdUjR0hubxFkvlAda6xLWzv21
au2DFaUg73fJpJN6sDjPFncI3wb0Vm3Imq4kmJywZvGyFfd/Qu/fm7xo3cmhmsa6
mVUQb5x558KYPmJ6uP9uETKUFHgXQX2YDT4QxSyh9sSg4KMEEtTWNP7qRwj6x5HL
C+ljo5SeUojj1hmbhG2SWKpOLJ1lAwoTG6ghjf7swHFSvRsASsTVvzhdRHQVXm5y
2Ej6QySLp/Egq+z2wCwJThvzIhZyTtkSxggHtrM0m74WHFiZnhwC3SDjWSN2tZDg
8or81f53bgUTmowpM9GT/dCPpIQG3HASr3tFlUMUo6Pg4peIvKIFR9dua4qG84j4
SqEZ0KsxRxmMUJ4C1SgxDcfAEIHjyUnOdRj8jwO0mv4NcI1468wFPchm0v981H/Y
wY0YzfLYQhQFJcobaL+//Zmz5jatQb2tn9XlmkKGELOwmPgoxc1jGlwtk1dcKGPz
m7t11MDAKW/dTb1eMSk4NHr1pFATLMVg6yD4yn74D2hYbN4kX5mEsQ2zuNo0c3o3
T8TEJi7aWTadC5PkRlJmPQGJtCEyhFLj+JSbvZD2e7coHhhrQnYYvysxrY7cDoxs
mPySuEvjBDR3IHutiu9jZgfNLmL0EQ4CUBfnk/4WZufFCoU8OcfUXXMl8SgwTZw+
/wThTW0J8sV5vOwuF9ggrEocv2+etc84p21UaWxg/J932A3cHn1uT3/dE5qjActI
M7j6rwMXz5aujm7UlPFx6k0vy/DazwhUmYeAQfuxZk3JXPGPX5XuNBK0lLA+KZTR
HvuGoewpt6AAndAZCjECXjT12mVUZ9uPeTkTvM7xD5X8axV+HSJY8HLPBGVKgESd
XbT9hTnfEfrOlWMp4UVGWvBye+mCwujgoIcqt1dMbT45oJfUWR0X9w3O1ej0KtZC
L0valTXgFn2U7785ftDxxavqmsEYK+13MuDfMQlUyAj6T50xc8ETqvWQCLcXF6zz
pe014LhjIkCkQSxDm0/ap1vKmbDnTH7n6LZ2JQhCttZOoh9hr0oLlpP7RbJzskvB
Wt0jrGKpNj86+270ye9vcwsXVz4xQ9KBiMDx0yqsSPS2shEq0FfBksZdB4A0bPDH
STXqrhnZATpnNdb0qpYj/E1aG7PrqSFk0jPq+G8RGyVCOqGiS/YSI24VML0WJv9w
FoO1QU5Rt4i28gzyD1v9tDVje7sSB990wstgm+BetWRTIN+uYTSUZlSRGLJJz5RX
K9wiCqZbqWhk36VPFS0dJn5JsqUaGawx4VvwOQKo0af2up7HhWX1SsQLiGV5jpx9
N1Z8OJFqua3amUojr2YDkcCuRSXnHE2CrJHlN6VlW14JujzgHlAJW3UxeKW6C/mF
39zizHFsqOirQeO5Ohf2cRxSspKmkw6TmgH/oWmC/mn1yBU/hEX3r9K40MYxSHPi
GteoLZEf5QizFVOGYl8mXci/RFTHU/Dci16qUjtZ139INHJIFH5KTYHiFe9KuQkb
fgU+LPC0CozkJ9yOzKADDwpcaa6/SBb4GbseiwAelciUhkvn4ZgWXWgSKIHJXLxW
oxY6ZyAE3AL5lJtvo276murn4Z3/ed6/7gcv7BJ9pJPgFFjJIQji7uPH/Odnt4u5
MCGNglBUKB6j8l3T579ZnAg1nhhLoyCU6BsKWbsgDTPNIiQX2XvqH9wG5gbSGqE9
w7SpH+iIvoUJthuXLQKuwDNbIO9GOKvPjdAP1VG8f5HRPa+7GaAXxVt3kQMLO7hq
0fJAkM9Ykz9pYsVpB2kVWyK8200pWnFD/RGBo96IcTOWkZb73SBIcPFgb0dkd5pN
Jrun4wEsJn5G6de7KbEn+FaWK3hYGUaPUfBZIDpEBCkNfzWu8wxsSHQij7kO9ikQ
Er7ylardHiJAKmHWc/yLHxiYXr/yr/Q7Xybh1DBIPofSQY1+PI4DNZPSz0Czt8Q0
obVYnXjAm2erIaP3Nl9rIJFMryx+ztUq7z7tLUullIfmuhWxU7rcpZhZ9bpvWzHz
lEFDK2ozwpC0G4KYC0hItVNRXuU2zXwg0qOP9WEy9wwQyfX4vEphtY9sQQmMs8bo
cnAP0Ws+kESyv5q+H5JY/PjzTk+FETO7mtSIN7o+7uqpXk052mVQeMcOPYaW+4zr
tJ1J3s2M/mG63Dt1XWLGNACzVP7StpmrgFkFKdwVrZM1lJPwW3LcAdwvUow3I8+C
/GnCjpTCclu7woB0EGe1hwtZRFp1ke2SWCJkCI1aNOuxBM85XUwz9P1FtqgZ1wMM
xrRGCBjjIYDbDTRFye1pysa6WBW+4G8mZDi9lBukyPqbUPVMM2hdO9ycPfzR/RYt
YKg8dgYRf3X9ql+aUudTIGJaVT6fefhOodCeBvrFBtUa0gb2SBSQIBwLYbzTRP7z
qLlAo42zKFmryr5mZQ8YYalwR1uKzeLW1Y2wm+7aKXP71iVpwwn0wUEVqVl+9LbX
94SRqNQoEy9gGaCzqArvpodpvgP/K/gZUroG5D5JL7rsVORVBARaIpXiSEU0hOMA
gEQq1NKaK+dl9qCr71bDh3KHWGJ7m3Vuj/fBoZECM4EbjZYxMpVtTgZeXLqjod3m
9CJnDz1/pIEVc5rISxWqjrWHt7wzx2meIZ6dmbdTJkAnVM/NKNEqgxKwYNW6gAow
A4dnGP4yHTVid50bZZJhzb9BuD0GVYvEPtghlxHAdmPU7F4bCQ2vys1XRn+xb87j
Es3xQLCkoyIV5J1RFdUQvkEkx1t+n5goe9zNQRv8Tnua7wvgk0f/auUBW6vsR8js
nnDaJZpJcO6tt92pVfAREtN5DTrDiloatdLmC/dfCM0FIkEf692uVyfaGIqNhQeR
IQ2nZ4SQ1ePGmnMANzQttV6BrIuSX6xVtnc5CpanBgpLjsOxy4MkMdE7FlxgXvXy
CAd43AirrZjtwiqDI2/Dk7vR7zpTc48+oa3N25lWbKZVr4VSAYlIaiDb/2ec9nGP
+Q94yXHQO2XsraJqNrXrHavrrDqlKCmSbMdLd04avF08dQG0aI8ewKfkQZflP9EV
O6s+9e2Spt3XD4ScVIewoE1V59PqZzsYurbF6QqahN6qH0SJuw9wcVGoHFWaxsJI
NwSkr/jPGBxk+eJDQpJmW8WuIHxlnhrjN1Jn+hOc+321g80Wdzk1ZXesR7TKhscF
WbsLUNbeCBRREFAB34gkCX28+D9RQ9LmUxPaAoBfwCZnLLqJGJU0jPZIQOm4FTDu
MYZmPf+OcObLRfyDy62DWeGv9Mb40GRGZV72uqVhypZykS7oE5RdyC3ASAzviNVi
6RQg3+WRvFyAgT0XiyD22SkcOrwADaTYPC8vN4PVtOxtaTg2Gk3nez1/CnvN11ae
S8yXGtiozj45z6d8CHyJaeFO0IkOpE0VuxjxVEdA19/rdp9k7qZV8q2sreIglJwK
KamTB9huTeVetajM+f0gSgvkKuGCaLJ3j026qmyOZiUpc3ocpNM6uhsPROOsVyMm
GEZusCYYBU/9zhwH6G3RXHCkoMmseXkmiRtTDuUxP5p1CSQQ/6t5nZL/FXzmbaN0
KTNhvqPg8v44+6z2kqCl5ugLTfxwjgAfHCS9Fg+Pkg3wGcC04CSyz4pypWIGo4Zd
VVR6jOb+aTQvRRdqvKZG4C5Xi01tfdbK1jrLOtE71T0yemqD5U04vfLTmIiekWC6
vX/6moL5stz6UG6lYw6XiqU5QcA4oe+toVJbXqRxJ/kNUQ4YvLDmawQTgaTHi5bH
vFmfnU/XiBbHBTqWMXqvKMPcKEHqm6BgBu9+bIljdSq5OXREqpRJrWAUWgAPK6ur
HLQKrbw+FqgTsWGlEpPidyURq3NR5/nOELtiQP5/ciMiiWoPlqBwptts1ogJpvZ8
DXboDp3QlVyzMNL0HMzehhaOIa7u0qBlwLtmSnpHfFc7jUBO8wA8kbaiG6kfZ9KP
HHcABCmcU+ELcTJNMYUNe40rmpWVJSjuxgbIRNpfjC8WQCW6YoAtfYqPcJFGvk6d
u6hZfoQOBWC8YmLPc3Rmi/5OajD8PkNwYeNCjnse475v6xm+kZfEebZZyzxofNdW
CyjIl80iMZdB2Qc1vkP48x68VDUzAq/BJ/x0pKFFMwFMJnCP+pyxoEP03RMbOJ5n
kQeN1wVU85IKBcpsBV+xTemqIMoNPTrqjuws+qd9izAaUHQe/QR9rXJhDzgyUPOQ
4pj66dy5TqSWhn4bGAFnQcOpelhpcfToXCpSSZ5DejFJGT/aGlnDox7wtNcbNHf+
+mMNopoL6Z+6gVe16pcVmecPBrGnoIvka7JDuT29Cy5db2LpejJVTXk+l/7O5Tr/
eN1xtZAWsCAml2Mwsnc0L2UcZz9k36uD6Q0y0dh99Kf0/tbJk1YHLzqdRIRPJ39S
TI5TDkBYg1MwoDx5kUNluq3xGkS33MLK3Pj8o09uDn3MYK76ALnDL0Ve2ug512hg
zaRivL4EnFYrOA9/Nyy2k7z9t7jGIp5FwrxZFu8uiXrVO0bXTPzwr59JiuzfFefH
PdFqezxUna3Z2Lg44vZwz4DXQjNti5r/iJXThsL3tgVA0Cl6sl0X1TeG6X+83q7H
oOXL/wiZJSFbj+UkgOa1TzKW3qrAu2SVnzXBHHOuF8R5iHZhOQKBrDc1NEDU3Ocm
gpp0POrmS/vlXZ7R/fbQkfdflFti4Rn1IJgRjyOYPif0rUIYjqKFtr29wokqpUa5
6XLBcVv98vy4FtU8caYphHMcSMBKD+ViVtef4CMNDs5WhIKaDiFQSjTcZ6tZWGcL
S54DVnW2GT9cYXOm9yfimZhvoYO7arncMC9lmL3OpBBi2asXSgSghB6JtTO3AR66
6HcmnqtwCKmSmHfoUXlhBDr5sYPHPzNE4JL7t17XhCKUo6+6y0W5hNJpFg130zbT
OmCFX/QqEdBwKOy4MJYXHdxFRqGpLsuwv9Zka3/LAM8vwGeTFENo1refKZK4cltR
bYggZ2tz7BRQdmzJP/dmVpi4VOoiNYtBc84aLNLJDNKLg4AbLO6I0iEo6p9XCr67
eab4Z3z1Mg3bIbqA5bOTPp40vlM6q48HwGIAKqqSK6j1so1hUrWVgnxMm6HrsJJM
bMcohpSgNGQZoFchKUrLL+7W9PyCNXTQKMrdcQa0ZyOpeaZUxB///1Qhw0cOoECW
IZm1HvoaxoJb0XPj9XcT9wE6Zh4IW6Us7ns4V8Dmct6OxOc0Ob5HKbrW7BRPSgSo
2qaojqk+kfEZrty8qypNIPPCobbjjGCwVLUMXgXCUqvrOs0RHbYHsw9I4g7T6caa
DZcLHxrl8xqBYf7e6rLyiYb8Ih8xiEpa5wMEuVSBphNigsPHyeHqiIfC/oXvm1Cq
m/7Ci2rxecoS1De7Sc3mzyKdF0nPbvVA+/tSBEbQi8rH/CHrZJviMS9X7THGA/Oa
GNCtuKNT0yNVwhS+VLKbxQBGdKI6Ok3HSsBSaoQDrTxLoaSAzT9JNJLrNi8M9bBz
ogvUv0D6o81LgXec1P972GIH2WCIz7v9ct1DhZ9UG1ohgUaPY6ZIZJO4oppHvsLA
ir3VeI/G2S6AljTPzPvo86YR5cDO4PN32YNwSqYoRhRLAdK52x9fbaU+vWpkScQl
P+ySF2GDF2qUIae3TMsY8Q87KTi6Bfy/ERnrGMz/h9JkugA2zB6Z7oPOVvYpbG2E
PYpMxelZFQ5iPsCEvG920eGzDBYEbciM+tgn3EajS9VcHPS85g0QFT0colExDx4w
HWpdPhfyRCz16ksDl2upQej3nZXajiUxxDwPYp4lsjafZfoacmsX+xNJ98Vr5rh5
tIpGc6qsAkWKZsVNIo6ByGc2iH2Olc+dZim5oOKDx97dJjzz5PkhrlsifWbkXYxn
uCS1oDh6Yak5g/q/B6BsXJ10NAe5tJfKQJwSNMUQ0j/uv5jDH+a1EyIhbYQ2chOf
FPgMLErHhELPaRIqB+39zeIA5fV/kuqsgULwhEbCvEqpFTLXWmSMchnkGK5myfP8
E8jA1bloAKOA9+zV7jurZ2JysHmbg3gyetS09aHvmCQyugNFq0Woyk4R00bxIYfq
5bZc2eLyQH0OldEZ4+ecTVOBaxkQM3dFUImLxDSD5Ar9T7K710O7skw3K2UE+7S0
pY2VIPX1pztgvNLXJzoUKAewiar2am6qLeUp3d7dvv/bWiQf4397sncOu4ngDaD8
VjZjPsTs4iJdQH2Ky0EyifIV9jc3hnZ9e8Hbe5v2UcccjWMWDBALEwTBVuJn7OvP
zBY2WC6847stG4IALeczOnDjfx2SNc4O8qK3KJvWJZqjllcZNYW/THMy2QoNVvCq
PQBgYp68WIZuvo+qZnMX6lqhoMRtWGQfiHBv8rSdNRiCSe0T3UAEyoITqUTtLIvy
pHWeZQOmTLl1g8jS+Mu1SONjlJ0iRWRlssK9rxjgmToMvXSNR8+ekOV/33Rl5Kp6
HfESNHYq+gNeUpD0atTqvJJGWk1T9aVLPpJhWDL78pX81wExzeRo/oaagex+1Fse
enP916RgctlioXaDRr3r7VnOyn0tR8VfriooLoIuWqVQSuRqHDCYWBiq6qy3O7C1
pX1G0Xxpx/dfq1NFv30cVP6BVxzE2Qf7HaTa024LrdUY6/HYErzKkKV3sETqsiB1
QbbTj3q4pelLS5O3shryLww3/Bq9zsFl44zCggsVKx9+fL3MnxDjMGn8xUPUlZ78
mP4OHMCHkBczl7Nu9qToy95nV4ZHLrqRtb4LcGrSAXbHM/edqpjumEawDKAt7Szw
v7zEqa+rsZrXWH4TPTo6uJlKcK5uM6dL/zS1I3mrPxoU39rDx/h3NbVqsWfYJxoJ
BR56nXu6uDPpMkF85xCx3qfykPwiWdxxtCD5hiZIyel3RwOq5tsczrqy/CtGQNYg
W9AODoxSMzhI/ROP+edLUMpL6hI0Py0NST6zthYWWY6baG1pEOw+hZPG9VFWAKMq
aLNadnsoiVsVm3EZSd1tGC19cXatAk61p3o0Re34Gn8vHA3bqfqIdvs9wHph5mcY
8sfnIdkx8CvP6awmgLW78u73AFh5avwblTYOqD1CPS1Vto79VSUpnOKPqimIaGM3
rUBFaGjQMGFjJcoPZQbXGEPHe5YjE4MVXV5v7Ia0Zxi2o0Z6bzLr7S4AcFkgAS9g
Q4E/7FzLz+xr4tZBLUc8duxHCN+hN0j9Ev14jEegDmA+WNTgzcOGQo/EKlzHSwdX
OB0Km26V+6Z/7fmsKTW8S4IqQlR4nsP/I3/ren+bxlokKsFFAoPoz4gYotgwY/Ko
45aKH2IfRKIkHF+kpPeBnK2dsdKj63m/1Pgf7OW8RtaqKY+DeDHvv2gI0JmYEoMz
qS8iEiNBKH+EoHXD4pljxD7puMFLvm026E0nw14MNJqsqkNKnOIbnPe6QRGfK9aw
/cA6mBXz8gTSc0TBkxdotIoD593qL8rTVP6b6StCPuQufqiDu1Vz+NO3sP21kZMD
NqrMmcHXOnQBrx0Z4vDI5f8qY9m/l84GBFprLhkj1mmujp8cloRxTi69xgXBMeWG
K/EGbF0UvmUJmvf5foipS4T1g5n+2CvEsBoePc+QMMHYZZjG8LXDnMlwVhYjXOdi
SA/sBLJRgPNS3tz0IX//zK/K8Iijsg/sfLjc3Gjl5zF5WEnuEpEmNq8OPzHHV7C8
owJsac2LMg6/i2STXnRlygpEKyhfEDtOgFLv5M22oZ/gvX11dscDEjbXJL0gVX/C
GpfP1wfX1cTBgVY/UqiqQ58ykXy7Eh9gtMLhPPHPxDHiQqYHmKagXcHjzHJxX/6H
YjsoIFFaGgQrCqdSZ4Y1Xi8RXmM6g7xc9/Hb6VNHznseTj6m9o3pWutEIJrUqVzO
PoQa6i9mLn44WO+udRxxkPIsU8v+cwJY13S+rr5c1/aR3GmMvFLZS2IU+W4M4CiS
mA1coUZLxep4vsS13078vFbj+DuMlPjq2qkaLeW3osoZnYCNR75m6I2adGJx1uCg
SOUxY8HGgEU4K7+jodjW0ZgsWbcxR+fAoNuj4w8k5yG1LWXScaat6HTq83/0XkhM
TctuTSz370IQB/3zPaoWZyO0RcaJIfeTuDAlq6QKasN4VgXzRvlONCwfaZjrIrcc
FmOCqWszwPx6xA+/huQ+pYESmGVAsdi1YQx56n7h0/b3R5SRaqSnrPcnegdEnjN1
A7B7NXaGdnb1elRP2Wfs553uDXidR/gWDMNBa4UqrbkMOOPRtQyS6Xk1Es/p+0CM
DkqtlwzdvC0aZvE179s7BmBRUzvfvqrvrzqgvC4tjf3RVOmnQ9CIfsG5DkOlARlk
e9LB1BD4e/9GWpxjLiFDpMNw98OWHWtw7jTj4Z51w6LmtWhPFsD+14TGXIWzULvM
dH/OrQQWWOls+XwxZ59qDbhiWKGZ8BQXEbIcZ/IxU7mOQfiT8j/jRHAk6dR3udvx
RFdjq2ooQON/wQmwb1j7Hc+dgHtUbmhnVMksLAo+oQvAK0uhcgcvuOLAxMEke3sE
iVuefvYJXbRcQ59EK0zacliki9YF+ltMO41vu60Pp1e/XolCFrMfmW8IIAV6V2we
+vCXWbZqSyRbewsQiP5l0rMItXXNshlRIveepu4V1w/Asm/KeYODk0hFFx4/VutV
AI1myZXqPpvw986JjucvC8wCA4oFTWety4QuyXRbQTwKO3KaTwFSqUT9WdkeN0lY
IugFE5TCEQsUgvE9YK/MlI7wSLDQmgKbYVihnbj5dsjoZIIKfwxIRQOr6SbHhFbg
Aj/E2FkRjDlvYcs3Uy88JjQ/QoIB32s4gE2xwZk/S0p1FBcwC9Dufaw/vYdAcRjS
zXjfMYvyZ07wtfSCntmlj78qwj41B1h21i0HiElaRiuSBkhDi06XsjfhUUEaY6Sy
vB1R/2rZu7cYJN3ibEKpshHLReOd7zz2E8i0QgYvxhEmwhsf+7QObeeD0k9fKH0X
9iAatgEo/ACum9NQe+iYA6jNIeBbLQsBZ57g1cpx34k8/a3d6cUj+qeJq3LFLyOT
T9I1l2n8R2OM+MRsZ3LwRsYWn2M+bIu8MdkYplLAwgGavyBMuD2Mdn27I+qzVpuf
eE/DvnzinrHwKFoVF0aKFb9o0w1txQMCinLUpbtGXmovZh+S0eEOGWJfY26ibrm7
O5kQHS+oApTtArGOUPTzVtMo/xHunZynlR7P4+Lussz3koFnSwiWk2bW3cc5VE2D
4jmjxH+3PEvYKylwYRMCKmyqGCrQqJzKWY772SAwBi9SK2FDxajObqEheuw/EwXs
Uwdp3xXYOoI6gNLkcei6xtJrpjwqnOSF1cLrVTx/wKSgr9NRgv1ohxTHTQIfUULS
nCLlokQnW8IY4lkPTfuDYX5Pvsut3JR88fcfWCuIzbW+eqLaAENJKF7Mnx71eQDJ
RRveAZsoBIsWLGbfH2U2fn3b/d+6DN0TpF+MfpATKlCxHLdjrGbuR3Gb/CkkYBYK
En/ZVvY0I50DzSrOFbiBWHgsAEE0G2j7rN5erCnBq9t9wYgd88Q1HXzGlThEbfxj
Z3ZrgrGfpHkyRkHZ0aJBeHfS/EI6XsJAfORIQhoT3TOLR53jw77z8d5XzaSg74Yf
VjcZscWet7xeBx0U0MupHiMfhzlULXJQmQnJhBnnOIKGV85cf6yA85TIWjS2XYnQ
o05EicSxd3YqjtUeg/PRjPIAiRZhDXjBqyZvoJTAt7hcVCgcdUW08cNBAoNTU7KN
Bi/RERKkbdNYRPr1rZLHSs+7fcwNw6ZKmw7dIro8clzemsQLIlhVZNqYHRtWhEwF
LnZFPzb9UXg4Nt/lz2LsUnPXuSrL501tApRo2fLEyjCcQ8p2yktWXV/qA5TJGTe5
wJrZ1CcCdt1OT03zapD18FDj4K6ksSXdvUN4cZP+uvtIv2TNlHmD5m/KgxjANovy
KtetF15I+Skd6GEtAvPLG0KHy/tP7t4L90SvhoC2b+VlX2t7lvN0ChMEdCcXgvcL
2eYrKHbJU2yrwRTAy3/zF1rxjWc1MOSwnFr9m7HpAD2zkQkD7RwLkJ6cfN1CIHXk
uuA6YUXeWVEqqVdBluh5RpvQGO77lsNqTR9cdq0NYAG2ZZkVFVUQZ6w/XD/pkzZS
Z4dbIbOHZY5Z6WbdER1NKFSQMJN8HaGlTJDdRLoRMPbPubg+OlX/LWQvuWxWyT2A
IFKKj8OvnRj5kvAz3Ph0xQ1YPszUqWAh6Id3B7N3d0k8SFuvim1HjbEypXI4SFPK
IcdYsg3+7izcF5XXhjbvndegEkfWaIVJk7rMMhhnlANg3EoQiem9QBDGHDpSSnmO
tJ28G2sG35MY0uJl0uY4cTH0ktIpoFTe6STga59ih9klp7vLAgflxC2icdbaTFmD
6bGiPekTSIMWH2njtLv9WXD3XmNxn+vZdiO5KdW2B7S1PW2h0NDrCaXI0TIubYhw
/DecIha5zD6nBj1vj7aAH4f+wBgJ9zM81QGVTzFl79XPBXww4dGRaBAvs7B2Cuka
RPVqnnyww+E9pFPkVULYuArwso4wj0d3ecPSZWMI3yIfsMYxTzTptgmnr6K7Tsku
urUcp/rEc7OS2Gy0KEZEARB/56AcThl5/r1D7KV8vwNkkijxYNtDG04fbenNpIn6
5cJrLREavBXYBRRsZ0X0Ru/ZT+NoQrvdf+Lc33rq5WGZ2J2QxTJMurBHl2C9yt8Q
Fuv/y/Kqi9RKTrlbH4GY+R5cKpmampe+T1b8DieDrb/HjXyQtBowf98n0su8JVro
3GrGO4E0zuD1licFQDK0PQH7pJEOOoraxzNz76EWKucLoWmdHWomAuFqQBWEchTa
G8o1apvNnNGK03xj+edaR+iqCG0v113Ste/RgJ9mhqGCvyUEFxsK+irqQ+Jq2T0l
YwiiT4T8HAN0UAT+xn71sueKE4/MukMg7sYh+3tCNIhlj2wd4rWlwOq9CdRWppw9
Av7dJIBaU5PBtiwB/eZSvAWYXzk8vziXJKG5+0WdwmeMRRRtdKiVHx8UKZ/8/T1p
ycFgj61IJaCj11IMzX4W0KVGjcrv3PAFgFgSFExJzCnzTT1QVLsgCsjHcV4txtor
fsFWeW00Vku07O73TENJxP4nWK8Y02ZImEx4rY8ihr59OY26HuNr3bgjBNfGPGEm
MGVLhcU7nsbe3t1e+SlV0+BeMBp5gZxGCWuc2zdJtF/qjPg338wY5edJl26Soagp
8jScpdadaqiatYhCzALnoA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dwyBm1SjTAx9j/sxZsG13p4V6dmmMarpti+4vqkeNgk5nW/oOt3oHVCgGbw1gI5i
kZnEMwGH4RtNypmFtD8XXe7EqzIz6EjAZGiJGQ8K+PzLFxVQkly4MZPvWS/2q4Vb
eBb3Dw9t3qnMTAWyGHHqwIGbUfv7gPPje/5oinm89aOmDQaoUn39ukJ1Om8SPVGL
Wkx2y6fRfremVTAHfzDu/kb6kRBaF7HW2In81Bhp/Mb7H1q451bSSfclxOdkdSwx
jeLe9G6+9GxP0csMqgVguzO/kf8UoW67cVNBhFdHfGl8UuxTVeMuhLMZFBKAouDH
x0y8GVahgnFeQGBbLhDO0g4hvD7QfR+jbxdp67WGS01lKmgnFNnqnp0z6oRlxen8
2Uyyunpbp0ZFgpUtLvwZH5ohotqGCK+x12JnW6R2a3EOqQmtbVBVUtGWNH+Erhf1
78YuxqG1q9k3GwE7ah6x+gLg9TlWfV//1cdHI3XBQKNOT3P7uiEnIT1JVW3gftH+
9ckKiZJ8nRbhhpSRbcaVcRJOkk0rqs/Thd9NxAgRvLh0X4xn8arkEs6A+LD0vH3U
ePs6PeOzsEKmx1RMQBJk6KD+WvFJWAeyqxT+F62uc0sZa5l+gTLk0zeU290AA0FC
Z3VjUr6UOg6kM8NcKoCeSstw2l9nPHwHefnoum0S1JMkz0clDeWrx2G16OZ93HzB
Pmb9SEGxjix9Qcwk8P2ThjTlc3JVApCFRnFugI3z2nQ1L2AvEqustItKeyTZlhbv
z8TrDEjX/dAunEGO2i/A3YjqBVHpBhxq2LBTZBVT9fwCea/Dm03hQzCWArK2ogGB
V+Sj0eoyiF5KA+w8Ier/QK7vmHRBPrriR5R+sHIRAzs=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKdT9vJgFRXdZIV7S6aW4c1npD50I58efiFDuiOWGzqmzn9mSbcWwaHpp2Ak4bUC
nAfkuIkYGKMOBT5Nudpfcs6JkFnKlB0VYzx2OHJOyseIwO1Bv+tjVep4CiCRDvWw
HuVBwO/iXRJlhpz/8Y0Tl9zhHQ1LIb37Ref5XR6ATCxU1/2mhddnAYjFGOAEMOv7
0dvlKs39iXx94MFOaeEXGUn00IP/ApsNhuLyyQoawfc6h+TDm1c7Yo8y+wgaUIUU
9JkE7sYw3bH2B9J9yq3FGLvVnZT+ELteW9pkwx5Au0p07CtrqQrGOpHa5a8013es
S6JZXa2oIPBmjf9gi6SJDiGg0roFjFG/BdlNOmWeNiBzR0hSoid3RTCrb8O/qIWo
uUpgjFg53XY0u5m0yvXBEKV9mjlRlJuEKivPwo66eDg9nLlfVuw1N73bJSvo7MXe
AQahmI5TnTmpooSkmDHyffr542H2mJh5DHYjdw4lgX9XbuTZQ1zJGQAHm6zoZUnS
mf1eiyKCTz5hHNIIvNPh7Vlrdz4bqeZrvmxHJEu2iwekPponvZDDGus1kCPredNw
8jNJ4m0xtZAjFmuaHJmQTwsHxdhrAvrL5Zy3O6HagqXlsqO/wfxEg9GnKBbCgZ8G
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKR17hDObQdKF8NyNRLH19HxD5cf2+VG6c9x0PVfJRf/CtqfBS1wVuF1BeeIwdne
6wZomYmFE3Mzv6Q3xAdeGNMnlY6TitG0rssCQMpSqlDoaniunSlifKiraYD728eq
QCsSQCnPJ6tATc1A3w2AZrkkbMEcmM5L/ZLbtxjUZfFzqKDe+ukS+eq3kNre1U9J
kfD2RmV+3ctz1wlWofDmK/WV/kss6yiL/oRH07O6IH67D9q/Zv3GtCn9jkwx9BDE
dOhTy/lBXTpI9VcT1rfxpKen20S2FLAHZuxMjEwidPsQisaci51HcSgo4Kay+PVy
R8uOIHvurD8fiPVAlsyWbm4S8TkcvTAesXhw3z2FWJb8j/+dXhO4/YcPGm9i+7SG
vwz7T67gScqR8mWdR7rSTLAa8D+MvihsubcnX7X/cNIM7WIKGR/IgtKuFykm2u+z
h0JcZAiyFVfnFbhr0JzFuhEQ91AUFUuVK9DIzfiWw+5Oj27qxoHSLLowpUo9YLGS
o7ksEc93wT/I5a+40JpbDR0DjDPCmPXrgKvs+DyCsYKn+jKzW6ti7bEUrCQRst6T
hnTIkJd0B5DMsNMox3SMHKMebLEqPkVorh8vmBIP7H+3LsVUPnXsq4LOe43drMuK
5lOK/wvQhBqeLPRryq2mLRCKQn0Cg4pi/0eofKauLmz03Tm0dFX3049ZT8ymp8tE
BsHjFdpLoOGwxKLUaXfyjiVxxhlHhZPtSqYTZmQOViKRzTt1V005pEhEk0v99DnW
mu4d2LJiGTg2nQyamQgBYBEcA1b+2SeDx2OQNqgofI64wr03dUELMCGGKtmBGsV6
S1DO9ozZSwQpdCUrs0e+mggzRneIaLe883AydG+6AA0XLUx1aEDbfZojkBwOO5FN
x4p/ObAZWNyevHwzrwSve9CQQEa1Yp4GCmedXCffjrXXUBCEiH7QOCSana5OAD3I
47TvmoBafvVvLA6GI9fJUL/zGt3z4GGpO31DEFtOFGhiVrz4wxU6DcFiQAkkFl6s
GSGnKWapjWahYYuoTeNVJm6LFxe8gy7rAYcvMoa2COvOwwI1m6/P2SbC2u3touij
jM/P1Tx0CeH2IQWhlgojUazgYupjVo2aozs5jq1kfKsMbs8/JE33Jl0Mi9bnJP8m
PZ8TsQBzdVJrMm2OwJ5MmxovnU2/Vi+sAouBsHQ3MtO1mSv5nHWwD0ayrWytFCuW
NtvLFw919ayigVtUCMjh5frqdauokLRxd1/YEYtv09pRu7hYVZwoveForUJ3A0JE
XwDlRHfe0bj4iAvlT+ESOoUXdxGqDgSr5UrCRPf5H4Vtl/KpMAlwvfF1VVcMN0Am
FtR/CeOykxmKpN9WOQGXS3tFGLrcgWUycP21FjrY2Gi06LUrHRPUxzjsh6RA6YU1
HBN4IKvtxPKkxfn/7CnYKbLVKA27NaArWRFFP6XsPx5Ye08EWECfoOMfz0lVkh30
WbKP5Nxd37uTQooFwGM9pjz0VQ9qo7uFpmTj8QtWDX0MZWobfX67tZuD+y3tcmWw
IjCqi6IZwhbCeWn4YIbNLWOLvozyMwRoIDjXKfTpDDCl8ImnwtuQb2u8S6Ip5Sh5
PNdB3kXX2+igpF0di6CHiLme+2TpE4iN6TOLDADSWdnz1ZE5I+Xy33yfR/wFn/gj
ypFiAfq+3WCs0YW0cUQz7yr5II+HN9Th4MCL07l0MnU+VpPKTxQa7iK8qJfnJPi9
OOEQ1g60jI+m1/+6hAgVQd2/G0hrfTWKosgwEmwnaY9GEoklxq/taAdPq/e/tjIP
0r34efXyRFyCE2+Ns9lzgJyE4PpS77C/J++xfMNcPUkhnf5ThF6UAkL86oqHH5bh
UL+/X6rJx3X84Z31QMt7YyAr7KJOTXV6hjojIxlaAu3cwWq3A3zbmYbDSU+R2zIo
bDV9YZp8OhUyDbUMlGkZ5Q==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAvDikmGlGbP0jO4lTQeJMAcObqPUr3V+xU9ar+HdOQdXnFuk1CktoyVKsqxlbbU
lVep9Rc85B8YhnRafgAXO4F6qVAKJihQHSk4N+odbG+Z47AZA239K+BRNcP/VdxN
6rNogzdSl35DDCSk/ZVHVEuPpeW+Ih2uQHSNTdR9Xb66b4hFQZgk0f/pZ63xrKxM
N671AF3NaXR43ZWiPjjbD0tXHAnUumUy+QMsmDYbK3XqapAjN4TOozgSlK2TWjzN
Uf04tx/82gCSDwWNBidDmf8zmzSHsbPQxvMHdD2+zaRJhcjRTxmIUdcojh73mB98
2Ztxuc1IT0StBHaWP6/4oZ4/0Og2Zp1GbKSdf794h5H4q0R3aEd1qnz5TVVGjGFS
n329cZa0PKDigL+eUocfDJu+zcsnmG1ZaRAzrK8b6yjtnKFBMiDtkhrbuS3xTih7
+Wo9CWDAwFjlSGRpOU1sYr8M2nf2qNMHm7bwNUhSqKpnPl/3l8lWclxr+znl6X2s
oomZvSBFBa5b6oxJ0Yh+pF1/evSJNsiOGKmAJv95ohotC8J6Fn+bbPklYqvSJ+NU
9ddfdwkMGHLe4PmzTgGfKk6QyGAXX7o/BORfYKlgd9gOT6xoXYcliziUOFHaWgd7
t9eUHkhzqs2C1fw6mYy1eKiZUx23hlNoRuVs5ZeKszbWMOeVT+up6Si8fOqChkGw
hk088M1zo/JBGDWrxqf7qc4dI+ZTZjIqSHNaR8XqCHTsNd+/1mn4RG0DFAKrqmor
QA9LE0d8OODcDdeu9gsTU0+oCg4MweoVU6LFMjOph6inemfz1GIsf6BRMPRcBqQA
fFcfR+wXJmXR6jJFJF1BTNCXh0h58waEz60rR+0x/op37dEhIi5mOrMFgVQiMl5I
EIWpxBmhRqAJ4rEKVEj1wcqS1tdSDaVucMt2ouqGB45Vf+emnJnG8St9TKP9VsYg
fF6KkX8zkL2m7C1lX37NfvZ6EJ3MKRDwbqUNKKPDUuzEAwRn4jVFsf/T0tzmXoZU
1qQBpD9x+wQcMCqUTq4Ow9iL1n4V2wcm86dNHjs54kZJt8sxq3s4fyEvC5TeME8U
Cpp4HxE1yhfdHl5oRWS396nTiUD3uvekqvyQheBCdCDnEgDNnSAJ++JukOtilO6X
30D4uef3KFvp21ExNE+M69RWI+F6gngzowhkeyMMd8UCuvhQFSRfrTxMRbF/xAxL
dn2XorGa2nTi3q4kVApBN2OKOXcmHyunORjs1Cb84tUgkeLY+0NcwIfCWXxgrc7V
CpYYtu9degeUXwZjU9eLGHI0j6PkQaBwSvzDl451z+L/3SuhwqbAMVL91/rd8nMb
BzsTE+t2xv0DO3AuE1pAcisa+LeTnICcNxhgJ5BXTtLlDn6mmP1QXmxR5JpwXaVu
SI+VZrsJ9P6Jx3LOVQZeV1gbD+O3vBnrm7yaZ/T0L/bzKOaGzobUcfoGpAv6szgK
vxIdFoz0INbTA2CWeSOrlzDIheGPOSH0PgLdnLW9Pc6mohPMp7TuL95enyIkImLM
TuPQo/m0IGGnbSYwOV5uGPWwCczc8QTdGtjfNouxENSVZZFKyCfMqRIGYaGiBm5W
PCG/e8NNyZY2/PkosvjgkQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
472S1XKFSSTdkhhZTrrHyl9qOishOdRsNCaKy1N1SqUaxOC/cBE7HGZtlG5DcWXj
8pW4/OzoTsNM6cJuXllUzlobcNqHBFnEP5bzsFJ4Tff/RY5q0+2e4WhU/LPcT1Lk
Wa24JR9uV4JVTvMvhUszM//1O6oNhSKiy9mMaqeS1G1PTrWYBcX//5lkwSGLnd5j
ylGtIUdPagm2vQfO+4vvvqWIJ+3gFBDh57gl6bvDUimdmBnPIU1+mqgkGsf4pIlU
KcGCwZ3rxnSKsvi06kJpcm7MFBx4t2DD1bAs45OzqP2zKt1QuvRSBhv1N7lSj9gB
ItBLYyKOZV0o88aFpQfe9mx76rbryw9oBbgJCZO+gmiE1MU5nL0ptFcamkWYAk9n
a6LGtdDSR7bnH+6ef3M1R3CcNXIn7Az8NyxjATG7s43hK8B3+y055NV6XrcppKBq
3ZeDuDBwv0X0+Xa+FEal6dj/mwQfz/h3OIMfpv7UgjYPZ+X6TRDwJjYRs1uoUtVC
6jDBIV1LfgxdvFjX88XbHwPgmfkyu5pnGf6SE9g7tpzQP6fDAMg4iKQBZBaPz4v/
qOsReE7GG1qXO/hihmLuGfJ+5yvUSzxcLuRmQkw8Au8WDTGB70hWMScKyc0NFFb/
DEPxVKN3Saj50lNW1HTYeYjKnBfj5VhgnV/2Lc0jfeig5U4HiFI4y/mjm6VrbEdJ
angkQMPRoAm34uYwtqUSwW/my7ampEkGtcoXlcn3Yn211CzfluuV4qqKhaaril9G
59rvoiB/phHP3+VZn2MV8VVHWga6cL9ObAbUyGbWdmzhsp1PuXokt9tWp4Fnrymj
KsyruOvWvXYdohl/V5kTRh4VNh1/vDTzbTiQok5rUGepIlmJ//zrPsxjxRnlMb2t
5LeeCIRpaXGJY8LOVVeHGSQAqDTYOR2SlUI8sWBPlrzNGRDz/l1yl4DX6/niNKPf
3eiuxZc0mdj2U7EB+bGJqj3ufPqEM+go+d6uXvs8Ge5ANXMCrPym5elsQCHMJ59H
IB33NZXiaQAcgW2edDvH/KvLHSYYUeZv49KwXbhqJRuhLZthWzhSXIXVUBc0/hA+
hGVmv2v+s8u6kzjnj+20Kg==
`protect END_PROTECTED

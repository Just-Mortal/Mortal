`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/NGyidR4cdEqpdIvhSq8zNPqAzpuOCXJE6uoNPBlHgVKqLhEjzbcQwXNGLUCtsi0
J4XNAZFnMvZowiuA2GuRtOOg4ham1a7rfj1jBjxDvYaeVSMuCqbR89s7YTGu7suo
77F4OBGW5nVmsXJj/IFkDf3KsDJFZTReW+OyyL3t7NwN4yegOglW05vCnQKi8PCM
m4B0cHZMWOe4MyYXlkI2K4vE/QY1jk4MRkBdq9JahfutA6duADYOz44EUqu2puT9
QHPJ4MbjpZgWCLndrmnU1AQylXDiyXyJNQ7rzLM+jh9ZPoiC+SWnEI0PwCeOGpg5
I7l12elzj7i675nVunXTKbgvpN2kq9XKA7cG0S0HtpBOpSDsYgmJkpvfeWUvjH+f
PS2xdHtP7inTbf6O89g5raWoSFQ+yDK/xy2n1KZkqgmhDdbE4HJChvH30VkXrAXY
IxkxzkClDuxN92YOTDP6sTSbwsBliMDR1b/qDgpvzLj29GXa92+JDxwY6w+5d6E3
+Xz45Z5lu4XmqJxMe6YkTkuETWx4mWlJCLSfat/D/KDHpt0suTa2yZz5MVgGdPeb
yW7lSG8fEN7jvWdySEbSQHLr8Rvfly/00KwY8MWNQfwh82/V9epgGbytzVr3CbPy
MK75Smz04n4Q9lzV0So8kCk95jbDDPcEmj0nDqPo7eWmzUWqgKhVX2EQN8vzW9PF
lqLhqMiF6HYYOsffzUB4xUS4+5cnqBeHkxChgdgKy52NPao1ZNHgpqR+32jYNcVE
jYMMTQqfNWFfu0ygYpTAb4KKDaB3+AWiFTMDnqeBKyortRvwF/aspGP7JRlP4Sh3
jthzA14kN7YkAtiz0JUzSMgYC6zYlS4EskpOeRdxL2ZxnaBkhTcLBdQGzKXSiHCc
`protect END_PROTECTED

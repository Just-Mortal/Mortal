`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xCLaTcJHS2D1FQ4M8y0s7/aUxkKfJzh1b7b33ScH6/agCqT9sq6ki8wm9S5xmYCO
7/D52S9fd3sMJPNC7Q4YJNuPlBoJtahE2gccOC8dfkjK82xZaEe7nuFTIM0dA2oe
tcKybAu2jXQdyBt4A/alO7HcJvNazGeMYlRtwOqik8J4wnglOPaw+XdzRVgoSny7
LCh7eyfvi6oULlsmzAfQmGMt41LSZKj2YrI7Qk2wgc2VE9JrsrWrQ37+1rHW2HCJ
FSnm1qeVuKJq+pf+Q5GSwTEd9A/xSF5N6gvKCItlKwPhXujszZG6C4ZuLjQWc8Xz
B/HjowaH+995MmQoZkCtX3zkMJkGPs5+9AVwrkHKE8y4x7c/UgqhKnKstQOuj+ZD
2fOJF9Un+G4PPIAAF4KKmOm3kJ92ocWrWePLZs5jZ7Aocss4+b9bWVJ4KEkmi/7U
j0/Ldo0z3hDs3vH/FQ20okFSaY05niekErPtNTA4ng0ruE1aWs0E2J8/r4DK82FD
KZm+auna0U7bV1todiuZeH4ROj070XmrVMiJ1h7RbGz43j/AENUIYB82MN0PeO71
d1/etFxINGBozwK0HdbtSuyED2JuBSwimoe1oCJuZwyMAuNy6oGcKZtWWd7ryW03
OoQaDYZNdZEqpQDnXoHIIQTBxQRQYW4YIHhOpPl17uTzMcmTL+nv2ZChj5ptwXZ0
NlNOczAlVW6fyJydRx720obJC71PeLd20TEv0okwLMho2Q1c74PQ/7V3dV7NT3X+
K83q2BBWuadexG4aCWTkPwkMZXc3YTuTQOS2W6WLVAJABMUaoj6VUe5GCMabzljG
zNzxZWlft5xlazCk5CND9eg616e2xM+SpEi0aRwUuePHCll7h3VUzRMcXGXPV5cJ
m2U8BFHlorVtwNA3ko3/ctcHDVnE7XCFvsU8YjSHH5PfnT82Q3k2gM39Ht5/RWvV
R/YZxmgNfVUybFnoBNpIrG4Oz0p8xFrhuzXpOgrundGJEqjN8ifC22mtvn6yQopd
CxAFmtfuy10VCWqmEBSWdpv3zUZCClxpG6OJqD6++XtE3MFQhBDDA4QwBWqjwxNR
Bdgv5CoXrAzsD2o9oItBXTGT/lexCgRRWF4wb/qIwKTZGAuBGnY9fz86DAauFN5M
ahQ9rC2ifMqhY6tGfrePUQTKSRm+65Kvnj3VG70uUxz+oDkSzrAUd8VK9oFxTopC
DiGjVegmpOmwzn8JvL12EGnGapeQm79cDLshI0Vgb6Q3d/ihsTlcOclgr/sfgoEV
erK+OPvlZAdRN+kt4JEaaHjtGF4HFkPwK/gf3YwSYBXVmvbLI7wKtoyOXqcng1l1
05KUmYlln8/tCWiptmRWv4W/6+QjZTS99o8Ahs2swAtwZZF2p4SqiIOwzxhDzlyM
lPQmQSJyVektKr4aDzi8njAcwR+uwQnPhaXEH4HoeTK50inH2TVv9T5jrRvHnx2Z
nDNaxEQmHkDiT40QKF8jZnx3iWmc6Ot4vJ58SMOGNjEecxRNuByFnd3YmBrWe4Ja
7n+1+Qi1Xh4tlqYPy2IsO8GskQgjbf4rzBTzxEY3mN1J8FcwrJ0sWpqjWex/8A3D
piSzEPe4i3IeqIb0FmJrPICOBsDbUZd6cxiAIetAKdhIgw7Ozdcy2tawGEZghmbw
Wu802J0/9nlvaqr14zC3prmj0Qrtw4ledtE99zVV1OVKK3A9fl0UXztJB1L3txTi
Gj4fQngefBxl4raFfZaqjzGX2XKrSXZ777SszOtgva5OaUhMVGGMlPkZo5pKRB4X
poCcfNnG83qAv/CQeHWkfAA+AVwbfcjEPCFU8uuZ8YRwgT9UeuRL3uhazzY8KTId
BmuMaKPl1flLqmWeW71+rq/uZMsUwQMfKpFGHmOaJOZawk36lGcyP5nIoP+LY/HX
dNqUAYMQwbDRX2ekTIH15xRi55UfzMZmTF3jlYp+QoY7HPQ5clXyqRcNS/yeY3Cl
I0V2FaboP1jX13zjFZ3eEoa8K/UT58I15EIxey8iuubYC7GtJKQI9iyPqXyzaLUP
XDxT/hl9PuXJnfbE5kthrDNGV1G2W32et0fJYlPO+cCdZmOZiHB6SOUGRK4MwyX/
tgQeUI2oJ7IK5Bfb3Xz1Tgu8GE0JvbamWZ2n4ApaJevF8i4jqiI1qCSZ5EkOP6U0
QHd24FRIHyTEp5oB41w+nrvgpCcHDRMJmKB700gMfCIyYEOceYeXUKjN3X2quXFW
Dh21IwbUBmry3PrpBhG9Ww8VxGG/CgoWy2Bg77R13ry+Cipdl6GFzDPCpS9rhAst
3Q9NWTD3zKhztQqZ6YtCN5EQkn6Jjjby3s9jVcpAaKBjetl1PdwGtwz9LNZCFNV3
RN6Ldk97aeFJrfxMxoSTL+YWCiRt//Qmx14FBqtWOgj96SyFlSZa+dW5QLKfkVE/
5XVDlIZwdIvedTbbX//FhPjubVSXwWmVetgfjCyYsT7cw1jivZ9ETBm+8uJwPTq5
/Y1VOUAoPXWgZRCRc0v8s8ix2drtKAZrm1gyE/z3q5EL9XF27Ana0PlI36EM6KGM
FrBcHspr01cRLN2giMwKynqweN5RTZ9MqPWM2mwbRddWJtsoEIPk4VEL0QjiAF7N
oRT03hHDdrrhadvduXDhdK50IgoBWEEODvzJAaxuC2c2s6napphOiFm0BVNiu0L9
CNxwEN8AAr/vFCyXfbLMFYoYOymP0O5UWEIC3sG8foLAo5u2ynieqZKbOGPoxO+S
f7GLfJ+sP/Rk4w7Sy5UQrEJy/+iDA2qSELnMuVf1JG6pRensnvw2mqVMC1w3uNyn
uHff76BPaRwyevrI7UneNDFM8GqY4JFIQkSeKWC9ElZaxOQJySDF/w7UO+JF1Dgd
uJgzrOW7OpxZEPfkoQEmum4mpmdB02wOAb+3UUARtZmK1G+epU/0Z94PKSThRwq7
dEo7U9Sa6S9IIfxbUZvf4PFD+i/+MO8KrpPu6AJT53ttvmNWUL6BF324zIaOVOeQ
yfL0om6Wc/E0WKFx/Ml9FnYtJn8mf9uy0jcqQM8gH6MT6x3AlUQ6LOUYz3ugEpun
5kczQDI79lvegLvBXnVoHucIXHK1Jv/kV7LotxJNDF+lI/cq1EghTvlJwnQS5gd+
TNOVgJp999XRxYsOgDXAX70Gj0pP4sT3SxTKN50efQit7yjRaPT3WC59JT9UFIZL
KGQ1bd3o3sQlTGeViDSXmJNRSXLzSTmwtlTCiyNKCRwhWZevGpE6a3NAkIn2t57e
Yt4iWhDIb2EU6nNDDDQS0aJNJTk93kMt4kZdeJqGcGxxbYFgcZGsiqHUpjcTxonA
kmZt4MvjE8oC8siGm0uackPTX0aUzplJfqQui9maaayrJic+LlyzYinJOtWf4VQp
iUQuOX6PvGxG/tZwyiUr05b+rJBBBKygfW+QUYLhxRraap7S2AkJOHJjhiVTbFaa
Xl4puFp5559GnxTrflVxmrvLOyqpBdiwjUsAcGzcO8s=
`protect END_PROTECTED

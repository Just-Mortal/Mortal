`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xv7E4GGB27aAyd/F0s7YakUetwsSWnGojKM6/3GdMDwSnkyAeRVykaPeWOVR9lCW
XfZ0oxAhRPjXJBkSmYYTV0zQDxvD29kvEI7pX8bWnywroNoOrEFviohS5Gfn+yRB
Y1/rwEZAMAl0hVw0hYUcWpkd5mlCOj4fHrVtRo6uDXLDoscxrnXgz9D3oRzOmFVt
P3aqsr9Pw08jWIb8qDoi1yUQjS3Oa435pd6INBfOAMPTvxRM4wkoT4Eb9+AO2rW5
7+DGwidvRtjL3QuBYRDzRimoDC3xx0eXSDrahvae7qzoWYHUVEw4Bd5B+WxSzhfR
Ibjr01jWoZ5GP2rh8MIJva4JfDSRoBcO/8yaVXya5DNFw+0quiDDd7zb5WJJEwc9
`protect END_PROTECTED

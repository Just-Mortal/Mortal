`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypnPpyDopbmNx0y5ZbpmWgMoiDq8gpI+joUIJrLV4AuI2aqISH8Uf9MjdvxkJYFx
3n4m5fWv48BkRHl6MBk0hoNKTlF8vzSEzh+ieqakLyNEi/QpoG4E+yX/GgvE9kDs
g2/XATGIE0JDRAUufwT1LE2C3zW8imGMv1wRuNKnj1039bV6eno4YjF2/m+/Zfjw
LO+Erwx0d4Iol4mGoYSloP9dPdsNO5y7ftIjfDWqdWKnH0+WNA9sutjyON9AM9mL
ybl1XwURJ2rOXiPowQHex9FFNk2xYG6j4CB3Ut5yWffe+jvUvIzM9AjAiOjuJz2t
t4JLdFDpJZM1O1BRjgBWze/t9F3CibJwrvU+s4DgdX+ll1XdBINIB6jFwRA8J5c5
MTrVb/0OdXYqHDeSrU072r2tgZ9fz5UZ4LQyHV4Apb9pPFV4BRCIlBEpsT3QHUG+
TZn1uxoUA4Mj80LIx3cH2/yRS63hTqsZHcuvCkjUDvltqoNVy72j7PGsRQKpbhcD
o2gVCgj5wiRq446pXoxB9YAbXAGcrNt+urTE0i/rlpw=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YHTmYWfrynsAcdves8yifoz1Ne7/zHwk1A1ob+TDs3C05PNqeH1dZfdCLPuB10XL
zQs3ongan9JA5/6lwtwHNZGK4CvuQQ+jKaL0X6P9waPEsM1act5YnIndwsgHnU43
sSSWU4J2aJe/nuLX9KbUyBgaxcRCNdFzi4Q8fLUa/F+WzEq+eXBDFoy1g6UrAw/5
8NuOUqLjGSuJceneA1uGGe6l4JwPFdJYC79D9g1MfIoVwSG1weyI4WNtUS8RiPgo
K3Yra/7ldUFpYgSbj6Cqt3lMwal6Nwx0PI/cB8EaR9p7Yp+5Kr1qg7EOb8Bi0SVh
O7PSYDGHAL3TuVdWpF9kwIpPrgfG+o+N4Hf2fZ1S4rinLi7EVpuNrwgkUT1r/jUz
meh8xR0vGqwaKhDuaHMK9pH+hd2U1vVjKqBqbz8oPl30N/K7qxc7vptEEIs3wexW
5kUjtfWO+wFHkE3R35A3n7n//7BlxmQczkBQKW6XbbDdWQUjuwLR9gVIlBD/2YVs
srcS4NylWFQlIKH0ByVKCnD8SM8PlVSOsOT+Lbkh9GtUQwUx8T8XLW5jsL3J1IwA
VyKUwELfCo/XvOrBiwKzQcod1oKG5yITuFD+VowU8bWnAYUL8828g7Ky1xhWKp0w
H6+4yInA0b8A4rmjPtac0XXQb+SyHUv6MPuQ5EDtwttgIdwmkPnxhZxGvx0wbIbj
7mHOBxW2IhX5AKQglqClNFKoKO+M5sgE4FBpYvIGSKZlbudSbKy2lsPJNPfWimP7
WQ+n5vmQtTUn5mL77sQFS+nBQC++G2xrxIOsR6QVRA9YFgHu3OI2u0GOAUxG/Y6y
3/YludtS0gTJw23kmbgiNcNP8xGuN/HCb0D2hRKftJRYJ0j0rixWYSRiCdnjmgDu
R9w0DNAa4TVFOCEmJJmKx7AsXKtYGQTLqE4Jc9I/+F+DLbojLZYsdVISzStsXp/A
ZCXHrS+nFgbPCocmPF0hiysC4t7PsYta8a7cfJtYk5BWINKc+IrsFGla3uStos2a
CazWJuPznFvyn4vHkdVYwdX1es2QxLUV4xj9ekBn71V7ZGa5VMD8/9a/LWTQQg47
xVMvAPl8nNl7AkW+ejBPk3R8ilhGmV8oTsgz5s9Ee+TSGk3nrmQZXrU8VmwH9tuk
mmjG//YqKTmCBCx0NR5eIt3mrEZc0qtwIhDNqRdwm0ThDgz4179HoKtsGthTPLpw
Hrsq08Vma7HSFmJcUYoL7daXXg14iKXmM7HMOuBoVdkkUBEl+ilzw4LbPmOpzVC6
cMs6xGLDAIev4SyPZW4/d8IjgtTYqkCi8KfpBu+NK5ex8UNlWmWIYptvzvfiAq9C
P8Yw8E+m8iKgaUNrAhXhA+Ii1GRSRJNDCJp44+CYc4D44NrZGWznDuvH4AHZFgP7
JChLH7qym4y5tmI6GtCUl3pX9z3kLprpiVQypArrteTq+wOIIWEk49YKhSc5Dfzr
HNK7f8FC0f94jUwsTraqfoijJUwmHyCpBLKWeUDDS2GxcG1bsXyosuoG+GaCHZJI
DgRb32rLV6dImQyfrVu+EGhLxV5j9jgmlbSB1I1gnNEICDQnLCQEiT2cD6ntN9Ak
spC0T0H5qZgKIAD7/wM7OtxJwRTdbGOE2gBSS+98ql1eANrACgipqFqyEwkl1uWW
ijtWyCfZp/yMOYW13aCVCRqBurp2N9vFI6r/4bk4fteeh69XPYLuFPdNnUfjhwlv
G7mYnWoq9BGMl03MpVGMWA72x/Eb8/qW8ticNOLD35PMZoSLpOhwTGFj0vdPaCrt
oeI8BgYXZJ5/XwB1DiIbVTAH2gbLJYzzvbTt8JELV7Xv2ITomeytW1Cv2+OIg3eh
HlKQhwUKtHyds/4gCBuXjoJpfUFR4Ph57Y2R3yy9UsKmwv3wIbiQ0tooWovLFY6X
fRfINHEKdUjT2C6A3I65Ckbph1h4CPDsItT1+fIaFT2JRTRRg8TeiWCt9k+gJAWp
nkoA9c3jnqdHA7S1r+brTYZfR7PGBe9wltEo4FYHzy4TPFygvTuDAYPGfhVFNdzw
IMviLmB1s1Y+vFB2PyVDkxxwKeLt//e8VCLNAdoVE/lin8h9k74VL65mjc3RR0sj
RsqJijNr7ZoaxeJHjHau8uyx2jd/p0GWugJdukBnrM84KX2oXDRVEqEGE2ED+us1
FCZD1G21ahR+9bCzVGYaQkUyWAcIfApk/ekri0+JGAjzdA8VkeIb12bSPvkY+4NU
/+xzEju0AK/msZ0iwubwr3zpBt+VqzSmrKpTLT6aSSS8k56MnKJXG9YKtMZF6vUS
Yy8SR9M/3e+dy5TsQPlAkoLqVRJUTsdoFxIrelKthC65bpXb2PJfbiUQzaEj3Vba
nh0s3CGF0As98EAO31DdJV84l9Z9f9ecocwscXVSSjYfw0C8oDfD8tO2Kbc4evbe
qKnE641I/wmSD0XjPI4smP9nQIXKtzz0CLpiMg2xYNOkopdGe32WkG0oO9VJCqxh
5WEhEOkLxEdYYiIbAZPd+jDM+pMydA13AOzXOAlN3o0aCYqITqee0T5rYFaQ4EEB
4UfnmVfq3TKYr8j5+p4iKTrqVXEci/wxwjqUEYWo0bGDehcvjMgS4WfnkUH5WO1C
LYkltakjVUw7jlp+ELr3RVDZ69XAf/4O2X90vJfCDnxnKQbQVzUVAS+q5B0F+9YD
x+2myEfqVnCPgK2JdFT3MoHlFp0A+SUqkWEV+F/Jcp8Tm+yHLIbsmmYXCxPaD9tY
tEJsfjAV5uZ9y0BWIv+db5oRsq02/EGKsYCsbPfM0MHZSAhDGXqmxwQ9hcxkRRxn
wP8VmJy9dJYhTj7iO6OI68yZ5KuUYOBS/saV/dlEFEHKEcVVJiwZFFZoAPEyVYYi
jsRpIMiBgNE3nzsq/ufSsoWl6hY7LhOTE95CVGtcwM4jLjuyaa9H07RV+0JfynAs
mjN2hNOwbSmm1vUoJhF0eAwSySgwCtOni1nxMGO6Uf8hmwOYlX/ccj/NzidtactR
hes/ikFVmqSBryGFluCfhm+ToTGGReRNUtLvYNbGNGd6kinY12Ky1yzB4QZRM5af
H1GYdkMgYvfRH9cf9LpmbAyPbbiHsHn91zHxjXKkpAQnB0WWQ6RHXt7mXKrM2Mkj
j6x9ZYf7h2cgRRedgraqfCBbl+NgpGOl2CnK8C3bRczFV+xlY2CaJNkEj//cUZ0Z
/YViUhlUrKhK0ieusYEjv9o2sXQ/NwIgC4+Qgy71h93oCIxLm6han+d/ck4m0ilH
SWjCGdi2SyAaturGogulCxIzWzA1TFCoVpj2zLl3P9DF8wOnnuA9K+ohnWdDaP+N
x5DOheBmx6BGtQD+MeJyJ8a4UZXMYSkULzLn1qnVmqGG2TSK/2v38YAwX/bB0D7M
R7J/6PVR8Ver2MvDlZz/JGb/7AUGZEQbOAiMWbBzXYaJVL30XIY7jlk5HmnFgpIy
llouBPDEWd7rgnJuvwohdOwLbts3L3NHQC486jtMy9YOtnQe2BGxFBzyEy9iH2ZG
OO/u+zUfmaJaWsjN1APf4vCVi2JiZDkotl7sF/XahI+pKKKeCH/DTSoOxLYZAk9T
+z8U5khem0GwWQrJXc2c8+/DMvJ6XxiQTMhdcqMTB3uGt2iWGHMhCcXTZzAZ6QOd
aKTlN5rwEinwd27uHOcpbJU4ESsQu2pQ/1/I1elQHzCxg5d+swcOSad5z2eSvsH7
LQ7VUhHJFA6feQt0wiqacQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MfAWOdil0U5BeqG8KBiPHOpDZwXqUybhSu69bwAGXuqIM4PBnlOz9ek8h+DEGkAV
DiOPiesyjwex50iYUhkrwpxjrlpnnMeSqOMVl+n/hIjJrXv4gkz0j7OZLsw6yDOH
XVmQ5EeDCZP5UpohjPBVgEFODSFcIklPjt/R3YYNn0/A8cyJ5s6+YrV6INtzjApr
Spxj0w/HDjlA/Addok41oxP1pj9zDCgXXtn7MSfejWl0XUFho+OTPAZy0R06OzNS
CA2NfgcnO9XX5aCFqHJSFQ5yns5Jt9C2RajgWuW9sez9iCZcbqtr0nzAvs9jjQ/w
mS0Fvn1wdZCmkKpq3TJYckT1YlV8Ehq3h6jpq47o20AqgwOMexNJj1Mi1P3XQr0q
+s0lM1J0w1g7kxJKnUBzou2pRHBbltemxSb/pXbZPxc4GZFIfS6yEimo2MTVhGYG
oLr1KuCMHo8R98hfw+wuWKV9fHHictEfid5a41vA/sEtNcdO9sbVzGwOd6i0F16B
+Six2QgSIRXAV9rHX4ohSghdDp3OruVSrbiPl9wAQztyBewC4raN2mnHeZXunUNR
/8Jo5I7CnhFQoExpiIV2MDzDJArWY4wkc1AAkEnnavjv7TkhOZQ12PCn/0gloQPd
AKSd+Yv/PoKwBd1PTfOifaf8TGh9GPrv1ZpFTHjarOSqHO2aqDzaFaLsqNuoXdfb
xpP2usxFdkZZG1UHy8JQdtsKA8yqOJmXueYX+0laV/fsTOR73nLHK4su5CuQBvqA
W+353QKD1AeuOwvE0tOyCykGTpyIXvtD+Qkl+dO0BHbDkHRRZ44MX/aIz3Kj+/Xb
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kaLaP3uh57owBYFLNfD6oTXU/DrMQaxnoaoL2Epfpy97f+xjRNyOz+H3AV5Ew+65
9VTLTMsl4jEXz7dZK/qEVLIbONmYWjBzYCsqgeeTc2D8bXgMHJQqBQX6awbBitip
xa+S1xRX2wOeMYuxQP2Mzf2lEhyykxlgCRshsw+9YEjmlAlgMrX5h3QR7xPjMo7u
A5HBu2gVc8syZzvc3by5GE59sbGmidB8ql3zPMsHkZ+rS6jrRSelzFVhMLkfOklQ
Z0irI7E9GTkwPhM/ZC5QrflEa96Eo0rNKOk/KLd0v4hkVE3WHRs9FNAOIsgd6y5Y
D8tL+cyw31Syt1QdcrRjpp3ghZtLjaVe2vhsMEvSL8cJ1HKSCNpHizriCyc2RZay
Ev1ApmpAvsIoQDyBYWpNg+28b3vYS/ygwobr3Z2TVN4z6QHxETKwfObf2iQCGqZ+
xzHPR5JEtcQZi5YAxbqs3faneu6LRTsq70Hk2Gr4xMX24e/qjy7HYxjGYFkOmHMf
TDI4t97T/69kymNsumjlopNy/cXaWOGmrz23qGMRJPlc9yDB+bymBQlwbxYteLMh
jsbBCuzuXedBbBgARGgCWMDehdHXqs7LmIEeXCEhtMfKlDXG7EuEF/jyjvpUgu1r
aXdHKMS7JTSUO5tBU5bycveF4zMS/fK6v9V/4pY62Q/3+y0gNMymLXFKrSFcTsz4
HCrfnMGwQGl2KsjoRjNzuSMLRqu6ybkw7YFwwyI9BFkBfWmuGobz4xi0wQPCAv7b
m0qiH1pSoBOo3fzQqLCL6o72y9C/6k0Pw1eaVjQBiVTKlVFsXWOOqfypw6ch83Sd
T6n8YjFWgo/AT7CaNqReKiTZUPpi5M1gXdhLN46E80HdbxsGxdlPmW/1D4Dmov90
oCRFEvfvCznX9yfzAeLGfE/0p2F/JRlQ1fGSFErRRSBaMKOiIx897sh910wheBFF
hdL9fAGy2Tk3ex8knTzQxoyPQqvcjHif/NklTMtz4fUE36cLyT9s2tXjSGYBcSWK
H04bXqwrUmxKwTYCl+45UsKvJGN+IXUwAu4Y+MbjpJYc+AwWdTzCHesnsE6eG3dP
wvaF7hpES2UB0zyp6MM43pRjAG+zWR2cuG6PJvZz0nFyH8GeU0OfHtcnfYaPy0c1
xR6Gc7lS4Gy/uni2th3tdzL2nv3hSUqipHpPYHadzqPGoDupEwwURYnF+aFc5EsT
P4YE3lSL0he+XaIDf7k3D9n+fYECZpPGlCeVsHL0EYf8koSZ+6esl7emjw14C7fo
k5F+OkZ/5HOgUNjQIJy8jHDn5LjLo5xCkWiZ7t7oXCQf5tPoItflnN+I1x+rKIVW
Ay0FcyPiWAOz0IkhWXStN2CWDwqzBadqAuVxJzJZWfn9N5sNWCn1ICeRL+Nsjy/0
c7clr+8OZ/DNpYkwUHk9doriYLyUwdMBGvQJ5kS/3Z+QfZEks9eKwlVkMhRzP1cg
F3qOfrUX3T2q76G3TimqQkb+87o8OLMpe4glttjh2JtWP+NyN1VFO8yc28p2TnkD
RelWQ9lvjsBol0e6JnvlAlv4LiGvRQJcTsnUUL/bW59b+OJ1cff6zZJsm8OAB3uq
aeqpTHLKVTvAnS2XmuCISclYkvdq9QOtID5sYw/Jt51V7so/UqxMlK8BAxC0ytH1
xgt7iGVNUvhIN/9BkcX2TE+wu64Qfq55nrD/vi2aOeUAoT9ZdeRFDYixfEN/F2+s
GvNSxLLp1JVfa8xMaxlxvk+nkuZ8GAcjgVITlUTb86eqlVe4AW2dBlXvyLTpg+wd
zNvHSWhSjSsX3fGVqykdnnbeZ3WSSbLUa+B+1Wv4D3usVdMtT+fbykGmJvpZgK6F
xXC6MjIxfSm/rrLk2UuvJZifBTxJ2gINEWyIPLVMgiSkHxfqNUQoOxEgH+Jrv25D
FjzoB4GZyTcmZOdBi9uS7619KBH5R8b6WHSL8PvSiMMeC/rYUlwhKlhD8wvzxKAP
4mRlrU8/cSptIuA5hf+nN4iQE+GhBHwVQPyMmL0lb8/TVaWiM2f5BltcyLi4OI4F
J8wbYq2DtQErKObhFyCNo6IFLEV8dqagSqnExTt17DJ2ndbGTDmFIxYMQ0PvTDWf
LPVll+IA5DOXqekCmKBUa2PH8UilXrSRYkpi51MkRhVqHQk9YHbN6vdZL3JRo80x
I7DuxXrKq+kHcT3wkgHvbsZ76kSMuTVvH4M+sKrCYHjOSqFfZIdPS0gZSSBJglh9
EgF3kDFpq6/NDwpAoHYJX70srOeZ0+T3cMetuh4TDMjWKA24nUGY8fN+JXlw2si8
F83R7A7TXgNhRSuTcJeJeZn7Q3JG8eA2nK8bC91EF2L7OUulfhBoWIxuzYdZy9YQ
2G2W8vHyQMG6n0H4Pz688g==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ySjBgQYPwaummac89u7AZdKy6g/YyrjpEJif5BKB66SFuMcs048b1aarqUgPUcFY
FfQKRJVW97TK16k0fmvJRRKp0i1SLjLNy484EjbpHM7NDSvyxvtNJhsCOI4/fbiP
QEt7PYbnPsYzZ5EIRUMAvrzSq5LjRh2igOA2S7tz+/8xYgAaKbh3U98ZP1qDzIwg
ULxxIEyQXdb124RadD77QRsGWU9CohcSHk1+ZVu4IvZTtpe9jRRfwhCtMWbs4t64
eIAOTD30dcjA+iVyaBLNbKl+YNQfSDZO/AnZnDEcDGjuFWS3hzi6FeTD9W4DeBJZ
KeLYINyqSsPIg0WvxcTTKYglgL+UZK4kphlYlHt9Qr4GhbZE5uJEAkCKFNgnh5sR
gBPoUms2T+/FduXbFbFDZWblQrqRS5lpWVDo4BsgiDkFT0qP3Zbmm6jlNQaA+5QI
+7GyWPAXaxPb+1/qurOMSId+J4w4t4Os0MO9rE6w0t6UpWabFi4pDI7S5H3YYfvC
Ru0JW1tFnb71RKk0aIGONvr2jFmKILfX0CSojteV+6lD/88bzYtcTWDjXklsilzw
VWoPWnoQ9lhqSMT0pdt+sO2RpDkqcstocDOr8eAUW5WOiEYEWZ/YrMeD+oxnCRgA
+Im/bCuzwy3DvoXvMYwJ/LinaP0+UBRsVJ/nnClFwKeX/dgivZnX6t5k8sv2xG1h
RTp0ES35gQ5GEQeythIdomu7ilHMR1KdN9orA/nJfUPljI8zuH6gZB2JhH9d4o0h
UQD5dCI3Icc9LwFo0O2ld6niwN+fV2gRwlCxCvydMmxm+Tffjjd1iJW8FOe60tE2
XUE7JeMibKxxJisU64Ant8Zu6T2Gx49N3uCkTNWFaHHdU67fa8zKet8n8gLzlk4/
uE3ugfGOwuiZgqiGXmdpAOpMrVGVAAV8NvmEAx5a7fVbMzbmXuRRTLKwyjh6HmCP
EWHi46qBWfnSL1tHi14BG98WukUVclYjWYHw1ofnDrjKJhqpWcWXxRhilSPReza8
SXn8PewSbWSottkSfKGa6TNP6ko7MWnlv0y2jUUoqtkIA7uSUX4Qfd3YUKdErKrY
3wmzRCGnnUy4aR10FebRwEhg9N3zO67Vn2Rl564tOx39cfGCWSHRxWwcI29Lm5IP
qbkjkXTejpLTImTcO3glIbxDq4Pvgm92sDpeaIFyqeWw/7vgohnSso4MTZn5DM/Q
lcHaI1vAsGWHJfCqMPvhL5SzUmjAIItO+BlU79ws93c7WQI4hT/euI2eKUVPGP8+
NI/rZux/Cu7Ytt3Wp6TNPXq1K578lDQTlYsz9X8JZmRLu9TnIhz8HxBnz8mLAVBR
8a7P54BDM5zh0ty5eBmlwwODlcqONN8yjNQfEc0wsy/G9JbtkFjIKV7xMKMxAZYJ
zkY19sULnCRecDRRVg9KsgeJU/SNixucBR5N8VlsFq9AdUnficJbE7wdFxyY0KAv
PDUwe9yIP4cQOED2vBM6btvg/ynyiSm/2nchtd67skKVJiAqUBH19GYXZQ6Vyy2H
Z/0iyo8S5fgZ+Mg9/zyjH7x986l6NWgQoRu53yJ+2OyvMzNrZpNq9b15AYQf09tn
oMWTV76H02OGlaW3RId8tB3dyp5KjRY63inSLNF6jzRqtFlc9ygGwiV7IyOkse5n
XYprn6e8JTaqxEkfQC6rWLTzIn9Lev/rznS8+IRQo3c66LCSMG5bksdPP3PQ5mKp
zkZvzxgAgsodAnqvX02rg52w4OSKwOB6ttLEGewNyC60iNOkIzUxvh6ynVYfbdSs
soDOrcVS21Xo/H3Q1YbV51YGtPzz8iyeheei/j6pU0LW+F79UdypY1pQubhvlhoj
aKBoFf6bevygKZIGHCvxzw==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NA/nPvzYGGn0GpP9WBB77oyqSVjYkN+q2bNBxLqaPVjYnpwpdK5YzbillPEoezVs
fLdy7Z4RFDrmnZfJaBsvFVue1jVj9xeePjysmaN1VgRZH6BgYXgXtCzL7AuVC2DA
l7fE388FRgMvx6du7gX2Q4iBPigNEzLwOMVz1kOsgUwytfhsJRuZ2bH2S2jnvAYJ
tsBiNJehHv9Dt7jS5y7nthALoYMIOGGCDUH2ql9fBdBmeuJeebzH4dfjtN5W0G3l
PoozweqipvXy2h5NQQv7xRzFikS4D4qxch0psAtIRRyaRM/KpvXQVj9PSp41YjT5
LMGcrQmPMMsBPUp9ghVmKePyZM8hIYOCXiK7hv00eifvcc8AGi3NF7e/drz3gCLz
Q5qeKFoHOnw3eS/HSzZgV4yS0nPZP+074HzxjNqqAGQFxYpd7pth0FdI3ght5ehD
OTQeu0dSYC+U9yt9AuXAPL6CTaSdonJFeme1BcDyHBaO3AQMav6coAABksYSCvQv
ni5cPu9YAaEmIbsBZ79R+htehwDX+Kknw+1NrcEMFplsYWhs/QfVpQNdHHwS2mW6
6mfDSnXsUl0rXDMzq7Brd1msz4GcbZ7PV643a3CXl2zD1DvBbvlvX628mwbwfk2o
fIoj8icV/jtkfGaXwJ19ESkBIWf3mxb9osecsm6qDtdMrM84LVZRfHUVFPBJ/MoC
8zpKIXafjd06zQnuNZHOoy6TLqh2dFOhG8n+vedbFGNJjRMLId4Ie42lidIyO7ok
ipg3ue40ZZin2ObJindDFEeBRIECTJjR0QZVB49YDRL/OsAoX7WSZmIl28IXMLxB
ByZLfFscNWZIBtsFdu82CCYGiB2WOi6fwk8wh6LKmlgqTCFR8ee1NzE5BEJLe4UQ
xCNTtvcjOjEw18jTybUFGWKyb1zfVXc5v1DX9oo7dBX0wdo7sKOuZZEKTHXF1/sS
qrKS5soN3FEF5EmTABl8v4APvPa1PnPzIPYbFDGum2TLiDHtpUb0NnOSY6ZURNG5
pZY4PVg7rzt0OhP7M3tlsEoJ2ZBR0eDhaBxG9vAzKPUvMZ8ifFlrn+F/kbNQ0YXO
FLrYQnAvoB8y9iIs/92Qo8C1Iln1WMuJlzrFhkXihdtGGPNmOCPv1dPWDRPBQDIW
O8a37XTrdQi98Sm1kXU/92P9Kc4AlFuP8OhoAPdgqzMLt2mInQy8rC5gFoCAY37X
vOLB/rZ4mmrXPNJqvT4ARd1E8snp1EUOvm9xhxk7//Nx6INK2da8F0tWpNrhBQPX
Uut8W1PnQwWREx+8Znm+tL1T8NP1Jq9Iy67Yh+I5by6BhZ+upeQ736fFhwCfHze3
bmoPSgfwOk0rXlilFjWisiLlTfdCQUdKeqntOOHW4Ys1UUh20QjvH+3M1/4nqdya
u/DEAvbXK0157cR+Ho9PL6kZe9xhGk++DGL8Z0x3TbtkxUpBtlfeUYCHUHF6TQ9V
LJ2EL0GhwRLj9AX7O2Gwg2+wzeMmMi1JwJ/rImAqja4E5eZMIqBXgDijZ84JBiAz
I3/9q0XH0Z67WCrI1s8/hqf92IhB81N4rPvGsyPW1f7FS9CZ1pKu+tNM5AXVdJc2
8SqXlflXIsgmtlq41dsZGABwygf5FyuY5lY5w4QikvSQ0jK43WTiyguZNo3AqcfD
+5NqldDYRN7hDcqQag+pq1FgwaN18W9hwNyfGgyYKjLUjG3RbKEISipg1vcIbdqa
FGtYJQXTqlbS8Ys500Z9wWy0NtYeavxl+vBII5zpY8G4DlcT6lAR3mZOFmF/bEXc
X5pzaCf0+Rf/hbu0XX48QgHdKCQw4ox8ev8m3EXt2gKs8RroDoc/urTcV26v+MU2
E30WgR4JCoZpbPHG6OHjO407z4fBzl29O5J93hN8gYx0RLzyLRL7W/nicxR6lufG
HtQnDTRN0tbkvLydwtO4Orobn6W2YLy9518DUNpDC6eu2y56Ac2r0dF0NQvucJCf
TEar1/TFGti9imhjF5O6t8nf+SvVSPEaIeaqLXqLTOldttS1lS5oLFgIuqhoT1cY
64TsgpHRSd17MeCAGyPFb67TGNkLcpL+H/ekN+ojnSZtQD9gwftktP6P5vyxlC/p
HZz4w99uZkGgLPthEwjTbDsXAOT8u+ytdu4pJ0xsKjqAWoGyjKQaQFIZVhfFl1T5
RldpXPcrzZ92DYSdyLmcfETIvje8Z+OeNx79jgxKeWj0kpLeZoUOioKwXJIHJNsp
uqpLQ3fEWwKhFGCQnfpXsjlonir5gE3K7i7sHcfXBxaEpp7jajHRlUZANZeboCMM
vAWq0/10WpmKHPHHyD70ahLblYYi9C7eD5GvqPNvEkKd5D4X6eT9JIEjOqCia8D9
Kz7Ifw91fDDqvDgHmBCW6JAMFh9wz2Ei5O22Ii3I2154QSYl3iOO1K58tuGLj8mc
CaWjzboQSWvuqhUdsoJe5yoJJbcMfWcg/ToSui3dMzasKJkbinGpQP1emFu+LYV8
IqcxJ6AFFxCR2H14JQxKYE0thcWZwgjnyuDQCO8dbu0umm0mRHguNmfp1i0Btq1q
BcVYxxpZ3Lr5UBJyQnGqIzxbqgsBZZVizQh9sTUuV2WdSW5YxwpcUkn+p4L5AcQ3
6zZtaEeX2ERioUXbIUo50r2TDzmG4YnwvikWaeN/uJVK7Hy9s6CrxmgwCa/QWO+x
xAj4cO0c42+PbrBDYarK7FLhm68RUBnGXIpnXJ8ljxVVRZs9469vI493YxwAP96s
Idorh60WkSsbWaPZDB/QuV6ftvo3wdnkYk9OPUJ7mpVgPy0QBhI/pw1JXSAqfsWA
+8+svxDUm7tpsHJeSWI6VdObLOQbUbVarvWSOEYxpph8+gNQPFp1eo2iishn1gUX
DYjKwTN9RLXpZ80bNs0SAClI/vpW+8qOc8kzPXXf4/eYGEMqq1yOv4259megeyxP
bCbnn35AOMmY0rPS17ewks/m5NPkR4MEthcQvrNQ03vJs3k/z1KR9TAcdQkkDJoZ
toFw6FTEvPuDWMh7pR2KN5cMnUaMeqqfQzrKsbALUftZh66dvomI0P7QKb45033g
c5mmAZ2s7DOZl7Csav5Unlzo5aMuLJZlbQtjvOxkIFNCJUQFFfdIeDYF4o1wgkEA
Ils66xrF2YIwEY++T5ZkPYNGlq3g1SrVy/GoyWjsgraRvckv8BAlt/tJwx8lxow0
8U7JQoyjVCLPFI6vXaFM4m8QEBVh8CQ1EMaftXsNceD18sR2PiQmY23FaVkOFUEC
YONoViXu4Mg0HE9a7h6gU8nXUJm6twQSX6yM7gZqtlgJubNpYlNKGQpt92iyvclr
OqaQYU9j2/Qt9VdPVQck9EJFML2lS/FxVyz48qIA+HBa/k/EQJFxscS8BfOhgyot
k9rOtgy6i/X8nxibhRBja/O+zLMtp6jp4xCBiMrNyufEs1JWVAPXKC4Sw9RUCqjQ
91zsAWh4j2qT1K8WMeI5BHw8+x6KkGnjKqRObJwtqT4pvwwvMJp/y8dGneWojIHs
0UduZ4fTU4Mx5Cz4NasVwUn9NDuFNFZX+kJBWAa8jhBAS8F5upR7DJZJD/0qABzq
GjVJ352HzOKVneQr/Th03ctcqPHcJYhfR5SPnpYcxRxG/6I7PEFjJRuwQgksoySq
xYU8e6HTmT2AuRT3+GKVGZhNv/IbK4vQKu4ErCrzR8KoD+RGngCIYSlYSKhIycDD
wBnIn8D/kMI+F4NBP/eG3rWGS3+ONZZef+hyJYLncxXcx74xStDgQCvV5kE44QxY
1ba68g8uI1kRsiICEwwfI6HMmcQYIj21uV+pYwMaOgB6moMdKF0X4b9Ruccmev7C
8157Kqyxjh5KLkkeSUqUrF/4bCCl8P0DoihbG6QeAyS9rqrzwDLSrkTB3qXORhh/
0gLda6txvbOxkhCOBYv8W2k0LlDapRr4pi/Nr3QOhNIhyw70VMuWJK/cDJ78FeRj
g3qk9klGvNNX2xU8o1Z7m8WJAMN2yNDoZUJLZGbvsKw3kIaeiQpVzpAmqBtCp/WP
vLJvSXx8W2ZSoS97Lc/bMbYsVsJhr7tPz7jKS+nDCevIafhzU4x4F3ZEDfEbafb0
qkSr2y8w7i1rPRHchyl5cws/BDnUjI8xZv2NlhPZNPpeJMzhPEaWvMmBZkRkR4xG
nGrXSdx6xRch6KhA3AiqQTTCpPd6BrDXQWPcFBCbr3faUQOyiLYmfpzNXcPacfkk
mniUcCl0as8n62/jiIRO581ZtpaEnGARgDQr9lqek49A8ISjnmyEgftdla5VmVV+
s3WfV26Ft24QjOGOWWVu8GuLnh9efSN9uN5V07SNAJ0boem99v5+eag/MuUDtxvT
2F10oKs7OhBuXGR9YujHSzmFMp5TH3g8RamBaZQtVZQBaPec/PW3dgMY6q5fWpUk
KW80P8c7NMa/yXPvGta77ZACWkGFpTtKWbTnvHw25CdTXpgWPPEGJiFRlSe3tkgY
QC3UE9VavIE012mh8OPwqxqkwBh4Q4VzOqH7/OH4XEE15bAO3JHh8YTlzCjgmGey
2O2Zrw4pBWDBsGpB6OFEw/vy5WaMdURxXJJi34jsTBPjj2IVF27bjbz74Zt/rADx
I5V1UvjqHAC0GafjEPz8TF7Ik+Ocz2GbvzpDXGpfsD4Sz/1ovazYEcCElwpHoEAw
cAKle2xLoRkwV2kt6+Wkfv97VuF1tt9DXg62ukHahWdt7A9OrJBWY72uWaqVLujG
1sB0g0ovVdOZmagT5JmpmMXnJ/jwsInK/A4ajvJpjaj/ZFzA/7plQR95SG1Ax35l
Ch3RYIZcvb84uo50ZpZSABsCvJ8lA/F6JpjJvU9V7MMJ02/ffNY7OdMUYBIE/X8B
5NmgOSZTRFn22ltZo47Nfhxo3zxZrb+QxxkDf0HtNWYDwyiQf5r5Rthjw9h6bpjq
XduEqjU7eP1gjYdXCkrKNi0czJ0rYTACHyvm0VhJpu9ZmRY2PASWrY9C9PAlcEM/
iMkIKY9lRu4RruHqIoMUG01X5m01vVP1Ntm/aZaEXCubVV58bqgh+9s+O/q7tWwg
BdPbKNgjFDGFElOHYPcCWKiHKay+LbHV39h0MbXRb990JX+UuYH425NLF/YlTdHg
ifD8w2veHuVVekKY4Ok3KvfsNgvCB1uucNyv1mRmEVua1PyYXIF7lbEN8qGKsbvh
W6sSrnILcfEAJIvg6uhZW5YzwMQoauUhJZAU57oWLNNXGYhgqYNv7pFWTUZq9NTi
IikpKTlDJaYDDZBUgYECwkESgFwym6SwD/EDJlF4k2Q82L5nzlIt0PCUKHoheswo
m71UDafj+3lEL+FXTjXvvFhQcUKw0pCGCPKKDXn5hpNXg5J4wAkWRa0RaiYfQsrG
dU3N1zLwsq1xrlYV4CJIXxEKHwF0zsfRlZpeD1/oQNsUdAdpXy5e17QB3ejbIqzp
VLZAJgrPkLk7po8y+oSALL7Z1GGoUSQNT28JYJPhteWhFR8q5+6OfsbWO+BV2vZw
9sQTLPHqvEAj2UlyaFA8C+oa0L++nJ2Wk1sOEB2aNdjLuYUlwYolGo5GuEpIyUvA
fRfkugg3ILeIyKjG2f5iOqzLInIwAaSGyJDcnJUWial4h8urqb10m7GoP1W4fxFD
Hs1lVvs23do8zZ0YvyBEzA6c1ZLJEYipyCPoXzyBf2gM08yYhekpkwAHM14blquJ
JPYCPDxwGNSQ+cjA+CAEo5AouZUXVIJAx5n7kAqZn49fYIanVTwyACehEPLYi2BF
bzCVKt6AQzeizjm3D6Fn/a4M1kXyfHyHPWExd4IusVwCSnc9TiUwa8cZnvmGkfUc
noSQz8wViBBWoCfZ5VByAqsnWjb8yamabm1NOjO2WYblg1Xy1rY4MdxDHMDwoYF1
2ynXJP06KI68VxlPEzBpVKN1JZeohOUBygOibHOkWUHqGeqcO62DIz04DWAATN7T
Pm+lQYHBQ9SqcidOdaJzL6pDI7v4btABp2Zap1U1SvyFAzynjrrYWkb853wtyTph
ZMA3N2tctwBPpdn2AthqmQ3RkpEB81GrhkPTIhZfEyMje39D5C7Rrfr5KszmNQTb
BVKp+AFDva7RG2h9sDnlqQjcByE9/pD4bfj89fxAj3/gQoHYHPv/eZzvOygudd0C
Y1xXF1mBvZMxrIfdS6ZO7AjdJINqHQvSPA5siquTiuGoZ9gew01g3CcBUN6pFGxT
Q4f1AwM9ynHg9qUUvmUjR0tgQEga4Q0Oen9VEYNae50=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ELB7rMY9MLgjATvB3gohVzfEotX2bLrRYddTRC+87E5b/CTM6baVm5u9yh7ugzbI
hO3UuvQd1c831wzEdHVesPBiloLGiGXY0S5CQmqOxf1EbloV1wjQwMPweVkaSoUN
m22VLtHMAJsNBQ5d9kcvmH4Uo8wWYLtyRLCDLzkXYQhz6jpfxedeeguPm9qh3wSP
1PmSxln5ei15biXMmy5Ttlyt1AXE9FsQQwkbOrBMecIjOEES57aBaYPQI+w5Ql51
O5fcYcnUu5xGaRr3WJM0H9znk1YaqVAKYoMCQFHxN0JkTp7QS4qUGfqe/wBDVmwE
OBnqvKEloPOZ4s7N68NwMv8eE44sNclT0AgyAtMDA78r/Pf01+G10wpzZOg6uLgl
7GFefxg+SMUJlwrY1fQDBV/e0nXczdFi9J2Rl3CWWsyLf6k8t4o6GqKt8MmHdRUs
hLnvaxXsEgD1vPUy1eOCWQm70HqlAvLN+pFTV4yNrJzFuXnnB974dnCha3AydToK
HiROqkNc7Tn5e0NlzIR7/mNvtfArU1UhXF9gqavXY8ecuGeeTI+VEQqJpOZT2JPv
H7C1u3wDl6PBW5tf5jczKoCAZ1/QVKLO1CWm87nUxMYPCvrTmfRZ2G9qLbJl6oTY
x3WkBPyXzwvg23UTQSmgJQfWqXlsudUl6RT7trc3ZJYHdjorGwIbD8zbem4muozo
JBv9GB0AV9dTP64jfnk0SOYtJ7YVGtSah6T1an+Zn+XMBQ5gqtdbAjyWYnlrcLY2
AEU4FlDT34yjI/Cw64fXzruE3iJPHsHuvCpIIMxHEvjnrgs8K0x8lmDzddB9NAov
Zt4Xoy9BXsOGqIdPBOT/Lqpmxj8Wje/myAEvec660/WIK89XvgdH54xoJzD8+Jeg
j8ONTsZ98k34RTwUamyjfnfNkUCTV4U6X4R9nfI8L4oB7yeiSq/h2z2bXHFfqPp4
20GFjN5kTst0a2nOnB8XEnhLsVt2CxNszYniGNKkAf+iv9dUKv4L0XAgV/vdUnq/
zJmC9nQVxiGVS2Je3Gr4XEhT1MiBkAEVuuIRcSTGwOoXsEWqlOgTmazM72fJLnJ0
GE/U79tskAbGp7LEWaIFdbEiw0xobqiZLymjqtTpXXmrJXTB+H0Z1cnSRJ39UbKJ
N89GNi/kI7+igefUuWlkgdApnbASfuG04fGcrhKdqxfTZ9ysUixYueefP8Y5Y+3c
4dOLfhl7hVzeLCwTXb8i5xOzlVd+3VjmDXb7UtncKXeDj8zMflVXujeCn+X/BHvw
atofFQYfbA8T4M8dAG6dUz/FKrTm7TljfXcbMoY5SvKOdI0d2entx/eQoftuft68
6IXjhrz+5OxiyQD+Y4i1/9sZQiYXwU1qXKjUYEFU2ep0wOC/jrXU2hkrL0RovudV
9kp3fg8O8rqrECnT6smkzvk4RYk/p8xmM49ZKyxJxE3DIL7yn/PPJeCjha29pI5O
2d3khEfWYcRthCvWDqlU60apTvIFZyA0UIhzn++0k9vrAfV8NeKE4LuxWXWaoe/5
ciIEzS9qQgK1HuZNKNwI7ogpBqoAQsX4GPdznsruK87lh/mQcIm4nq8NDSvrqzFM
3HFCT6m0g0qmatXC7DMmmD0zEq7gqc2A/PSrFUCD1SDGRVcksLkSw8VacVsGcPx4
lN+x8zbiSj6Vr7Kz8urEA28rds4fYwRioPm0Cui3oCOZdbSbIbSzFBPSKo69CRk/
qmacTPkBu/Khyq45xGTKYFEPkncrWHSV9Hfb0MC3mO3Z3WX3ceVojaNiULuTXM9g
i00MrW+Kyp9QGG1nhJ7TQ2Vm7DuMYHGwy0WFqF66+AGh8dEroH49wl60wTZnWPfd
v55quD+fHAOKN99lgeEPJEU6ep+QK2/39i4YN/UJTTPNcEFTfu2DrwQ3oQ1AoE7u
FIEI63NSyPbW2MGXyMgQ9LKFDejlGku3QPPprgsG9CMgs/VNiHGS7Ofhv2FSW8DN
XA/4oy4kDetpL5l9ImT+fEghu8kMmJXBqjVO+0sHO7/e8pMPA9srWFaha/Jqxqzj
qj8hERahn+oxUSfJFkkKCv1bs8ubFIPC4F9Bvcdnav9xMoObJ6ekSgl0qJB9hl5N
5CLgo2BIO/o+yFXf0YfSu374Ioh88ZBaNBQs0E3BBd34+MTutT7LC5od7dWkmNon
UDLWWyigzp9D45gd/MIrialZ0n877CfHkhaMtudKYV4RXiw8oBu02tTX2GKR6S1m
OTom/rQ+yfvwPSjATfPMZWpm3wkb1G3EUie4NCFs9JxfTPNclejf+EcQWVxlf701
N8rkiV0GtkfBC+FARE5qbTgvU0NvybrnbWgp+jWUMDp3mYmx+3S4cfM/RpnpdgPj
T+efKENKxJIrTktM9dFZPcAFR+DGgcazl0Up+cou9iX2dm+tRE5ERwTJOpDSU/5I
vKG44+o83f5UjnLwalVIKqdGaL4zuiARnR1m1fj9Qx38q2bUdzb+Wcac38ecrAUk
NJzByuW633aqHLnGXT90r5Wq0/RmSL8rA1vrvAZ8E1SQrzv4G6tjQsy4xLzSH0Qo
Un7Pe4unVHiGM9KGEfO8gMIWNmB1/DBXN6f2t0+LXJREt5pPA4yNSufvUdEbKZRS
PkmMuwTa0B1l7gWDFb+13vPgj4v5GYW0ztepyH1qlS1M7DnBwLA6uiLPRklLMDJt
CqUlvE7swiYnW7HR+aWQVoU0Mz1eUHt9TBIodAXghNOyhYCauDrkBvDcP7IEEpHO
UpLEVtwnlao0iXNGF/joSJFkd3SLHCTQkmY7KVe/vxmlAgxYQUFUFREEauOKUnU9
ai6uyIqtWuCIpLHAoeuQ/Vyg2TdObrKepmUfJ/G20yv0GZ0jRXySPrAUCP5fe95+
4MWkDwMf7mTfhS1Vj8EyL05S6j32BR1mIrpU0UGSu14p49glP09BonAQ6myPla70
lyY6zJ7fwYqIU7k/3/ZmtLo13Ei1Q+YLq46oizmapJCIJ/Xlp4pdZh0I/w79hywt
`protect END_PROTECTED

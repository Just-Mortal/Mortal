`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQb2RNxtkofwLVB+zt11LUXPXjUcA0RTp1VNxx6m6z3+yCTvev3FbDf2OhmRxwK/
+djOr1Q+LyzebgdLoWB3mYo/FxhN2KCjK9jl6JJI5aqHUOR7x9wgHFw+trhkW4SV
rX3r+dCKdxNSnEsM2JeSGtQTez1w2O747XsFK0Ff8d8q5J+9BDL6fTQftgzcOAKu
t0PCt2CmraIubzglaFWnvYgbX4+B4Nh1D6UQ2am6su++IdJDnEUwSU6Bv9C97H0i
0Ggb7vJZgkEBpogi712Ai8EFFODlrpit3qndnZeG3W0FzlyfFFRHiop1zXoDCmUd
vAYiv02tx6GqskLliThQmT8kmmp9EhWsMvBVKRvt5UP5iSiXhykah5yNmB9Drh0B
Hh4P8ZZ6GBu9k6gxDSqXD07I6jK3ad3lZ53mE36SkOEWb41wLmx0xDGxmKQyVP8l
pbUmDjKZzPDtme8AgaXzV0hqhRduBRZuJMlIaiKKYozikpj00ialo2Nt6+ZHa2l8
4OH9Js+xo32/9FkQKCFHr1omQT7JgXVavxGmuIAOA/g9VkuB75jovSCS48TVaNIY
0O1GPh2SxYLMklrz6Pq5TQMLbyqanEPWx6TJi4CGExY+MSKxroaQJJe/UAY8LErh
0iI9jlqAYYIqaGnrhGNB7t2Qy9g2SE5606l0yKf5OsdD+qUmnsDsKQ+PJW22urJa
px2TtcdcKQOyBFy6gQJMr5YqjCoXW7VWCqj/IswUzrtMkP07fhDSiaAiKcT65tzv
O2T97B4LNBukTbivOeU17XtCw7tSEN+3mvxmiIblMYXlD/YOqnXrIgVHrw4PtNuB
viq4YAiSJJY9n+rGPhDl+UUfng8e6LKCnIEG7jk59LgcouLkvMFRZ1TF3xpGa/kn
fikQNiifLew9jBOt1afg373+kfkJJL744EUNZ5o/DiWP31wE4oV87xmPWF9twMo+
eI9LQ5lciHxVxhFv1DsHhyqOFU9rEKpDFRDWP5l12b+JRbvKIe3hHOm8+Mbtn/BV
ODGx18jVQHfl6hwCW+xPRQ==
`protect END_PROTECTED

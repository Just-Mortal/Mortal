`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yAR/II1kvaKuci0vH249EUbHs+1phfUqzfGhc3lSQ8USZfbCDPBhL7qUVPDkivGR
Pb4SOVp5tYWpluEUvVaVMFCi7f53iTyLWxyenNXv991HLFhFIKm2u2LlI1p9/ajV
J2ldRg9iLdUzZ0RKCAzdSnjewKqK70L0Y66JjyXg62qcZxBuxIMdMbllzgeJL7rx
f067lw8mp/kgVEptfE4JG8rIubKpJxhfffrSdp/qIeqLu+qMcTIc/PgJAZpNx4EA
ir8znWiRvZXhYCUWleLq0dJteSFkQ/gsGqAyjCOGr+t9J3WeX/2i/Ylfi2Lp8md7
GSGd0GWulcPwPFvFVWDeZyvVV7BnucEPU6owHniWTWfL8Q/osX14hfTv9S3GMVux
IbftsJ9RQisP3Je9kbTpr8rw4omT8ruT+32f5UA+TWvcn7K6q/hiKSeqnZnOvL2q
PIytMmgaoMHnIzua4FvBhaSGURWYubjBU+Ik2BPxItaBa/zBL4iXisbkhNIyKugq
OXKH1GVirDYmH4zRSdgiz8bkzzeberau0B1568opVfRLO/MvkbqKJp0lilwxt6u5
ZeuD1WwSmRVKRqubbzQ+m2RKWVnM2g1A4v4jXfV7cRdVkCR4VcwEioITfdXvV75Y
LzmSGx450IJIQmyNfLQ7VBOCi9oFiE3uQZsLmUfBDlixuESLdUav/sdmbH14Z6fu
33UrUrpkZaR5jdiFa/2a9RpujX4XNF6Jr5R1p1BiFfDZ6uldVYYq+l60WAI4t7T4
J+x1IOR5W7r8QDdEwcEgNx9dDSqaaNRtwc6fO/4ksCGn5vEgyQEU4pp/phfcv6Nm
1m8UO/ldAYgPUMK6LiB1YiEZS+aSXB2nWRM18CXE2pEWqrkj93jvuuPr5y5vuTDt
dT33fP6V5kIPFp6gZZEzIz+D8Vq6Xpc2MY7/jB7gvs+w3TnHc0iuV1nbEriE1hOL
6zihy/7x2Wj+85iD17jHno/1HbgazBEiPzg8yXvYhM8Emg3u8d009HU8ZiEnw+Cm
56Fh1+HC9VPKR56hOsHtBO0lSGJqOZR1DNxckxntiX0l0WGHEl+YmOxVzwsiuz1r
MKkvaQ/HWYyNwpaZNBYHQfV5zl6ebww69Ic39ubNnwl2Q675P8wd+OmkmuI6B5L4
w1VB7ssdIBvbfU/qJxiHVCjeMHH7qU9lzRYpI/ANh4H/tixQgmLGQW7n6E6wiWF7
KMVRtY0gdyc6BPl748CUaiUtbgF6l3CfSgUHUuGE0M4jhh7g+a5cjFJ8jK98hB9h
lSuqHYc8YYJnVhE5NCVJsd5kO5b8nrR6zy3u5XqXIQtJYE13Xo8FDXGI13lFdWOs
LehauKcMOkjV6lfXf5VtPRird0Vhel0GQJBSYD5D70RewyVaPhfQy92KW0PP/6uF
jHh5WWbSbTe/M9Ad7zUm0raJZjx5xOF2X0llpeQliZGL4K2pTpi50gHe+PnS0/ur
Wv1oZwMBox4N/LyRJBLICxY/JqsncbYHSm0lOdYC6P4gYPvsK5BW2aZZzbNDHb0Z
feas8autpl5DwZfKzdmKzDZIe0bpBzZL0cm4wC1eHnER2AkyBMhPqIvzMCPDz2IJ
JOAhFr0QxAT7iDA9sxUm41V9t8ZXtA8df6Jenn+G1AMBqxOoTlROasRvUym/aJtq
eyGmBj2XMj6r0VzD/vwwD1mmsyyB9eZOvfNZr/iP1IoU9Q2GjOczIVGaHThzF1u/
voW90J/2Y1/tY263vJvCQgdXhnoUHO+dgTfFjIXfpetKqQk7r/J3B5PO9RCD99f2
tbp7o/leB1xTs+dU+YMpvtkaNwnTkH/NuKndrcdoH/P7gQqLIfHrmAfrkq10xsqs
6v8tvS9HqEEp1qdnO78XFO7kNRJ+N5Zh8jJsP4yxRG5cXSqyLjHuLTTUXqHVESq/
seg93dMf+OOg2JsJj4oXTH4npXXaIe/34qnHTNI7wQjM5Z4ecl0FDCmnFRoNL9gO
td9FiPAhsp39M1GQj+cYhReXgu1s84WVKA1udsQOmpHBh2CNO5TgfWhQ8QptJw4E
O4jmiGMOzmc80T871JVJy36ygy5ZSuZcRiPPskRggNAoCaESNFWqzdeQGVy2LKSw
cEuwpwi8KsZhfliYBZbQVGmQ4Nae16GXW3b2rg7LFs5tBzbVMxFgUsB41FpxsAmR
4vPvWfoFO+jiWEGMWc5/K9HY8F2pne8IKUV2DZNdmPqh6C+/MgqpbPsPJEGFuPAP
/b3KUX1Yc26YKDDL95LKDftSAFLHRjrpi1oilUos1MtSHy36PtfxT0nslbJhBIC/
Msc6lYcEqPX+vsq9kpyroF+Lef03Z1TKelqt5CyR+FSTdThLygLX2L2nm3KiKVF8
+JTNxu1wpT16jgKhQW5bvHq10dNMND7yvumTiFpPC/Bbq/JbHppT4paqKf0OAZhi
oSHTG7fMSe8LsHlvQEMYtJXhx9e0PcYrTttu+pA9zR3N50322QWs3mzW4hQVoweg
BSp1QsNL5V5K7lIbrUajcUIajAbrQgatyzZJejKnQJTlJkul31xBVWxlKdxI5jlT
y8jjvDhOQJcZaT1Nexy6FuzFcEkJuhG7Bb6ktvUttQhEFNyt35DR5c+bw1g37Jub
heqh5EzahRM44DsCbkpLStEuRbhU33c3XsNwL2PTWYU1hmL4g02Fst4k57e2fzDZ
mwHartoTjSG5R7uwrRn0j3DnEY59FZRMYVARYkR4snjwvPq2hrZ7+TFgUO53btFo
ns/VZDh2WEsjyum0kmtb6KdbBGrvlpCuKdBDjqK6LVdI/JWRbJksxi+xYtSdq42K
BKLf8ntbvw2SCbs50SJB3X82bB8ObLX1+pd/kf8pgXK4kO3/0NnczKhjE+xUVY1f
yMUgX9cFuDH3odW8Ap5YyNxjQZHya0i6vjmXoN+sHZ9vAm+BpgGKCWREC+4ReNs4
T05911O9bpkwfZUIT2oIk/gm8VG4xZ6EfcubKV8Glprn3INe1BuTogsK9RcY5O9A
7+y+zbZBmEI6QHL9yfuv7gZjnnN5UfLYMX2xX4nOgl6T7w2+nsZFi3Ke1zPmSOhA
OmGpwThIYZP+FlbKDr6O0Y7kra4Qiq6qj52eiH0/psaRVDYLN3gceDUd4Xh7gatN
ODTDi0M2xF2AajIs1/gTtdqBvZKHNqb+UBgiECzyhMwdRgo+BuW+gAVCVXWP+uG0
QHs29KBH0pmgirl4vfypKTYQ56bOYkaDSvVKlt2X7vokWhyhuXoIxtViAqhXJM2F
v+5RJBZBRCLwrZhKsC4NWEn7iRmkne5dyFUAKCBJ7Kl2v7RQZinAhQRodP7/rFSo
ALixS4dwmRiCN8JSWnNuTsYzgWYLurRJ2S6IeYKZ65D/w0o4kjDguKIZTQ8KQNWr
mxJV9trfgKNsCS8ONerm/pS6LKk8acII/Znc/Q4qXrWvONPtSENPCIfqawksaQ3s
AO+PXMzl1anfV1OOcCQdmC8O02bb+hJtcRM94fciV5bl2KCAtqFc+TpzbCBROVaJ
mh2bnvqw07kHfoBCs3Gv1zT1eiBUEp2bjikc+f7txvXiRBR755TtX2ibSwWkPAdy
VUQkhYWoXoyxw5gLiBD0MC6GKcWkFtWbYX9kfv4n5ISvnTlgAbtSh/dXXX8Hafiu
lgRcnU2XzRxc2RX4Bmx5fvJscY6EHEdU7nl5/nGrHdlZaIjIDFW93NvQDxwrA1Pf
psIZ3mxXz2CPvTlmv0RZ8hjCvhO4NdmbqnBqKctOHUoZwNUQUtB9FycAXRX4LzdK
44OydxdTM4HnUq7uJRjEz9zzL+xuQ5bPHTnUnavtNgC/+D/SCcpb0nXdoY9OABNL
vtBZRuBm+OrlWCAIlM3Utn4BCwaIjkfm9Eqzk7KZEqPs0CKaopbm4xsLsHKd7cvU
1RMXM7DmzOhAmH5hul/IdreCB4ud1pAjX+/ij/DPwHqqSbBuxSkEi101z43cuQk7
hVMWA3CR4tFoGCYcr6B/V6xOgyO32+5D50FBuWSAykWXbA48uCBUdkYZcpZBH/8l
HGsln6wdZK5g6xC74iPtvFeqzBwIFCQ4UPx5f7ZbklRPKrgYBrVvBni3OO6vRHvn
j36pBOkDPJ1NgYA29A0RBNEOcG1IpXc0LFTrKkZOArmcufJbgWLfPeuYr5aEm9Ht
ZcmLo26EUSdwcXxdsUmEf19WxlZ0Ju8qN7X8oktR3tTMzuwxOmd/AQrrswrGLV2G
MjJtRzLBDv4BMGV/aO44faNY52Up64vrZTZG2alvAmERgh2UHkgLBEcoJzWOk48i
AvDtRqiORumLb1I4L5TKE34INKFAxy95YzYYKHLoq8Z5flw8W6Y3XTRlZjjOYYEl
dOPn+DBHxFAE7z2dNPwoVhl13CmnWF6XY/Je5pAmf6BNy4JHaHKmfyHkj9gpVCs/
o+jqWh3HSO4bFbpr2/ODDwILxd+f6Y38WlIJGGHfWRp9TH9qqPJnMNhvLcDYp1Hu
LcdIajA5tUvSZ8Jf/qAiPt1fYwkBgfx+lshGmCTrHI9HpbwBp0yMQLpXoVk25gSI
kC1d0yqm9IA0q/Qt1POv+pT0E2iez04RNihFcaa6V6Thqu1xk6aF9IWCaZqQzzT6
hnujm3oHM/W81txg0NmG/tUbNpjx6IyznF/Vyoh9GhKL2B1L/8oKhNiZkkkmvLwk
Lt10JRoCg8JJgU0rf1dkBZSt68k4joJ22Lh7zUnp1Bu9ZhJBcjka3WQuCqp1MBcB
e32WLUYeFk/6PNzg12F8ckDmyFGtkeuG31RULRDw+wcXFyrcY6f0GcWc1vo/AdGa
yXaEv3b+ugqRHDE0gkDXP8rK6gDxJ1HvqtjB+/qcV8D9uEGIJUP86pGDjWlTZDzG
k38B5RUULMCPTaAMVy7ZCflITFwh8OwEsNSkFp88O9eDxxFkvB1zBfia5sUEMKhN
MoB0Bc2pHDCeb9SFAnxcdGQMTr7nVHIJqVTV53yzPa68j6H71OYd+1r1y59bGS3V
OPD70Rwmn5QZ/jA4Uw2hMbao2v2JkXtTNUD7eivIIt/Qwtc07tMFZiWDkve27Nuq
gDozFN3ICfsTuSvN985nQoJsCflmt7L83eLgL1Qw3BzPUkqt243twb/SqIte1ld5
xq/QNOvKJy60GK6pxKtV0oZcn2i06bsAxONLo2yr1KBcS/ltH+klBwjop9pkrJMc
pDjr3BTyxsLdMdB22CA9G1JcDaCJGd/M2moi2Lg+UkxThLXvb/96CsoN35Ik1L5w
JmSuSJboobarrvo+sWKuAyARqhApNTPcJCSapSXBzYGJ9x4grdZ5w1mV5sTf37Ni
xRQEOGu9E04+dLetXOhBE4aIXZ1jc6ssEwD94EmWMzyPgYGp5Jbm6iYHVN2WrJNx
4kANZ0MLXLIdFFxE0ihZ7mNpUoJx0fAei78J3gOhk8VL4S8Z4HlySVPBF5JZAqwY
CELaPzxHux/tpV8CZcTSB+/u2amxbflucR6nYmxYuc8YLBcrdFxfFWnd636WtJJW
Vhh5B/HlXz04ddUMiUt3czkinBZugUhu0R7Yr6GwUEG0LoEHvvYJCr+dRuwisUnX
7Yem20rZGV0dDlv/NdEqMHZ78vs/xDukX+V+oMdvDmxApyGbTWTDKlQkbFcBuJ9T
Il9YjHRIqEDkb8UrWwtZSHuuL0+5ISN8MO8473bjYBaapcjL/goQkjPHPc0zC6Lk
tbLyZqjb/tY95Ocxgz7XNHNuD+bgydE++aTnU0sEITqX3ZCzzQiHjxawmCODooet
YUqpyC+lJJtjqKqbFLdCHfUQb6dPTVPdt1qlQyoK6JKH6Uns6EDbgNdGR3QGKol2
9KnZ/+SdQs4Swikpfm2zkqnisbjyHmRWXykx33UxudQFBib6Io/YKRXwXGEcc+cO
cMlOaSX5fQwwFDDKpukzn7QkYumbrUBnNsaUilnuUaysF1l1EZrxuW9hq8UXueIv
5oEIWOxvLJaZwFFT3nW/ry6Hy3cS43D+mrTyhvaNQJjsNTlfQL/0gJo3MTdexFx0
Xmm0EEKNDCgocFFmQxTnHslZFNYNKggAg0NAtMocTrAD+A1ZTphZj5aNf7olJCZc
U0a7SKKC9w44J5iuwAf61mQGt0Xg0Wc7eq+qFbdPdg0d/4G/v1QAzLn8dRl5itoL
33owrBRu7Pr1xbPRb3inazfdKEmnCfTszRx5za/UqAzhSYx0KB+HTcxfo0EIIXl3
8SeHzZzjDAvlnsVrAhmWVvOLlpNXhF2IcZWbu3yPurrP2KAaSwT/28+2ZvHeA29Q
FMJnKCPOvlMtMRPwhxHCCw1a/UAntecFfQJvrqmtWs4dWGnMl1isEcIjnJg2V0uO
il+R/lLQDzRRmjRhlySbel1ZgN+MQpf/5G2hLqTx23BANbMQ4QkEj/HFiuGQMq8v
HIW+GZuGlXLqPPVxSOdsy4Zymrv8l/TmmLhLxhN+msZ0ru75PiJ62xPJHIqUG8Ii
ptOVSoC9pRZqs44RJ4BytJD6PyRS6Yp3avA1kYMbBAEgwz2s0kEI0evLhtbaeqZQ
nKjfIg94ZXRnziXF/eOWAyZT4VViGAasyMJ3VLIRMbkBqrUST391TucvY5BiajaD
hEuHyanO9tN6wf/kXc68ArXRnB3pw3audSB//qqP3vRR/d86++lo/9I5f4O5iyjq
cs7G7wNsnxAHxdblBmaDCU/ADc12TinloiL3WCglAANqnj0Fppw1XdDovnVGj7hT
jko62xei7YRNvSdoeZhQPn+ICSLaypibhbgdsugDdR71lnGXgqGAQZlpmoXE7MfO
QTJLeykPXh8SSZRKKmdfaT9LHPPR403CTYZ8Ic2axqud3L5D/LHl9y4fO5w0b7KA
VajvE/VzY9wUIayfP3C/h05XIjKr0b2r1Kv2EGFxxuY1yo4fdlephnAu2dORXRrh
vyLvGvE4ymfnEmAEqZYAUkI1jkpbSyd8c3Xmn7RhVrxKaEFu/OHBnltvb1M9ehSN
T823pTLooPjRD8z2w42txGgrfVIoL21JQNREbdPfO1gOE2FcvzGqroUzPPpfL0Oc
fdhAQb8GvI7XErvDzX5LwO4PwyP4x7HGclItO0QPTi7jRbAlhxvLoCFYu+c+Kqz+
5R35Uy4xEBzd67IXiboxaYuoHeHSwTgearPN9XfVmc6UXaSsF2nxxllizzUsXJ8w
XjZyX7KqOOCy0rrwWEV0FMWyYMI5TEBMKej9khAx7BZ3HDetrNYEJWrBTP3OKKAJ
OHCexfiAWqD5lPjcAlu4aE4xra5QFSVp3jW8EhOo5PdiCSrDpQJ7GdK/172LgVMu
wtWb6Ag8I+oeyAOoWF11kKcZEpgM0mAadL7+LWEG1xwi5D/1go/Fy0c0txM1u6Zo
afxWZVIfhntaQNfUQy5+GoqXlsC4zhtC9T3U/JmqS2GtjuNcHse6rxXDwh2RJWEN
5R3GXf0d1D6gRrkYsUj2CegF77lk2rajxxr4oK8qwWlEt6gUbbPdu3HGOFSod72g
IMw/QMSa4O3o2vsTBSyK21wGbiIimS5mED28kmtNdRJFb3OhrnCdAFMPkNhov7Mb
MX1ljFikIbfymIi9aRn9CY9jtEXbDd2tYOxGYs7taMKeSafZ3FP1XKVBNKurpx9Y
/SJGURwLLMk4nPwOpRJyC56ODEH9mJe/p+XyXs0/fgrGeh88L9isLGhCdVfF7VqS
y3yYJvxX25A7+GKYVNl7P/YsdWqH/G3w61jK1kJbV9IKotOusOTlqdn6HO1lznP1
J6m6dHSbai3Bf6KzDELOpNUacHG21d7+gX5XVcYdAgkKqmtNqSz1fTuVUyfuAt8Y
0iKqEHriCCefoaIjbhMLlpHkgBbxQdWy82jxVEuCzs3HlAw8arrvguyE6X1jVvpX
k79WzdrHtXZdI6uRP4/giUmOMGyY2uVIKaVz5566nQCaSacqcMxAgTa2+R2zALtD
czEt12IQHSYpGbob4yV7D/0gRT11bYhNOjy7gutrHm8ZM/WTcEzdiyF1oWBJUOz5
IpwYlgd8vdeeuEekP+46dpJNBinXXeGXSuOGrVudKcsNZ+UWdzoHlf5KmjuHg66D
gHVNBOJpO8QX0DO42apayvU+6iOeyEx/UlxfofJ0MAlSQuNeHqNYO7l82x9pPymq
oA3mjcI1jxWX1Lc4kV3qYCde9vB6OLv90QHwbGOuNzD7TSRJvrV4fxXfZTku3TXE
tXHN0tWCyApZxs6KzXGJUpy746B9Sx3v3HGFjTRIvCGvN+l36Qtijf19IB5wV1vU
ck/sG7082b5ahao0eDmmKtCTPWBxDDI3PAGJRcLZEd06Tvlc6GWlGvMcwC/Nm3Lo
coygv9/5hcBCxs22jyT7HNUkDSQq0Qhlxp7UA8d+kmh01ZXLu/35C9GDWb8x5npZ
BfMrtjNMeNgOXiLGoUOoulsy6Ci3ZyKHvGV6lrEaTTHrulDI8TK5/Uc9oXTHrLfO
9VC36HtyLhd9VF3soo9QzjexsknZullwjPIRXY9uIUIYX17JmQVTV3jS5S26Rimp
0aztAOs4eNVWViPj1Hm/NAWkZbyrPlRy3wMMNj7UK691X3t9bXWQLM5Ttr5JJ+E6
wcfyACW40htFHNmxHFS0ypPPz0uglp/YgrP6b6IRkbA9qPFI1xpxPnYELIM90wxI
k7d/+G6q+DGq0iq/mvM/OujFUW6ySfLmfWd3/Y7yb8V+zcIVMU9E/1CdTlsqenLs
O3C9bvsxRFvJl2wp0POb2BpZpy+f4Go3FxN32X+XncRM7m6XfLCJ7C/DtJwuyoni
iJ+kEnOkK+zYpheWww7bAt2N51GKuf20342UY5SdZZoYCuC6RilBq0i0BrVQ4ASg
sbCHvhZGhKSioCNLX9QvXMlaBFQaQPvKpdFVFPJKJ5ObruMl0EY+tMjjwLN++fIp
5hiCl6+eS/0RXRbbH6qZfkbgXIxqFryn9N8/TjYbDZtETa4p3KIopJqkU6Sh9J9w
oIOpmzgiBJHagpbdlv20266TDfq+3Ln4Z0cGXbNvEPE08S0/DsVpxkJ8tznW+fj1
d3iqtF/H9ibrsvCso2C35HUXafr8nQQwLtBlPNd47bP+ib8JZoCvAJSmi0R4J/ZA
1XywJscljO8SOdgrNmNmVu96R5v8S+DjvJOH8UiuRmvQzHCC8YmqJSDt4nb/YGWZ
DJGXvKZb47zLDH3CR2V6fzWXyRQAfXmuGHcf5FxJy6nMYIUBBI0DJGkC684CsjFg
oAP1DLY84xRTaAiILkQwL++C1zgsgG1ftdHPp363EGpnSfYzCtTw9QLWRQ1gRLFh
ZvAcTIZYFzBmvLSE/z8eATrxYmBu2i5sA3GvDTPMdBxihjgrqRBbeZYjXMTEAlfe
C/IDA1L/XQ+VozL+3aNWJQJoUwrw1VfALJv0bNaoy1dKLTRIrJ2ErSYIi59PrLsR
Gbwz3LIXrjohAJTWneDhNWCMMvepDNq2OJSdyXd9VHmXIlHtysflfA8o4fLaPXGE
8b/O/vDESM5ubxIF3Osm/ptoY0kcD54twxMyKAVyp8hmdDHU40pp17Q37ukSLXkt
T28rF8CzXNOJg85v29ZB9Ebj12dpaMlpfw67i2LaBKUsFRuH59QyakQNOPhg/lYT
KvNyxKaLFo50C6rhoMkzykEZ6QzKVSlWXYimvbvDyJHYMXXqhTeIpFauHHlz9clO
Osn+qHrC3qIYD/7qoj7L5BkUA0z5a1V0HDopx6UlMKEuBPcXhg96FVQAp1LNDp1X
0dozUJBaNV3mUvsZxnIKlqH0WgcedEdMvQVarbFe/EO47+PfoZ4cMr/gc6ZJ8uGj
+SDj2z1BH4e2Zw+t+sv6XOoNT16qXc/k7uVdl8RD2U74ZQmyw2EwK3ddhGVxqmlz
v3cOqOGnb5EmBlvlDjfC40CEzKbNyfj1UTGhzFHoks9jirF2YrUIh//xbYfq6Fy3
jK0bMGptcFPRsg15MaCmT4gxqvNriM0BItTeQ9Ushw85wQeEqfnDnvBt1ZzGCkDp
3HTui2DxtYvLNeBPc4g+/T8xEkIZfdSecnat6keXJVv5zEYzcBsbowbiuDvnpqDH
qLQMCwWR4NTaComavS9sL/f1QouAeiT/C/54nODxHcYfmn/G+uEqSzFV2WzZTe7z
JoVEhP5FKnpr2sRtiDvPuIpYKlAJePmLXLkCf1mmEh0MeooOIKp3pIfzcyqcFPp3
V3rYN5wKWvi0WrxW5EBSduMzCpiwqT6GEx46YNemsyYIzpOJECpIOnLV3Foy68W9
QUmSLR2DGOsM8ocpeOpdc+DbXJItwWbdOpb9L+RKwZfjwBQvqMFbc4JEXD3FNnVj
39H9+BqVWAzKStuaHl/zf5p03aQ64N+0HhOfCrLrxJene8KMNWJykwWgCWNz/hfH
zY2QnXPeKVHYQM+NW+kBmnJiTU0UyB/uN2OT0f5bLfVy9WgOMxz7G4NEZ0OTf3Xo
E3CePBCyG4f9PFUbKTcqY3YT+opjJ1fWZ8gjpKq2SWk9hVuNs8ijoUpBOvLDVM43
3LCO1nhbD2GZwc618OfGVSLsaGfl8uhZI4TwHn/dWlr7Zug57xqiBXPlUvGDMOgf
l4tluJq5OqqFO6QWS3kLmR1nHSZ33D0eTebisdhLBCrPHyeMWc0UeewsHoJmGuJ/
pv068UwyYvDPAhAoVeO+ggmYuhR6YYr2KxVRjpUERWRx0LoSHIBLhi0YKl+q+HpN
ztXXi0E3ZuPIeLDtfjZ/KitlKC71iUUyY+Bq3uRPvnC5oYq5xwUUh6oDu4PoXOOn
xIE0onkYOUMrtmDbKPu8F8AqCTi20P/ytVgBVKwgxtaCDWGUl0DHVUIAn38j/8kS
o3xoHs9ohSb0i6nQri1leJywJ3l15M8OusjNwsRonAbzclFQVmkiLGGBLOsa1fU3
t++GutI1ktDL3kj8DtwMHcQs3JXjWaURh0W7mSi4qqQFg7LBakXB4qmyzmN3ZHGw
/b9Ivvl5kNp//ssm2g8VjXqjHhjP7bjncWDcZ+8/x44kgTo0zjKImQXtrwqrgsFQ
P08lmwGzQ4oJ28GsSuRINLsPLbITdnApgbimp4KZ5OjsO0sF8ofNHY8comfYIsKE
h66ojDlrKY8Y/uHHwmCppO/cPWBCSp4J7xciP/SUuzuazFl6BkPv0o1fCWbKicBI
bkD8zkEI7gaxh4hp10plXFBaXXiWgrfkUqBWslEL2G/ehfr9UMNBatgLiJut4Mr5
Lsv8KAiLzdJEdvmiXO1vStMkSLZyOyYplTn25E+ZCvIL3w967m0YEnv7JkZUxIHh
PxkXUsIp/Cb/nSQDpRRjvhZVKzoTMrrfQhKqwE2K+DJj2Chlky8eFm10YMI7bhWl
TsDY9io1minj0H/TPmzM/HnZnUuIj8yg22W7Zk8ct0HwYrQNhnrbkp2swwBsOIQ+
Ewziai8s5PtkRvDFQ76ECGvzbUBFOYZIInaft8FpSG9F5Ieirwbb6zAyrMsv55we
eaMjgQVOUe6wgRUu/arK814Gw/v1fmjIBvE8qam7HqbNYYvj1rc0dBBchw7Z0gmh
REstWbDHsGerqASW7ISXpvFudIb0YnWtCToOWTjTfz6mXD3sqHrK1Rog47xwOshd
L0FqxCNxIdAV65CoW0FnteR34ccYhDswsNVPsycuD4d7wEVe5dVjVQ3OI2/KY9Ax
65j7KKLSLr7MyHr4LNjWUYRHosxRbv351dzgbhyOtxCDn1TtVQU9X6M1q3gwlq5H
4SkOYXhBSn94avgNVn28fI8GqTtZjqfr/iumf57H8tRqdWAIvOhlU1cpOFY5+Z1B
0U9czJlg8vy2E2gA4JqYSeOpOr+qVtK1NNsz3RyxV9C/PJC4hgYhie+QeICEt6O3
inz/TNI23q2QuS01eO0xD5gSEJbwHe2I+8iMhdlZI1oSAiw7dsyH7JJWMIn4rn0C
5+qUy7iH5un3RUl/MwiWx6hft084PwS9mFgpTXuLjd3E7rD4PeJh2/5HATYZ6ct8
fUw3qaRuwqtgMlx9S3sq6O1c4D41tWZaZVwi0w5pbKqj/F2yG1ldzVm0bzd1frcd
6HAWziU389GpKoQowJCs2kZnJdkOoQ03RGEJLpiYwf9b9lYKPbm5l2Z18ZSqphMp
DjO4Jp8XU+NrsdsC5Z1uUsDbZZRYjzelTYe8T50ctJIVNA/XzbSiZwuPqGIlYAds
SrJ1co5r1w8SrRZxGQqZunLeAZB6wAeniy/clW0mDCIeol5zx6dwzmYk+TXuLCIr
SE2mSesVzVmB+k4iniNpc+nJiVGRnHYiMg3Fkr2tS/tTqZW+0DuhTXJUaGHyz1J8
wAroH+YNKcFD764KPo0w5THFsXjZbx0oXdcgc4MnR4u/vSO7pewBrGk2b9GXpEo7
hzM2QNAJv9pXCgihaglyTIsHoDJdX8C1BcMPMbKbC8iflSEsC6D16tIfxNx2K9Uc
ajdmsa5QJPnQN6+gBkyiIk96WUUN8A8Vz7aytBAVuxdIIOPpNgAuhddzIOynqNJt
FB4NWY/Jc+Y22mFgIvHTjFZoeA5vKuR2ljU8yXmvZN4xbi64txqNcA+FQ8IYiEnf
7kZvpAK+qCXQoLUu6P1p6vqirDsboxfONXS0832+1/Da3U9P3HVHECnAX+b35Sla
d9reGuCNSxYXvVJn4D6a/56PLG16GH/nYWJ/V7cOv0C7HVcTiJBiISETGOKM4z8s
W35Smf+WyGskB+gcVaT6iXU4TyYEWoPAndWdIW7UujbplqgV66UwZbCPlK95F/1c
2PanqAVQ2EVkDPxwR7F2wZ5UdzZoBDgmDuWReXqsHJFRqL84Lgjg65YQ5E3cbpGz
q5LFOTCPov/W9XXz3rZOFoc5ms/E4Y9TnQEtOHwqSyFFc9lmjtqfMwpMlme3hpxU
pAtPUeLL6eM5KotHNTo3xrAh7GbZfUlxoZRrSgiMBlR7l4uQSsI1jq8a9CVUOrM7
9h5wPI9gjPG/4MQSR1ZuWT3nFWD28ywIBh+gW3n4Yeo0pGqk6QwE6Lb5ct8preEN
pbXkvZ82NMtCNcJ4V39809R6UxJDM8wNQDl6xHtqx4d+lFbPJBMk1xK7332cwPa+
QS+wYqKu8GAY3Pd/+G+v98sNZeyU0Zt6hYHy/biTNjo3K5USyJRxfmqeI04H7oSY
e0Z8BCEjFoMTIFAIfeoS61xGDvWEtL+Y3IgAF5vWt2+KypxaEwguPug5DUiJbQn0
jlPkW3sEqUCMGwZp5IURncYYSu8VgRBG2EpjlaUn7Vg6iLQu+wlMxz4afx/rBTfB
UbisAlhxeY8CgyouGaQ0b5qpwqGgoK8PeDGQDV4rYCe476MhyES7tfNUErPAiEKk
fBPXKvyjgE3hTZn5kc3FaibhQSYJP6juRpyaJUvugYnAsPDrSoJz6KyeKheWokTV
kwBmR0EWGbf3w9iL1iesXjPuzPQ+dkDgW0ggXp0zAXxDSxUngHTliddLEEh5E9J9
m+gY/yxhqpupsxdrmV/oIiWFZ3GM53KAw3ikRTe+KSTa6d9fGEkNdJslWH7DEbYk
XyaEbzFe1qR+ZJWvh7BSW2O33yjhOuZQCUVaALOBw7kMiXA5CwQP60XJIJiSYq4r
DERNSVNJqvr8vTFaf2SsgT3d/8Pn3cNu1DYkL7unOBytRn8acFbFkuldmDKqqZVA
6h5xP2Anhi2vMw2/NQLCDJBsS8YZK6pMBPgX2D36KRCcu3v0qg24rxYgf/8qCsLC
hDeax3c/EL5FIkYrRDCBPKQsmSj4z/dYDeW/Dzx+mE0jDxa2ryUEU1+HPIOg9g1D
W4A4xwq2WjlzvkFltrJJrdMYgB0hJ8guknn1miLTE/noKVkD6wYreILnfzjWeNEb
wp4Kr5Qo0tfUuL3mtjg7LPUJ0k8b3dj6L4mSnjJlq9r3UgD50HJr0rVFFp3hYxi3
eW8nmMxzilrWLNKe5tm5jIMTLKkcvIE2SnRDmQ4B7lHafomB9HtK5b+wOB8JUpWm
D3gIEfHZQlbnzLo0q7hAplw2to+aYMEaXXvZwoiDtvPABQUqiv5AEYusJmlBuZdn
jQWr8GeM8IMv+k0+gLlTW+LRBanig96Tw21h5IFyeHYOxeAGJAS+zUFXb88YtBR2
4GeEaIMS4ODmV+IoWAj+s+fQX59/cFLThwAaQUKteEfF3ScPLQI1EsKDKFZwggZY
WZZWXwArpeXQXtsPI1G92ywDxzJ+upWb6uCIvrFmTupod4v0H+xoZEbBYkKaIdyu
R1yXn27EHolAxLCKzYDoUGFLdtxiWx9cvBkJXQYh2WHUCWftZW+WIO1Vl4664ztJ
esak0uhTEwvnEYR4mW6vM9RrYgm9/dcLDailj4UVAxgbgmfeZFPBnDkpU+V28sHX
2zjery5maOHQ/dYs7Q+pc8rhHGsnvmiRgVMaimYyxQNXa4lYwSmEmsza+qjAQFuQ
Cax0VPWLX0alvo7kzw4mK34Ub5dp0ztswblu8dX8cz2QnOlZy6aNrJUCW+Kep6pi
kNaF4hnpI56ExsnqaiqI2EWjN874wT9DM4I/5ZkoLZHMt4DpAF0q5LsjrKYSlmIu
yinWJwHWAEknMC/jEv3N26oP75demKkAuSW06s+oK+TXv5kDD+VPlPbkCknpuA0b
L8r4G9DNxJWH8Ifg/hqizhA19gjX7ETLvRefDkLOIzJTPJA6KvzvXHh6opnyLSpa
rWZCTLVNwLzUB8tJnszmprVutAt813s7MO9GoH8JQ+Wnh/6+NixV8thv+zC2h/UH
PD/dcGaKnuIcOGwsdWfxRwJevHxJAN2MbBpR2Q6bAVOl26wVEzkC6GeNJcWak93v
eNuoDaPjrjwfLpV8J0Yrkjj3HbecGgBff+1Iqxp/Gzhcn4lMxUexM5vEWhk48qcA
n9fsrQD2QKisGYr2w0s7ORDQKatAVppUvOPkCAZEckHr39bOsQILKCwjzyQz/eFr
iL3K2IrKadpFBx+E5J8V019gzFGHwuVUsoeKUxqzqh52b4RELLW+50jRb5LX3kSz
rxZX/dr6jrFhHwhtEcn1wWi43nbSnNwEFjqgVeTYWW3W/cwQji6DCWuNdKmdDjVV
kmeRVzKVX+ECGngRxTVTZt8rwgByBQKo1xhNn2tiTtG8ZMLwXdIF0xROMP9GbamK
lEKRasJrgTLsJlKiEYsNW0nuMfji8AphCXTP4yHj9QYVRY766rm7h+uYWI/cGICo
q7lo9ZRQTwvxichOzFxS+ZLJInbMb/DJu79aiHBP5VNpVJfzJm3UhuRyWDUt+fBT
VvWk901whgg9tHLjnt+SmV85SWNhnSSt5OKUbaYMkNQE+41gXjA4KzAT9x1Be/S5
n934rIJmKF3rG5PUSf6vrb0nChTOjy3QmOq20uXo8L0HWs3Hj8Ff2UlyJWBJmeoe
xKOxLJLrMP7PRDq4b7ohvG+IIncAH4t4wzlUKutCMtWZfcgYSJy9trWg+bvQskeY
JousBcRt4twEpLEjSL9PHS0vDoRz4GTgjS8iCCvp4A3q3TZFeaKYqcWAqV8y9kXB
gV3h/JVpJSfDTYSkEnrQ4bBvcp4zB0muZghUZuUrjG1noQgW+ejOf0twyJ9yvcsj
pOME+vt8kp455DV/Tjm1EPxFChJd7ekC0pVa8A6f4lBgsDGtbWzS6q1K9UhwBQf3
rzkBqNE5eeSrSwrZKIUYOr+NUuLec6XROcOW5RvaPUsRscc5j7zFPn9p/fiJ6RNS
K0UqQeo8sO8bxTe/2KJvDeoQqqIConpZ50MaRSClXSlXTUH0Ofam0eH3HFA+F3dU
bdtamDinKc+ELDBfRKB2sr9yufNr//OF8wo72pfniQOrhyhHn2lzum4PfZaug8v/
rw5D20r4F6pCEerwzQyb0jS6Zhx6huSHMwL9/F4Wu6TaaT8+OWw69SqwET+uewM0
CICrgCxTWPcEqtm0S5tqkFZ6Maysrid20i3VjPnQmC+XpmZyAGKI3jrAOFyKD4OE
9gooI9r8KjlBUVsSt1PHmZ/rDgRnJo/AkAUWXUpEgvKUXrzDtrmUACC4CjxH8DMo
nSAvv55JYbcWv7Q3DqJo8Rkkv2wHNnnYcLDDJVgOTvdYth4uoFwD7QTd6jaQ+N1L
lXNr8TKjc5XmyOqPvdxc7T/u9J/p8qC3HIdYdj0Tw19VG7aQpiNCa3CPUyq14OWm
XBt1FMYurUkqqonaBOgVkRyDKBhW+zs83lHyFwhEVR3AeKSwi6utuzV2KbpkzJLK
7RUewdP9+CmnQDJkEqSBqq/fLDxY4cIW/zVqBIvhRGHNW5tM8ZXpR2S5bEo04us2
hqbxNV5cZe2OPwscKe0QN0LmwRtKqWa3iZ/E2jR2cApfR7ILmH2u9HoG2c/Uuers
JmDG4topUURjMVlT+v7D3JK0D7p2OjtOAnaLNCz6qaj3bY4a6YWgOlv+Co/kYJCR
yrhbbFqE3AnF0arFoWC/+pZ4C4tu4qjUofbb4Ov6wdJdzRL7mTKtZzIrG8jxBFeA
fWY4r9bqq6kIz50YwIdkqw6/aandtOv6+TTyWVAqROr43npVUDzq8WoDSSM3Ptb5
cwLZdltXtcY0088dGGA1oR6oD8sTe6i7QxRWTv1zvAMZMiR9MOwDG8wj3ng/yqV8
OQqa0/eJL+J2T1ysrFE00P6EN4JZ1XO7CkKMiH6xvmF6i3/VKc2GRRbbFqY4sX4s
QBTJ262MaVgtjqMHmzYo738pXAvMYvSHGlWFRTM8xp/3cuFXGS0vaeWzPOPTGSNT
zHMAJsSrZyKX89b/nkLmqEMU50nVjxicKLb0yWgAcXwI/3dcIG0xmnpheYJAPOtR
y5tvdQLJuxcM2bqDdtq/Hz8d4a3JOzH/Biyn2VFIK0lcE6TFKBb8BtLGjOPc0hRR
EPFNCcZFeZa5UNV3TT72XvWyw6Wq2gBcIyipUexqf/AY6VYXgcpmgGcwvv+HbkXU
YutuigJyV2cd58WpZcvO6IoadYcvCVv1g3FhYA5gRhu0a1l6hvqVYi8lbJPN50NV
iJW9gP0KfrQfwho/9amc5TCS3rnL1hayEv2ElOOsWvFRIpubFhrV1cbaakB1GiOY
7sPFqdVcTe7h2Qf+XfNImiANcJAV4haruN1xeOrmFUugSdv7jyZyzGKUru31fN6S
EWWPVzt2DXdFyZiXaJZNReZEHSshXP3ahzx8ZaK6U1X+9VM11xdwbq2gddPt4Y0M
US11b058P2nANP/jrkZk6ZSn2P9T82P0lYB5FMrFsU2Vpn7ADmGFCTJgXz9dslwF
3S1yNf026QiRYHLhbTe6i3Rr6rX7w9l9F7wSDLwOsHMeN9O4y3wdnPhmnStl9aeq
Ci+uFpKuOBsZjYp7zZB7elu+/tRUudeLaEaQJCnRije3+K9E1pgBS3cps1Sy3z18
ELLYMhOcEcD7hjkWUPsosZIrH1Qkq427yz/7lGtEA6GBcdVbTAsJqI9CPdZX2vH9
lTLMLHvQ8JEb8zv/wJi+fYNn2M638hBnxCIZHLgUPt2c9kjtivDddGl/Z/14Y4Wq
QBoUpPMgTEvsd+y7sD8I2Y+3juakgBMUS26Pz5M0o6xfBqoEKNw8Ze6x736DJT5M
Gm89TXDAx0aGwU1Hj9pv5ePVTpJbGd25bdjG0Pkoj4xORmSqDXzEkfshumCuk4Sz
y1XMrXSb78SJyHIYxAwBwlPQ7p7lewaLf5A27UsxVXh7qG4J7f+TQudgk25jI7C9
op1PaFUdHKeUDdKLyc6dVu1RcVBGTDFRNlfmCDgJq3sEj1oe5EYEhCuWJEJ6IZS2
/PipR3G7mokl7OpythfsSgXE5G70fyGsEC8WP6TRS5XUZRprhogMDJA7CQwfqvCw
lUPVYOWLjG/BgAYeexKdzWOVKRmIX3u05Pmd4SzTwNjYf8xe8X4E3lagcCN1my49
UQn0gwfEikXpbwsG1yRDfDx17c/MRqArAnCVNOht2ms6dWKk87JYMrJJtftUiLap
9U/Pc8q84ji+bvd5aWdpvrITxpJ2yb2nb0JNnsmFCY7uao5wzQ5xHjPxVsFP7pSj
SEwE9hWZpA6l9Wu1Ekcsku7uwUbzVE/j8dTDN8I/3qjQn0h9xNQkKDXbpSRExoYq
PJuvqWedaPh2jgvvf+v0dFTONGGZ0cZjIRi1Fh9b26nOjfBDzBsbkkuNpbwQta4C
OmwY8e4pf96OfyRp4HhMryAhV2yl8H7lArwdccnQhoOdbZERH6DQNXV7wQY5A9Qs
PAfko62gcQlXNMnvWpi+Uise+j8Q+pM65/i7IE9cVrO+cE/Ux6ZbjhDsRAWHI+oO
SWpCBFa/tLFUJKxxZpAkmzqtbZyN2Roh6vrnwnaXujkjKyPz6wGNWNPmpoK0QknD
ALbInqtX06iujf9jgV9ctaqte0WW4XQ2Xs0rzdEb76WmupAEV+v27ovbym05il5X
np1oPcDvgTzLPU6STESSAH0glt64ax09MpUjYRgLlase/pbP13B5GxD2xX8ddxoj
4plZetiQkpn8aJGJw1mkQBfFswijivLC8DZKBn29TdBdVRkjW7v4fnRdDu95voXz
fAc+Fccmb5l2y7aJwjfVG1WYufrkX4vaJ7cpUEzHkeKYACP6M3WtS9tcSxBctc1/
L2Wg2IFqlinpH0Lx8hVYqNnluyZTsXLZKkWDzDYxjB90X1SVrmE5bNz5kpoZVfAS
I13+1HuZZ1Yhadv8cnTUwJEe8P06f9SNpFuhs5kAlznsmIYvku2sf64CjlAwoq6y
ffa8yI+9mnOq9VlwVuyUBbc7xM+yCmt7LajzDV4KOlxJCJIVRzgEvrjpQQ4Or2/+
0zqEjhKqVHoU3oy/O05CNFBhrPngA8y8dsmMM7VwW+1YiwmyuxEEIN2MIKxaikIM
N/KO05pIlHifzuaV2clwu7ChtRgTg4VG85H0p65O+FL+uYXBX4mU3Sc7AJ8p5VXi
jwCFyQ2REoX+GHZO0Ba2LB+CLDBRlAFeJSqCeLeDPVH1Q8q273LYBQKx1h3LalLf
tEFsHQ4OzxMOKo2lpidCieyCGFGm+niLkx9R1A01e+JIdwGtlfFbUiC4T6FfQyCe
ydc+1FdvdGlHuUndms/DI6/Z3fRA66Y4vcUVp30YGLWh3d+PxLhJtGlPCcuIsVer
Br9FkI57E/Mrkv+o25smjJF43nhLA3mLtS6vOiXpY03Qzyb47ygaSm4NbJbdN4ZZ
KB5Xrp3uIm0csl++OavjFh1cGJq3hobI7QjYod9bPXJAJ7FUtuG7FhUvFFkJadOP
2MyXRLhJor7HnUDJfX4dVSUg86q7/mVK5N/onpY0bAGxcorBzQIsvRE9rbdFPR+m
jNoZ6iuyuWLkkJtMwmkcOAnYV6gYk0V7zjnrV3uu9G8hSyeo+sPOtWMUsxKFCN5g
SfuocY63v2HXCBS0dPF9URArYWDk4AI2+bF19CCskBv+rLbi7DWtrvOnl7DyctiD
xZ1VIlqxaT74r7nBXdlUj2PtZLJrRWWf1wOY+zXezkJUdB27q2KzyimVEPgr8Ki7
Hpjoo4AuvUf2Soix3PkEZSbSiOZGSnZvJzd25o3V4kyuc4Rczt8PDSI2dFLnTgO3
aIiEGgafDalvnvyXT+x96P1HlIoleIeRfK25TusDAj0gD8gmtklfyUgiBzTbHV6E
Pz3Z5OOHBW5yduE6Eo+4VoPqN7cPJsApRL94KbNnRwYv+Dq7vJ36mIUiPPe/bIOz
i9J8QT+bGH6XGzYpXkVE+j0kRZtPcKh93tYA6zVzNW7psIm/V7DZVedlnQmkbLIf
ghSerIpiTtutjpqFkb048gVwZU5X8XgvslQFLutlT/0ggq/aaQL0DDPyoFGXsrEI
EixP0K7QvrcvGtgNavSU5Emtp3+N1SlVRs77a/6gZmICGMTS/Sy59gCqCNIhWkGm
qcnkmymsnSXdYzf4HTRanmMhsu5T4ZkLKEBwy5bC39AFHVMU7gpugwSbM6xWAH0x
fgaVojuljSMMp5q30cbMIaw3nCeGxoBI+2vaoB0Ux3ZqHywNgponwmojZiiQJWCg
bWJz51cnmvhjX1QEjwvDLGDLJ+IxW575DcTMBcSMPeaKiQFuuENpjD2FAEAxlrqC
eAx7EEsoeoqKMuLSGi2Yj0u+zEc6nndvgzFxpB4KOZ2Wg/Uf0IKhsUSHEkT4bzou
SWPerjsNxP/jTnno2gOY8nE/5OqKdgMbbpp05P2uFMXghrdDoKl+vbwyGor6W0am
NepQNdsWlqNR0G3eVBLjSUASv2I1zivYEr7gpdHSvFP15ex908ZdIronJWe2BUj2
XErgScm4HNQmiHagF3Rn9ZNbILML0HVqfGr1118U3l9/HjVn5rE6H/ML48rejnZ5
0b4jYqGk5wKgMJr9FCDmT4yDJi6dpgWW60DCf2uG9J/ve9W2rDIsga4lnJDdSTIK
vsUEqRAQFLWsmQRPREXfxM02dEtR/W2pHtvszSfM2ZCEFZGPOq16+RCgxKyHoQ6K
0lfco+gzwD5mLSedsV8nTOxNwX00Du4qY9yII7GUtkW/8Z50K8AQLMn0SoijEPZX
mlNZ1752TFTIVfiutAT2ZpSP8pZRjcWKBLZDAW1bB16VqtNth7Bu3iRmXLzBdTKl
0s+6FLxFpc1dcTogwa1oOTTjcftLofCzrilN7aWcLTcjb3L+wbMla10/AD6fR3O/
2zMApGuuneRpw47gHbGmzcRQGECS4GYTdy4h2B7VbLeiXekPjMSsrS7vbIxQNoZ5
Ts4UKXTmEJWWA3tZcAeB8bhlUA7D+7PRnCUMp2jwYuEtgMquHkuHi4r9Nr90eDvh
ytcJD1vHhXIJTz+OIeL00DhftrbFkcr9q/GaqwQE4Rfrz6FlP9wNxfiE0r5MpWEH
8I7kAu4vEzHMtMI57rSZg73kveLuSLY6p77tHn/48KS9bI57q9bId0h8+HV7WZCV
M14TN6o79vwC0xwjOcsxkPjDtg617P+PFJ4phUWki4mnZLeO9Qp71BDDclBjS3m+
HaVzlF1Ia7Q5oac7w/A4B2i9wSGkJdCvrzvQk3hWikQI4IuTsOVIwSwr/TQeiNjm
p07dKD5dWhg7fNSbRqa8qNPnH6/Kh9kLqQ17V7sZx24jeBAZAQLc5VQ+buAC7KB+
jq+3TYRKHSkunSVAGdZ/MAXA56eflADH8a89iZWHKIGJBUVOA5y7be9DuywNbOmA
TtQHH0adu8BRm+6t6WNp2hhX6Z1D9Q40uiWPfKbltG0Phvdsrg6Bcwjgggjrdy0T
E9eIHvdo7Y+8ApaYjyZrYZ35ev2732CYZOGn8f8tCQCCXaez/WrKicX4mRUpbERk
Rm7EHPme87HH5u/a3o2v4xx85xcVaRwrQVIKiLwpRFu8yaR+HOSosBi2peWBqa0S
TdWT0o1U2orYicjSa9PVPlDCIOdl60Xb5YjHxCQi++YFQOWLvdl1xVqfB00pR/md
icvJ8DSbkB4NRutmoZUzaGtNlY02QYSt9TH2hfRQjVu6iuj27/zDl0heYPi4jxJ5
iq6bYj1rt0FIY98TDbU3fidk7YrglWPKe/w7MRAkFnXUsBPVR0YvCzdThkgNKL4o
RlIuaDrNivinU7jfjBvvdRhDXrzu1EB+WlGSdItcxXsx+QOKRiOFaC7Klg9ZoW8r
ry1wpEx3zrsHB9v4S4bZ2WkI1GTfsFbpUyDUH8KVa1tKg/KBiXe4Igl+8VBZfP2W
dgWLwSGGCaU9i8rPxN9yKnGTyMfWLxJUP3y+ruhzTe3ym+td6y4VFRYJWfqT9Xti
Pka9oRlqgjbdwm3PHrmEiUGjy19jbuO6Efm7WjTFW/FePK9aGYZU7+OfPvRwpyJ8
qDSIDzPMWQ5WWnpbaXkSQ64jIdN9/n8ClRWQCA/IcEKOf15J/RbTTG/S95gMBAYR
F91eXokhZqlUaFiRnk85iXRl9yVnVZkZY7S98YLW4V36A3/Q8Sp6ObmPpnNCWkga
bABxED5r4da564TInUhgzY1KCM65Q4PnSzPah1meefKprKR7uRoBi1Zb2uKl5ZEg
hx+spTVYCA8PDsFfOmbOBOYpNWQb9aBl1cTBWRfk8/ZrGGVVJIk20krrh6t+8rE7
fn11adFh8ocwOBsuSLYWrUWn+cqFmlGSYnoa3V/Bqsw9JWXeyT/V+dWFkNogcANB
TSnX0mGkA+mmvHLO9ld4EUl3EMbwWxGbrN0ovvE4oiY5jo2WdM8y93wTD8qJcqLq
lXFMc12sNTELg4urv9rsY3iKpTXrPRCLS7ErbS0KSUhSmIeikgVq/hpi6if+Jylk
otDclfpzwGrs6bX6pqFfpKQLlppqs7SXrJlC6kyDkN4jArh4qflUty4ddajMYIyx
jlu5SMefPfVaT0OGVo9zSK7vxY1yI71QmfliqF0R1PhZJFkRNzd/4hnu785K2mZ4
iiijb/jxi+j3h0x3eqDo0w7/OmJg8+epkmpd2W0+CQ7qTDrYRoz06eA3X/3KeIXP
uoAV4fXMTwr2Mj5IptxA9Aow1tG2AWfhTAcPrNsmKT67v29bSOcf8JJe566eu58l
xUFK90s/xcxcmoHhIMyLciP0tKBvI/4MSmwQ4D56JUvUvCjAU2sI3GEVQsRDECc/
LGxxBOycl1hjt5N51nZ21PT+d8BQCUH9u8DwNArL/Bu9fdTQwXAv8rrG1DFD1C4g
zNtLbdewMq6pL786cMSUM7/psSWH2K0ePIT/SAoBZm+N0T1nzN8v88vhyHtauPqE
ujnysE4uJJV3Fp1MCLRBi92FbbVNXxCYvocK6RwZJK/ni1whDpOq+J7MzUrzNkRQ
ivnZeiF4x1olV3oezTSrLKtSwOW932Nni45EdpTkeXJI/MraXDhed+20TG7LdWue
zPRN2ki8X/rU+M0O6RpLbUFae/6CHu1soOuMUWlgnxZOPFluF96E7uiyTa34jsvS
zE3lFDKw98mRmglaN9LJJ1m7cyNbZGOTMU6k7tlWD/zwCplcrJ36LPodlDjfXEhE
F/OV/dGPVwvKnqzvBnH47NmqG0iNROweZS9MFL9ldKiaRP2vxv8OFYkaC0R0r9/c
gZkZ3Xw0KeONJ35+LZpHmHLhknGGolNH3ne6zPH0KYklOH/J/BGSvBzOvsvfepqP
TSAV52Www7NwLaLUd61ETDBv61eipHslMOmiNgD0v27QXkSaRv2rPvz1X8bxIO2X
NDXbsQUnXorqgm2jKVu9KcjFhc+5Vj6LF+e+E5858iuoz3fv9q7oJr97ZrAHXGDy
MmpmA+oOpTN17tba4/7p1dOPDlC+NN0RTVVX20hTSMQphhZsN2who5WpAlhY4IC4
bh9YJsHmLvJV+D/p+UIMtni4qKvkeMIPU9dG/aEbBx4ELOLVPXLbA0xgIlE9tpvE
72v6fCgK9Yo595iRBxB+EL5JRUTBR3pWeN1wYTaz5Dd8AEzOopo0YiOkH/5wZPeH
E9W2rUj6yFBaQS6cPFFs536d+6a6TB3sjWiVXoj6Gfe7/uuvm3JmfuIbcOS/sOiw
JozXYU+iF0dOlRkdEko/5rFwSLLBBZaS1+P519/nMnMH/01qMqU3Ovdbs9qhQ9XR
9JT82XuftYIhq0UVF3deN+VPwPR+K8S4fH6EFR3iLDPQ05YFvcxr9Z7Iti1kGZCo
Q4yfVc2qXezbevicx8qtHPwBcb+ycL6HskRXJVQJU4WnYJ8pXkf/pivEGI75GUs4
Z4PU73VwJkIkILVCcuC6hpK1QYj2FsJGoi3EZEPUDP/Ta44RAJ81EB1f7I8Ndtr3
vZKRd8GJqzOJNDAmSYkPEu2+r305EGP+CAO48mSD5qMKpWlEoE3jL7LFTS9UxfVg
67wA5Sh3+nL0ZJuysZnlVDWHeawVQHYq9jsloiUNx4j+O4AgMwHTZrrZGlw5vmrw
1WJHsWiphJhFj0yAettE6EBgt7Rz0TBS8mcZtpN2PWE5u0dt1fCJJKzimSIhZks7
n+0M0qzwCVZsibckC2goH/CyZ2tdsm9w3o3J7DZNJmRzDWJ3PBrkANKEku/WIZ7C
J8wnTsbxDSygNB/Ocq+6G+GYVuiMTDMFCWTfD7m7QTp1JW6cNXOxf8Ikk2SsI/1F
XE4oPruIRNK1IgA+K7IqSyRNYsi6Oq3Qy62s8Aleh5LQOazgOvf8GXDTFqICzR/H
paFMqMG8myZbqEgH+me/DHL828stiyzFe3Lhu+XpsuKBo+Az4U831UPC0zwvH75c
tG/nz2kYiUXwA7RhaITLJi6Y3uWv1Klyu0E2R2CzXjsUHPUOO7f5/CLgTTeIaKrb
mS+0bCi5Bxgz9RbTe4HaNGkFpLf0B6i39nublfCBmJxQLqkHO3Kads9L502BZP36
WZ2Cw05P90w1G18rgaz7FK3OzcaeaFa4CKZZDA4Z2PUkQovaGkxADsyyQQFrbftf
qiAintuIsp9nP2Srz0FtrrhM2BMOs0ZB6LHzus/wNt+DL2fI4O+lCenA4RbAUX1X
MHzr01m+BiwI5C21ih93SgmCglpdrEe8TlNGM5qxE0C4jlkDdaZl/dPfmtEwcL1Q
xIfqYIzjj3wH+baJQE4nNVT1zJeOCaEeYemZrshE4e2JljG/Nzgq/mwdmE1fhV04
iQq7QJkxQbDttPJmkBpb2EOHVKuWvRTeEE35OQ1xQmvSqNfIgzw+jjPvhHJns1sh
E6jKaHBSFd+nTbDPqudeMttQ8UQ6Xv4lWl/zlSPd/wOEq/C/8JUTnqnwIWLVfhxm
qFWuQ84huBAKRhqzzuYzCgK8PlvI3xGRAlnomEK9pVl2/E902UPqVqHxEIcST0c2
3TINdlyN23nciKsYXPLBiuBp5txnz5YUfZnrAcwSk2RNS3cx1nrMUs14mnqiJEmo
T6fZS4LOSuV2PSvyHogo8prOVye5EPTXXinFt3ybReFTYSqqEOpD7nhPpfErfpMJ
TkJ6gjO6zsopUkmgzdmbnq6jO85fAmGWMb/2p61J4Xw0yV4vPkdrg9s4ABoAPzEP
+7A+rKOHtxPS1t97B1lOA2lQE+k7MemPCI/+FR/9rB93v3znrLOdjYer7lbVKc02
a1MO94hpTE3esDNtSAgTFrZ5G9kG7gP/l/B+k2DAOVy+CcjnbzNmzZUnQzP/xel7
jhadBd1Cu2DeBiuFSByUmgz7pf9MeQwqof3mIgfD9x6VW2gW2C27J1ks8LoI3XKM
WzhQ8QXRtZYNL7MLX+3ez1HgeCeQQj0H0+hMGchnGsnWFuXyteZpk9V3HguCiPwp
v0/Ij2hYucT0CBV9tK60PmlPnhPr6uyg17H2Jjq6YxAXpIOTOLfQZnROBBiN3Hlw
G7gRiGo2g9BT8d08OOqf3+WPBHm5TfPRucFYoHXBK2fBHCvRTbu1PY/1QpnPDej2
uocgWrnxK/88a2iTtgyJoO1rh9USdjPoqzIQPXEInTir9LGlWFsZyMIWbejTJr1S
jU37pEgEQv2l+twmtDlumnooTV69KHJ8RgPsUH+yjGy7+D6IOakm0Sr0ENAOuzi/
PvICjsk4QrXRrPsLn67lS0vwmjaEe4Ai8VvCPWIQGY07YQjDerq3sxXIIsn51Ub3
neFm3QWGXBtxNCKRKKPFTG8MagFsj3BxDP2QpZBqHdtsdXs5xZWsA3g4JLrM9qyF
zA9NyHIDqFkTmMAy4KXycLETOChg3Ku+bFXFfNYsmAAFuOSKGxFwCn0cmFwN2Wy+
K5sT/kdSZKXp5PwuoPR7LHaoTMoJnuKNRZT73joS0IKTeomHeasXTlxf0jsSZkCn
vCLxDrLWkV8Yf7In4hvyyzOqH3wl+4QtRdNS4hxHbwYd7HPvPQ2gn5JiKdFdJ92f
otxImHqGyRR2kxjcBrZlf5qKYghNagHF2Yj3DelqbvCvLDmS3FuCamzbIgKaidX7
Sw/4V5WYpEc5+PSww8Nv8UZ7b7pVu6NREfo8xF76sV0V1DP+PoUgzZrxo1Dv7PDY
yVd34sk1ELREBsoaK9d4s0GV4NqJve+pXY/MVgm5i6feJJhRECZ7M273OCsTTW56
2NVxCuv9EDVki/ii//eZ5a4MVvsDtDGTpfmzEHYNb/ZtWPX6PnCMUFgNUvqtD97P
OQIjKv5rpFP/yxnsAkdcFobiPkGDLtqxAG2R8Q0hKQHPPUrm2Ro11N76M5LoQQca
X6gggHuGD6bVwtSV3CqKFTDJPnJaVpAGgPjN1awZBSnPbWoxnik4eF02/RcT3dxZ
rLv8E34sg2pFFkuBIPOPUlRRM32rFwoy225TlfjVs3CWG+pkL3n493leWRW2hFLn
5RwPIEsgTgQZe13knhBK+DxjipgqGx3pTd0fKm0K6wrW+NVuCCvEE1GMOR7hszlP
e/RNCkhTqYb8FJye1uaEXCKYE/BwjpN3Trmfmvgfo0DPRhbPpNpecP0g5UeQMI+s
v8G3/wnuzz3W2bCfU1dQdUMLMNqQ0FQt6OOAWGjgiCvyI8fLBO8CCF7WOjI3aQh5
m0fRINowew4XjVu4vBmU0PeLwNaVaiZ0MJoBOjeQbRhtEnURnDEp8IAQLHAk3C23
EGxxxBTEQfAlsAPeHgDzzA7pnrh5Dk8qjPI0PpV/tQ1H/NnGNF6jbnhid2ur6yyy
xUHlEd/Iijk+3q3i3zatED73SALlNMeWfvZ/Uf/Lfl/PJQjLimQ930SUdq2f8ZgY
odwHCR5gd2jzc0VW/8c7kXeUgv8vax15H6LdR7gjHOpbbsOe31hWxFB06stWw/xS
rrcGMmcdTEwiKaix2+5K0fWUk1hldRyOMWrUK2k42HmgNi/c7O3FmdLNMeTbdQjD
a+l3WG4Yheea2Uby+H6FGt0hecT/tA/418Hwi28ZIs8BelfG4PgdhbkGlqVRYP7M
bDgvHEI1Kfh4ydSMfE2CSFHSKEEgk+0eeEWsnRLIiybriar0nEs0vbuffX14jCQ5
JyPeTj2z73vnm0Pai8k9+8pJ0BjPZBlrm04/dEpZVUDNiowq8sdZJaZRoA5BVv+M
ey4olEBU+nxF3Ag7qJN/CdMP2AJki+I36n5o42uWznuVjYUNr/Y/SRs8f2pPEVgy
A2Pfr4PRyygr1cCVQBg3xovmgPfE99duScjETbGpWEvkCAxJJo7S/n7zCxm7oMRo
6uxY19PiunNa0381JSEvXc/j2R+zc0aZt+snR568wWNpn9PDIT3aunhtmB1CMi18
P+Mc2y0ESAmNEd+CRdV7e0FacCSEE7155seoX+O9EB7biPrC5RXafFtDGXP8g87i
VPcjGJ+wkotQrz4ohfpWISZAXFKxWP3USiXexWfaszG3f7iM8tuH76v/o+sBdY72
pvs8XZfRpFYqHwQD4N44145WsNy9qb99v1LOjjN0JNSZOv1dbdezn1bXpQlhvnaV
HikQJKxIYTgqIlkVt7X5oEudFH0KNDTzGwqlaIPnKEldnh5sQmFQkL2UCG+Au6R/
7eaj7G4yK3uDbm9JmLWqF7Nt/up73cLCZ0/eZNx/WWPfFST/yvRwM5i377/1XouJ
vq56OWVPqhL698QRrzny6rtTG5Nq9YSTJ5nJtJGS2obg2wZNdoZ6OXK/I7QmcLc7
H/qFNklRCGz2ZRp6DMLYdD9FqNOHYj+lBN3zP3k4Okb4Uhn7B45twq48KGlGB3+R
KDM2s1Hl0SyIzEyF1a7OY4b3vekacq/A0/FaypAoF3/iW7DS4bBVNlDDSHBOqyhN
W7Mm8cJiClPtSAumE6bszWqvYS6IKf/U8YT3VW3jEJMZ2zwRrAlgJQcs46nWx2Pv
jB3v1JC/jTIfcnw4A0Ms9Aj6GC7M3rR5U7e8E19+EZZds3PJG4Gkly07mcpinh0+
hCB2FPgh4m8latgf8IQUvl+H1yDLyD/GOC/d11cI0r4ocFDDKC5POB3Spd0HWmJb
j8YqrKEltfmUKuMayvuVO0G+cZT8lhat4oXKYfYWkoGf5G5sp1llWniF4kghnSzm
v2vtR+DE8vSHa97rp7g4T0qfyqZVAxdTAN4HuETmTWJEb4OLEyUNu+xLE38KTNtO
rjeoOD36o4oqETSbqzcMJKuCCbX0HwNo+O3QOOgX5vOu1lgXb3jc9feSGDR//05L
aDLM3jTTMuGRz+0KzzpgWj2wEBLOIcvpXNNKCIoIkF5LmLIp7VSTWSwq7A7FF1r6
kkK5jO4YFPc7vSuwoTgWKwB1DetPCq4lz754oEjvOgvk3/b0UJ8TqdFFx169q/6h
oT5YEPumA9wHFSNb4fZ4V972R4odYLkQAoC2sX6bBQbZ4vcTvgJ56WjKm8vUHuRP
IG8GiN/0cH/BRer2CSeWJhtSVyynWksfs6HwerFYs6MfIRsZgESOSZ+IT2WMoEPf
KanhnoLN++M2ug5uo+AKzomjaXBug7sDUgzv3NH6QrYqBZG4ULtjMMuqU1mN8tbA
NBsepsYLIHKA/HYgAROpO4KH/SMBHNkp3EGQm/JKfu8FQ2WDwop0SVz/xsB1ula4
by/22TGVBAnC4Qjbfg/vIgK0TixXoK60MkLtOxr76Q5acX0pLR8HrKTN8aOxYdls
xO0Xuh9dGgOMXVHOiQiy0W7m9udT6p8ID4clxdjyIzwvrBwqTio32Eb6zGENCeMT
3YW1abZjxqIkryAKraTRUth8DbYiPNjyNOIsr075jrGHLC7gONuv1H5oBKEKCb1S
qNlHvBHQVE0uoeZjZ5fe/jjkDsKx6KmexWMLINVbnlBTi7vAe3WiynPcJ8SLzaMo
/xvy6dfvmYF/U0YRAAjKswW7ZN5Ym9GnZPfSiDNZ5vJEQxvKE3b9MzXxeCNohQHY
ttd+I6SAnwiRRQaiXceLf2a1cuXVb6k4H0VWgxTK/gbg1pYNVSPkYuY6Ll78Z01H
jBlUeYHM80IRj8B9Pqb3NLR2kDYHDtuD8EJzROMcn9dvmlNzUanb+CzYpPyKJJPE
xEoTlfHfperQYxihrs2jp4T+jX7fOKzud941dkMJ7FzelVChZhgTit2itTLYHNME
OPyE6U/aUoX3lbw52ZE5x2n5pcf3NhWwB4aFhaHG0YQGMbXCZ7g39ikB4H3W1EFX
WpTv7NAm/qV2wDF7515gxGnPJi4VM5z3vw7veIvDU8ZVJgqCJCnFtlDwRQof8bBO
uozS819gkigqpU3FuH+/QxC2JnnVJzZkfgzJqrqRG+vr4paIrhxMDAgU5ElnbL1u
EvmPuFAaGE3bYSfZtjvqU8BLs9e5BCkzAydlQZ6jPjfsoXzGCaTBc3FD9HVD13E4
+ehmOgpYFWml9KBXBxtvGRR+1RoUffv0R4mFH/xdlpZNv6Eyzk3S9ITUxtZErV/p
qM83GP2/XsUgX7O5JlDejsCZLUlVXTWFnfJvmyxeApj+Am727DITd9RMPXE2f5dK
ZxWi6GobSKG/dRbIkSKIMh1RcnN4AQvrALpNe+9gEuFDNVnxiDuI6o8XHBz81hyS
QjiRSOO4OLvu+yGOqMZ+oIIVk2AGnQDbzHtBPQ8ih3Mb5EKSiVsl8BRsm3eHToYZ
ZZPl4e+oWFPMAhVPMZeZEGVG3It8BU3Ena3RX+aARrRs0OBHsGcaFO51xGxmnOIs
N6ZW4wW9qdIhGO/F6haZEijGwJa6sjP0QP8VeXAZygR84fHfVRQlrbSdIUWaac+J
x29C7l5eGGRcgoHQWsGvQMqrZFP68qsnt2+1tOEOgjZbo6DWs5M0Q1JqAX5IRDP7
qmST8aCdj6DCFm246raq+SCaccexPERIQPxtRZITHJnVDYBBDxmEdlBrg8G4pz1z
7i+4+ZxrVYY6Kv8lBSu8fcWh1dl1KUB7tIgnZIf4Yoh9OMQSWIBUDcgCiL56x0xE
np3T22y1SVvdB3U425cBgCFqJ6oLkZBGHK2EyL4eacslt2mij2qf+d4anZqc0nrr
OwmH7xc4emzYyp14DAbkg0T86XokJsYkxafey8U0ZHsxNcZ7Pvod3VP0bGxcO6qB
nplS4V0LCiv/9559ijzBf0RwxRVJH6tiLpSe0xuRJSnRS6tgaGaQI1gYYeEi0ESg
U2aomD80eJv6azsKU8y0Y72o8Mh9GJGzqgH8IyElwW56Pm4XExKKpkaMu6YZjfjp
qNuxq96UXDNizxfb76r5H866LGQH7TQw3E5kC6jj3VddQdxaV80A702mxqn4tFbO
OYOvjapRyapWin+cVmWNlzNEA+/Fxkfhj0ReX57N1mR7YT+oUO/IdHgey8D9igHf
y+S6VuOwoS6QjDMVTfl5Em3i3qvdRq1JELjLtZPgU45SPsFA1xFum0zqbdpXXQ5E
jRrUoSj8VW8hUOdBtDcUPdQ/4GXBwz2SON4rExk8JkzR+7K/4lsBdtiEMcZbeSmk
KEUc6VpMvS8cyiFTfEsuTdu1gYiDmpRHLVnQT7HHE6d9hTxF/0sQuBy6h+lr8O8A
+6Th3QpJ+LMzk8DAc28Ij2jAaeA1mbMQsVmXByJ57PdfuRx7ZxOOateUjQKM1Mz7
eBUSJv5yDx/UUq6xS0zOObfCpA+IDjW4e7baFMmnZhFEliyocDPQ7dXHCUorV1pW
ByhoVHbK6zXbaqLDCeU118MvuJqrKda8aVaIn8Qwj7AHW2XClcJwctMBkk/eoF2h
N7VgCfxIIWCBg+ZlqSA+2hovarFx/MquM6HpCe+Fb30/K39pqR0z33ios/7VrGDD
xQP6eaKifaCg++nfCjb+XZLfCP98c3zXMrfSFNdvjpdz+av1uHIhI/KE3+TV/lwd
hRE0QO1LF5dNsa1g8v78ccVCspAhqG5TqMkf8NSwMdZ2CwtVa4PKTusvddgsGt69
oHFnSYriEsMMGLPsCQA5sk8eqeW3Dv3a6EzRgmjuwhsadJYxQMmRDhw7TitVwN9p
034m4dkYNDMEkkpXFolMpZeQhmSknPbXhlXxnexzvUcSEiy1SRncvzLaTAPv8Fe3
wViTZ5bBqCLagJ7jhUWAUpIRqXfLtl2vToCVJ5tEp8KrtBCXT1HoxG23aPY89j+K
FfclV/tLfbmgk13e5OoV8bLifIOYZcMmg2RPocRVEwAVfNQQHqJrXCfH/RkrHmDD
j+gIVaPyHr9sWvgGtloO2bUreRFF3MG6m97dcmrQUN0ZRWZ3Pfs/kk/WVZ4ZWzUi
RfwAVVEDcDLeX76R4IZrjz50VR3ss5ybElUe7xdobQSd3dJKQFdwWE3ltRsF+xi8
qNMaFSIwDP8p/o17QhDSJUrTCfhajns3eI4EHPiGBIT5cjjM3Nr/lT5gucwKaUIc
MaiPmbe6cNRJTWqtPj2mrphruiEPHwrYmPLCWEeSDjFF7djY/GSy7K+Ol/Uf95WB
8lABM9wVGQiG6kukZJArDi65xK4cc9NMnxHzVgMAriKugTScTg0Ts/mWyNioe1oX
JtRmGvJvKL++pVVLp56XZ/WwcL3ZdUilKcbTrNGx8EWFmgOFYLcMc/hw7ts125QP
Q1WIA2U3k2VnBOPaAjKstFiDiBVhPG/053Vn9EFe6zE9xDOmaIzMbFbV8GKOrNQt
/qmRkdz7FuG4JOaij+GNNXGJvjafGO+FCQxG1YB8ZFn7zs8/6u4RBaA9YpyPxuRU
Pw8Yk5FCxVRuYycYYymoKW7VGq0Xi/uqws5eRLGzZy4EOm9vUOc2jC4me6YKxfX8
f3oM5RAXZBJBfhaf1qQw319Zii0I5Ue8CTjJOF019P7SsLrZEyA+sLc784fjH0w3
kCeuT8SSbZ8ihdbMQN9JbBFYGa9+lrgd7ZtkiUVDddBsY0ksD0TKhGxyJDliwZD2
XZHSsISl/iPCd8sIGT4HrfOXsn5BFwLqxm5Rw2b34m/A+BPhvJdSH/aEwR2Q//Ee
XLfGP+yTWFj6hbDlZUuCmE/EpfhZbSHHnOhasAxGJ7YkJxH3CUoaghibsM9W9Tsp
mb/uH+ClPNglM4LxAZj/v3GrIo9GWXQLydrXltRO0zALu01nuFLvTIQprS3Wr/ph
DN9fyYiX+obgtEGvafOv/FW2+1rIfA/mjJojbjw3QuesdsaqNfcwsCfJEHdHx/Qo
XCsMJbGIab5LS9OkzyI3XnDssu4aslwdvJFk4Nsf2h48Wuvg0tqXgoe2Dv306E9U
ENVDIRM0hcAVtrpggL0syStwFJn+VGwm9QEawdWsnUmI6nNBOAwvZnbSXuoImwIa
os6Xi4v5ibPfSmSbY7vkiaGibLwdrWk24WTmb5LGFnJlgI5iX3vbVfjO2jigaud0
LgpzkPDgbN//kLQRgyrZBt+LkJ2lqpoz+C1lt/jUJQa6lAkuZaJnVaFotmEfz8eK
WJtSEYrsnlTRKDx6F6azVxS+FfBH0jAf8veDoT/T6//6MqQm3Ae20yGyZTwdbjjp
+9Y94Cy04VQnZ7rzVzRv41kqkyYtA8NHvzhHZ8lLc2HjmGzb9yW9dZKcFCGosMKD
KS5ccrTADoTNnnJknttKJYNNLbAtXujTFbYPQe/D4nkrqxYjW5MLsYAhYs/RYRcW
vYujv6laCHHrGPb23aI247e2PZY/etp+1OHc+gf9xdJVBm8osoo86Lg4k7XhANII
jA5XsrmW7n+FlbBH1fLFK3ntK04emxR6iazEkzWQIqH+2zpwFXeTBdaqP2qFc8TA
hQmTUJsYvG3l96OpgOAxfe+qa3Eq/HWs/zLSGNam0QKK98CvkjLRQ05VI+Va6Km8
iktJ8b3vLW/DKom1KBx3gEzVLbSfMuLvvjDBMQTd7DtCZrgNAUSARt9oz8gLLJoc
KSIvHs3bdcMsOypVgK3EotN8wfh20As0zW3jYi6ulNiOg1r5dlkqtltBzaI48Xxs
ZwgeHAqhpp6tPswyBO3Nd7Yf8xC36NyMlzbCSE3uPFiMdDOH5PS2UVErYQZk/8Fk
o6PTqetHJtn/kRlQXhC/UeOIhlGHppqQXIygOU3HQpf+TnwVtJZ0GQx5mzbAg2B3
krljsUEcqeddAOblsVxWlJDbmKy6hoBqh2LL/DLPvgyzmgG+fXOkFnxEcMxbMfh/
onI7Xflcz0J+GK7ySBK9e5TN6IFfd8y/dmCefHMlXJmFs7HwFNwTdni6Aut4lkUV
gA+EvZFS1PPe5/EQQPy3sMMuNGmNZvcyXHA+Su3xRX9YWCLWyR09W2yDRI3leY8F
mbfkPjeldG4I339v184kqYNTcz6x9A5RPTl/aAXjyAQAZnjajJSRYtpSN22oedfI
xmS4vkpcvxEfn++1fI7a37tjUN50IGTPQ+iznYTK+y4Gv9aTaRgUT5N1YEE+Tvnl
oJfEl9bLtP0rY370HBT2URYxYR1Lg/OgeEPx7jy2oHh9rmwJh6v/LuLPMGDR9O5u
aREAQsklAw2GIkiPprVdTGTPjiLvGXtLN5TLSmUSo6OtFeOHj0DHafIXmh4B88mp
dafmwtumdPHvX72pti+ZB/pj6l06KI7G/INYvn1SuwgbcDCGSJKgSkYUFSok5xXj
/0KB2ilsMEaT9Q1Yke80Qz7Ne7oUXFJZ6gJZc9BG94T7G74gBgbEQdR6X0iJIc1T
aCcS0GHStP1Fl+3OcKrPKyPZgZU96iI8SIhZe34MvvbYboNFUZB6NG1YljnoTOD4
TsYWtJrfdFGklxerLEd8iXYDRUAr50JljSSviZDiSq1qwpACVNgIxxAPhz7M/9FF
CWqIjR+JSaoF9vcrb0ApQrNOZ+1LcEdm9hbSfVMM3+iWqMwD4NWnJuHmKl1TRJvk
JsleexFFvqvgIhR/+xmLoDckz232NulbacgE0dIC3r9spcHJFcRpFpzm31Scy3Sd
cyvwVsd2YIUAiaS2rtQElbQUeoBNH8+0Ldz0C0XZ66cx1W1oMlxEiYgQQMI7VkfI
Fl3iYZS1reOS6B7lSyxossKBSpahQ4mo/HXWRMHauLq/ybhtkk4mCP7/NC1L4tpI
UsvEX0XwWwQ1fRLDCWURyuL1KoxDYlmuTem2bZ74KeIk1Yiik9j/TlW8SHIjT6k8
1XSZ1co/0we02LmvGS9CiwGEfMqMgKWd4K2V20sAeywyBFsFV5IxCKWScxc9SwYn
RZW/MSWnOXy9yCSycf6dNcrGrTdDCRGWA3kYknb9AkFTrekJqNIpr1sw81Z7lVch
i4NxiTuLp4wJWroOhx5UO2stAhZOF2+DISq/CAxAsuOg9HiavAQkBAv1Xl0XsNrs
5jbehjnAEc+DhSPjNlaSCn13qiQoN4pNY6/+C+aNCqEwO01YCGwQkNm0+woEpMuq
hivmvquTV3scZUAfKk+JfcHeCnspm3dG4LbOalGP9gQy6y+4lFDNefpkCDB3fx2C
3kq9Yik9EJ+eEv7kdP90mdeqcvBRM9SwQJRdpdCIgwupU4uJxGu6jOG46ASw0Uhv
Tg3kOkrwATU4u4Qji2ZGL2NHSuzP6LNT1bgLD+caT6A5YnI2B/ViN4jsV8wh7EP8
vd++N7QrJArTp0rGz5xFWVuTWdHdC41jbbQVurNSgN2j8jZ2FYKZAFRk9n99W+WC
kyPVyLNr7hBJmDq60t3S5/JUbJqpZtHC+5TdvMh4BIw9XwaSkbx04EPM6AgyHRPz
ImxhXv//8qIKe+5wuY+VVU4th1BijAzixfRM82h86lx7gBEkEHcQZOIUQFc5dtJF
eL0Cgf3kA9+zyPCY4PCJkKtXC0pAuaSeHv/VNTd9ntDCA4d5AtG3d53Dr9KXqT0Q
EU+0NZa2jehRZqlGuqqva5yOMu3uXJXRl2QB+ik02Fdf3Blkw+jC86P+MZsR14Mh
I2zVMMzPUbWujm/trsAos9bv0Fmk7IihdXNepgPvMonUawSF4q0BqW2vXkC6bjP/
FyYWE4RGmhckaOjTpZ7f1KD1LXzSmcKMzbg5+5qOZuRmucmN0YTOKEatZLbqy1L/
wL9VlLkfMOGEsTdjETzBk7z+pWsqta5PD34/oP7F4UT/5m/adxC1oZZXEGqMN+nv
e2w3aGAp3p1dIkeanHGnI74z36KAF1RxpcjG3mteA7ouhqk+DDKmMmqokKLCb68w
dK3ZFIh6QmGNilL0XSdLU37euIsyDn3tnOQXZmLXy2Jid/7OEtIL3iyQbsjgt2o9
PeCZqWbjyf+8et0L83d4nNp7HYkNXPo9gwHmDk2pMh5z0zwEAquzL00Xk/bK8LBW
YDpgUERw5WWKS8RnTqYqyA4+SyGWhR31lnZe0N3YW9ui6WlFnkR9D767aPoA0jfp
aVEEC4ASJ90T0js47Ebi1oi6wsOzBXqCEpbp0xgs3SMCjHVymUkWfTlclRPc51pM
P+NqOnV7vdMmf9VmsqYb9iByildJPgwsE0+jebLh40wMiRa69Vy58FL3s5h9bKlj
m0/WQRklDZ7Brp2zsy0pGHRyRIswotigNiPj7Hg1YktBLg+OgIeawdpvKwBALUuj
4AF4x4gZ444AFdjc5p9henwyDMBS8aSkA/pfBHlYkUCPA4lHmJNRnOI7ZXzQSNGr
oCWWvulVf+Oo2Y+Nw/rGSG/VfyStoi7BHZojcEtB3HlGLHc/3QiPHn4YXw2iGwMN
BPAuZZLpYwFC2wn9cALGaI0QtqLgze7JBXMe2kBIxXDe/WGEEllvabaxFb2Kx0j0
tq36Mzt6QUmA+ECiAAaAYPnsg4Laqu9i7gTWigejAFAKkqTBvj1OIltDtvoW7BF9
fh5ZyPB8JF7mIJDaLGPPmyviJy18PxUchTnk6s5ZxcPUQyDxEX3p/WpRvIVJgjoj
W3jr9JfWRt56LumAklzdBfDvR2/09w0i/Cpyrw0q89CWN36eEt3YlLR+1t38hSBM
C15sCQojBZ2H0op4vtQ0PnM4tgbKO6IoHrR/mHHb8RDtCwTzJQ/rDqnz6krMyprt
14uPYkidAQ/0m2iNyTd7wOSFJSJsmN71t95wyVRafOboEckF/U71qek9KYwg+J+4
NxwklGdVUmkLxgyVDOFPP+HCp91XBhPzt/LxYPimnrevj20DfbJOsIUU5Tve8JOV
xp0TronG501tUJE5arau9T0LBAeRLCyhkkxYGl39t6+VNBT5LawT1xVFFcRw85ZG
G/Fza1EdAYXHywXLiHcC9PS7tiONzGQ9dU5kwY5Cm8JFbzXCiFTskVmuqPWn+XZ1
3pfgAg7ZOH0nt3yvC5x3DiWmazNeA0IwRM8lxGYtePnWFGf4GsjgE3hjV1a9qVpT
WQY/dpP8xkGF4ZTKVPSuNRmVP7l37cIUmKN62eyEIOe8v/vkifUfVjRG1BzoyWyc
0E+QPtWpdlnpf8feYtCZR4b+TX39m01tuzpRgSzHESKcPXTDiPMTF5ZcG7ZlCULe
MQAJMfaXgwFUqrbO8kEfY3eVGueGq4mzLjs+608+n3Uj7HaCvQ53/aMT9L1xaJZ3
jjh26VAiXNHtcsDa/wBYjZhO2TmPiGUZq5nbwGzRlz6hizj47FQIRsfbLlfbzlpf
JSHuA3zGmY7ZXhvrl+HlWg/r8lHAhXz0E60kcG5euuAGeU6R2ZReDzJ6tHeFt/dh
ETmQdOAHGdbvEn5fBFkmye1iaUFLSrU6R/e4nKyJU8eWODYgn7w1H/pIpRZCpFxw
xAWwDxpAe1OedffUVLDApQJ7YatLA74UDP+Jy+PKGtwOBtCy3zrII18lcbsUSRK1
t/aBiq3uEyevw/uNw9tNXFKvopjJG4zbwEn++1zW78DsaeOL36OklrNZ94Fa99Wi
kDlIlx3KMFkbTGL+pVOrS7NkrpNkN+d/4rJv/Wcp1NdyJ7kgChHlOebICO8ctRd4
KKglp0bYESQlq2kCzzHkkSPrXKCWWkSwd9zOqe96BpTUPTBKZZwp51IuaHTAhTQ7
9oQt4JFPY8Yf7ztWnm1Bsfi0WBDvzBxpDSIovYfHnd60z9W94BcrTGiLeAcy/eDl
IW6vRsYhCWCQseSh/bymY7RlxCjt4JUd6HKsPeMMeUTV5S8YLXXTIWINIq/EJsmF
LPax7OlMDTo43FP6uOOAANZz4n866MHD+i5OziZMEwx17uAS5Xi0X53jj8c+SbjV
TtceT432fIhvDH7MeH6qCTpGEqkKMNsvrslVgqx2TcjF8O+yTpY0elWThe1CgVi+
+XRRTJ9MEk9GvtDDV/JtaQeI6wmiCFupNIT9qzafBJlEA81s6eDUvlpyJXxbzUpY
rP4obkkz2JuirfMCE5cMvXhh4haqrdUGpfsugZZlG2t5/osgExUGkpy3JPyLANoV
Pb47pAtF04aoMJpff0Fg3j3tfiaklB+7yumeA3JiaK431ra0QZfo48Gnf3NiLjrP
Er1WSn54C+/nZ36gJGKE+w+OJBPX7UducKNX4mogTyaIbo7/HcIRQCWp3/ldzxVG
PwA3vsEG6uJ4djxoiL3hMDy4Fhz46bF+MYKpj5IeRwuCovixDtYOPHQNlReITlF0
3IzcP5jaKSDGSQomgXoSPDX4XizTbL8m6kcjD+8ZDM2XxeQdwdksSWeeg5kYA1bC
i6Zi7N7h8tIK5bNDmljXuE8m/w2hbV3V59jYWLzhWy4FByK0g2HASEWTTyAIyRkt
ancZXe9KQHhZohVqjRMDYIllxi6Mzwbp9vhrwVFP1e2ttja/x239mzdIfUCqLbax
jzfCB+MopknyqxSNQ9ydmIXu9NhkONY8IgdYzEaCDiO3QhgOk3jLSx50g2liKQc4
IfPvvgOm/HZmfKyhkjKF07WRVcvufVtNoVPL2AE9F2JIkRWTWRJRQmobSYh16f3W
3eto2qrLjUE1/fhvLbVBGS6yy2MqZ7e9F8U2VGTJaJWIbWRbB53SrMBDnsTOjWkh
p3gVUI2d8aE8SnMGaxeOWNZs4QWNjlmusy9VhJB2vJwXIOEAE180S3TK3Ug941r4
TSbtHPzINHRRgLEx0dj0BpEKdiA7oPIQuvLNughDyDbRx9y8BFh2MHup9PO4qpdl
MsRVPYQLRqvdnJB7p/NnV1vEJK6ja2EaBFh30DFvE5OTWf1wAbjVGWzHv+sOpsVV
RaspYBN3jXgC+DQLU3AlONJqkxo7S3V2qW3JStN2CP2LlMx8HtHxLdszHuO2hOsP
k8G/Ydwm6mYRKyoxFsGssRiVmKyYYTQ5nXQD/3oHoj5fgtdWu7EoL4KwLJxoQfJV
2v9ndUs4+UvNJRvcRYStn6ihJPWEbwyk2V4Zv8DXkrT8Cxfc7qqfdCeWirlXFjQH
p3RgUBuHZ8cTuN7i5JwDZuIVCiy8UEljnBiweKKC6bLYMT/j9TI4g0MAtiZO0nKD
fwiHTEeRsLhdMiZTkHm8bMTUDfHlAkhCJh3u8CqJ/R9pLkIPV2u9C6+IJlmLpUZ2
/tHppQtP0DM17fQC4DNQEDkLz3QMC7wKpOLgmspiS404WamX9mbVdbS1+Gf2U7mB
xPcPcRdmxOXoF87z/Q523t2gHCefrQ06dqi5WhkypdD53lby7eo+b1P9MR0uZz0A
No95eyoukfADMlnoPIXggvtTty7JfPvY3Ex80HaN6fCftYH8SjUXWR7sRbK9Ti3u
gjlM2KT8Sbm/g2PCzhoEIovGbMDGa8fjz7oOTGMG+VTVb0GkvLdQU3RP6nn/9AAM
9RATwdxsmjNrMFTG7PI7cilGoEyZtV7Dn39W2qItizEnj9RQBLmt6rhxrg+r+eQK
CCBTUV/o7fH+fBvSNTF2CNv7QI2Z6vQHVKO0W0UnAjXaUhc+O1X7gdG28HXKoxf6
8ktRdlO4uu4AJx4sTrPmEfFsdcSUuwwqIghmV/kWXbST9EHRiK4N9ERIZBxzZLSy
aYDv80lVNpQeQ4KWZt3JfKK2z1mAQDz7xcpR8IdhrUVOoV5m4nwUp3N/k9KOWvNZ
h+f6rO4m65rI4Yd7ghyOBF4KPoyM+eprB5pdUznJy/klS4BhZwnJqYE1XoaTmQWv
Equ9A6WdO/jnvHdMR+PPzT9mp3ATBY4FmMo4FWq8JPWHRQmout7fxzvt4HFIKxOP
IWkIlW4eKWjuovTQYvBdoprvcgxEmrwiNLNSiU70VRlb0IWWp0pYms/bbRuWyeba
aHiendwFVEQtzzyBUruF9OePD3x3bBdqvFVYPJMlO8qUQAW+9GPKH0tQxq+GvqBL
poUaYkOSNL10ycUh1GJeB9yANqdmTeVQ4/PAZjoWruBpOjPh6eP0IiOr8wXR9vVp
hW6CwhMvP8akzqPLmBpkdxIwxh8N+YbdfHVEKGgodovLdcN102j23vjcEN96+LaO
WDzUF52mI301C0o24INKwSiZ+30cPq+SrfHAdysUAYk+kJvHNGDXwaOVyRZdP0S+
I4EhET91wf9xaRMoj8knqNyNIfpsT5ZurSRXNbhKH1YZn/Gv0Co2V4bZZgYXd81i
kiFH4SOfJabsBjv7+Q77GI2H52hjWWV2Zw8KfrfEh1lMhhLSUYx62I3Oxu5JjDuX
yjS1eQjBdNSkCejcn1TxGYBdBhqbq1iCZBIF5E0ibOe3rTnAWYbbPuZ5UpQoPwJI
Ftk6Vv4cZsaf7y9u3uEsSQFTJybEq2Vq50zoccE4fWhvSUFJfZ6IXk5BOelSnqzn
YeRVDZaWL9XDlJYO3gbg+UzhDqAhEjlw/ZiDvTMw9mub+N6+cmOFRhzcUKn42iI0
qMEKdfXTQmT7qLGKP9Qk5nQPUE34dXNVGRu/TPRFHLHkb7+rSkimf1TXueXQw8wM
WuN8+SIJcW1dEhy4wnkTMYVikwrNEa2uMrfJMCRZlWXRZNZPh6LzK4//wglUomaq
lVaciB6q2k/e3xTqOvkoc5Rf+/d7dkxvCI3yiEYWWicCyKVAKH9RJjw/wkvtWmjm
vB8qObsWr42xQsmypGM4os5+bVuhP+Z5CwIBiUpXDXDXYaunW5qmtpGz2C0k1cTE
4jaCylkvmEFh9HPqSnZBROdGLfoNyC7PEerw9G3OLrRvozQZvE+i4XgwgPERrc0T
DIfUkJ3rZJNu7hR0SmB+ODpDWg9cJ5tD1VPswZrfXV9DBv7UZ7VlS8IivJJZju8s
qw07HjFOeQDUqDsw9zSbpzcekPcjXRallwYb1AhzTDUe+EJGji2die49TUN7cmd9
GnGDwM1K+TQKaswyIFYfHIegRY/079Tg3WMg5ueS/SkziYic5j7YWZC91NfXwOhS
AwFGZUBF+rYEJ/KUyYv97Ylv6nxD5D+dk54qJgpOH23tj2htdi/5s19ckBr43/BI
TgqQkm0HRrHFvNYmRiUdVvRJXsSaDjVgGeoJoXpP1I27xeyGmohVBplDMpYRFOwn
7aa401OP6lqFaWhxVDrSJ43s6S6FUlOZ1Ea1M99nc9WyD3J7lcaac7SZVrL/RJIU
1STZQIhMS92AYjoLHB3FKdobRtXEmdUumBY+0/9U0gDVdAT+8EdjnNHQYDHdfnbi
uzILOSWsipIKwOZkK87gFQN0BWcZPDVXmfyYPSuXjChCLrpRepGRinM69NUUtWq9
lzSW8xO0AxGsOXaNrqyUlczF/ISEt4gaPA7bT0XtyecE49irRf4kQy0Oe2cpq8U4
0jEcrjf0GEHPz3TYmTR225Gj5Sqs8lOkQrMYFPfEhgGGE7yxFGMAJRXs3T32X+tW
IGT9E0IVbdfqPRuegnFYQ4208PgFcN7oZH3FDR1ricjVHjyezeD2hESQn/Ibzu+y
eWkXEnGk/ejQNb9gjMY07itF3sYPrt+M9FlXVycbeoyVv/miDyppu8040LgxXCai
GshqUuIgqn2BNGLZJZco8TjTsyTzJeADe/9dmvgqsh9vAHGpFZzoSFbvGZ5eBlCL
Vcrkakvp0QYp0XvALXwHLEHzqIJLB6LW278FVuG+s0Ofm6QejznMRkZIJBQpvXBv
+q5HN/7U/pC00bM7Bowrcjpfz1v9WJJxpWvkQ1Z6+5vXJcaKLDQKHt9LJ2ePEKlL
6iFaxngGsdYeQ3M0Dp9Cwv5JBR6PcQSC3hGSMmZBVLvvpqb52f4XWCCO/6CtzU2P
kc/40sa4RZSc08pwUl2z/4imgbHdY6Q50gv2JTAM+j5rksiOkftKjItM/v0v27Cf
XMQco/Cb+wW0CtclU7ml46T/N4aRuEG1zr78xx052L0BhfTg+UHhYdhaiiKAs/UJ
cQ26eW1/7dL1mcsz2ldcHVr3CoGI/1WxX3lRtDkyj+O33TMSqSnkiHMWzuIr47KI
q4HW5o47lD/TJU/UKQOakGIPeMLcJaPDOzhxAlYIxB7JYgDMxe2V9An6tU8QjEjr
+wakFw+2t1ZeuOB7683uGq1IBumwJfpUPUZtWf6TMGxxMQDW3OqE8NQXA4lIMxPJ
D+7QkqPQgUTvU0tFQYMM5pt8OTSqcgdz7FHtrlE5vwJjXt/39o2V0g+BUjSRbW8c
fjbXwXHq52HenRAdZhs+4CYsdFmD8LdY29lFVxX456SAOXtLcc//AlMoLJ4W+lIX
v6r/mBEOiHrNSU4fs05jMFFxg59Cy6LGAXwaOo31fThwqOsEVHb9pIrbwh4b3YJJ
5r+lg2NE66OfQWw+Wmys3bWuuCs01vWc3P2gM1eoWZlh8KsHR26Uafic8nhCsTTs
E//aCIElAmwd0lKcmNEOA662vwqaX40hE2mwlSk76zinru6LABYa49VelKMoQmKv
sdXDHhrgFsY4Rah406i3D+QIf7bv0jZGkJv16w8HnAvBtecTRPULlpG91DFYAjBH
O/6Q8FqgYPL8WzYo7ODmGgCCqCL9ZJ4Z+PQVGw160pawGwoi/w3HxpsMddrvA3A9
fTn4WvmhocGOfUnBPLGH4Q4srMpO+CV9CGX7qhq8PvPkKPZAXA5nTuumtFHvLbEJ
RfXIjom8CSvFIaNOXGxx68uEsvJumW8enOo7pGWHvKejXp5R8kKkucbvCYnnFhKC
BumzrTW5Xb4CifucHhO1R2SlvKQeVlQz3U0Fit4mZPNopozxGKR1SnuReoDsZPSo
T3oUvY6NrlM5OszGkrDrcu6Hz8Ka7ON3Hhtu3xhtkgaVncAXyr9+6JS6qKlo5WfG
Ub/6rKrbrjc6S8FilgEalviZkFhd3qklRAhNqfegAdm9J+wK+6wxh7jld9vhRx1u
KE0mkoCk4X1OfGTQUQKnfXFQAATcsorRcNkfua54khn7MzTwoWo4dxRY/kW4ihYn
/t9oV5lDt+vu19zYa0YMIHkLzHRi01R/h/hLBp6VYoN90yulH/6ota/FlwsXogUh
DxQjFUwo+jDj+xBEoKj5IHHXfYa1F0fkWmrOE5F9posm5yTXZJUxk5vr3RN/xQEi
Ex646PL42nSdKWcdPYslBMTysZRbwWVosyWkWe+TuF7dYmZgkvo93vVMfnlXj6kX
EirPmBfdgFPdwVfmd/0/hhvviiRDOnk0YrJZzqsYwHlyi0Oha/r214Lcv/RmBSDg
59ibhfF0TTv62zNHVt7RIv0IxTUhhIadYxLLzDvSXaDqUWXSjT/2MWilylJHTHem
s9tFDsfhJVsQI/+YGp3Mn3nggMSLRCdMtHAs9tQb4JddAryStiq5eMH70c6e7zTx
KEfJzQw4IDCw0lWB96lSWjPBX52/qFFtYhBtmmh0Fj2Pt1o9uCw1dRK47BbyZ9Nh
2nVcmhwc+vWr8cgS2P4aqB7dc9AWcdOcY+UJdXqU4EuxC0Ren79faexNNstKxiZe
dCM6wjxlEO7rZndPW2bsoYQg8fUYnwf9ETKBY4ETsQCuuLAQzBzBchvTA+YErNpi
rXhNpOF1NKgGbtvDoaJ597LVxx33uSa0NTd52UxMSLSb+CmjUtqJNsGZp793CN3h
P1WwYblxjKPluTVDUs9UZRG5XWOXYID6syXnK5e+jSMUsFSPQuV1NKbI43D2cAdH
RNIoudArr3RqDtYKz9g4Jd75293vCfUepccNqWJG4DtdXdX/PlYhvt+2uxxzMz4f
mwqcSp434pvvFguQ7TVH56/qFMNWi8WOkSpwW3/CbSVkB61UzsWTZZsULRutv4Z0
rk8dG1QTNKBrArslknfQOiZnibl3K/i32wVn9oN6UxoPYL7gl6VcGKKr7YJuzcFI
U8ySVWJgfn3sO4BjwVE6hzZG/RSOtrsGROa8I6JcKbrtvAtiPQt3IMdEXPWWYsOU
VkiLfTDRmWUhtTTNWhXP0BudamENr2iszDVcJvwHpJNuUVfOu0s4JeAm0vD/s29B
kldch48IFDop5sjNpaoQ52sDcWX2JR3cAuLGUv+obCCLyMFMrO1GstLeONrumx9T
Ht0VxHHdeS1PJBbWX7wJLOSZjwtENuMw6WMGQ5uRTRKwzYJqfFLYXl36sbNbSOsE
7jiYTAdLdylWwhtY2LAiij9zWyPMVDkiw32T92yD2n/w/vOp6qrqW905c0r6e3PK
vX0dMrrWtGdo4XBAX+17N926ZRbuw+NuEkqWE8DCoKr4wSJPJQXn1U0VgcB750s4
Lty0WEVqZONtko2B9e19yD8GmExE1genyXl2VnCyKz7rnDsA0yVpTC7VfMpR+19C
ndgVdHcslmrERp38SGljZYmz92xEbaMr0C2/2PJ1zSt5lO4WufhaOzyut0ZVCZhs
aqEWb2Wdn/hRqjbwToRIpToAeOqdud623E0nbmfhjB1u3g8rRWZlxMPD5/XVrAtd
9WgmLfuPpnXLFdZGIaAWCSKfjqgm1EeqtAPhqkjMPJPUw5y43txxPs7q77zaS8hX
FuRSioXK/K6wxXrA4iWhyCr6okJf9RVJ0Cp2Q8W1viUHy2Ch8+v83CU7JVsPDpm/
ebo5tHQMS+qwVEtXVMsMgEdhoIA29mVSPfNuS/WuZ4jX3DR/5QwiZH5df7Rqkjxb
korRDy0OrKLpgf9D0Kn0PdrY6EnvxySiKHJQ6icYPBp3HqmoeVH6gP+M3pQYAanH
vHlDDDmo6oCkC9m8M7YDMgQ2eHgGRDRUxuW3SqvPmDKXP1gNJjkVrb4PR3hJ7WYq
ImHBWHjqavPZUDiiWoY8keBg+/iF6O+1s8Q1CFuekJRdv+aXIT6jIBQTfJVWMXoB
CNzJV+A034U5WZq2VQH52u9hwgboWaC9iFeHYa/+8+OmE2AoHSU1L9Zaur4VmE7z
pp/19wMVPphKp1zukm4qAxkZFS4a5BtUaWnpM83MvuymmDz/tzwwmNcqC5kFQ9pI
/bIfobSBKihN+bYC+dSuCBABnJ4yDF527UIXPA5iwfbS2HW6ZHMeIOe6gDyoI66u
H1vou/uGn/Ai41BysI1AcDL/h2aOkUmXm7lNhl8YZOxAExm+XOKNTa5o/VVA9RZ2
tfNZD9QkwQc/htT8svI1yHROVwwrybj2mZPQO8NrSkjlTAqXEDdpiz7T034fFJkh
mSXcA/4xQ6TAtQyJ5fWIXPiB0nyjqcIK+25YbAtXc77SCKIuZ5HZuUMtlxFHBJkk
mFWkh5y6CCnJpdiGoQnVQ2tMu5yRQldc1rLMFueEUUpYSzeQ59tDphFMQvtymeWk
7N0d3o4cu08zsEhF12A46C2LTFp+SKCvevOUTQurwH3y3mHrs7G2P99chTXKJczn
I572mF8RDfBo7jkbosVgVh0tB+Wb2il2E4++UpphFNC1ZqkgsUuqCAEDrTtUt4pW
1s6NcTiwP/BnTfRJb8RNz+yZSzEF1JYYGMdfG1YKmqWFLLW8ZD+kOecaBqCJzBQ2
PhkJeGvCTQuRTFlbP15+VMABWbn6xcdbRZUiVcLALzvXXp7gsiIBiQlJ3WiB7r5A
PS77Kbl+jYhWgbABsKqkiKGtXJdv0o2Ty/oaTm2Ysz9zfs/A1eEP0UWhhL2z6y26
9YaTVM4HdTIrtqfgIhNcQ08Z14zoWlA5XxVOOFKwseHREnQs2jc3SDvdd6wo7wyI
dJEGIQArN0WUHr/RSZ11QIhMieLAmDUpkP3WfgzAgMLVDOs+qhv7RQ7ZLMJ7bMDE
dFBvgi+Fcuz/hpiegzlxVFBNP8rLltE2ykb1zB3Fjr9LOTcCVeL6GVpMSxZ3X621
WPF5t3ndGCLNIal1G8/O3J4ZIku3zp9SEhFRyFVArKW5zLtGODmCNSxT0jBZnRbR
ewmCgroFYPz8Vh59kKVoDNLhts4PpjrDItwniTP34Jst5J8VCd8OwCKEJaJd2xRx
iLeglF0rBJm7C4C/GfP84abk2x4ua6BiUZLwzy+6E308UtWK+2mNCPuVY1x7BbHl
yBmVYAIH6gXMOrL2uV5H1/duNnc2m4MzSwcvI1SY49+GnzH9b2gP42kQzIi1S2sQ
rtzWavzMhQbiCCUDnRTESnGSlnk7UXW7I6YFevR8G8Wv+3Mp9K42E81oGedn36nV
+r7bZQsUxrlqEztS3vgT+IZDQ/aqEkXsndN+OZiBEO+IujMt1cBrG7ZO81h1IG+n
V2rXX8X/jwua1z507FygexzbeHlOJomOf+oP8YkGFJc0N/cmbaxL29Le3dYi8SAB
6Img6jvqTYw2iTjdiSsgiorUIOVqqfKYYIb+ikDW1HhlxSvRRynVjGPqMaiII/+A
+aw7TUPMGkRemQEjqX57Nw/jL5BtQ7Qa3HTLOb/PoEzCzMjL2A+vRQ1Vq6ARWGRT
2QNnoRAEgy1Rr43aMY6Fbl+Po6JTPyKqUlVEJJWtkXHZDwU49cwFHrhPk2JY1JZ7
5n8SX5dL4iP4bjIowf/Mi2ZKBK4rR+DhqaU7A29/0e391QUfxUZp7YL3TDvQyZ9n
EWw9bIwVnMph+tYZ7XSavLZtWMeaI9haqRnX1qeKz9jabYQ6f1EkjwDVouMvRgMU
H32pnxEOekRT5cbzFPjfJEIBoQKTSCfGNthGi9nZW+KikbgFTCbuUqOxaBHsWR7i
/3feOjSR7tZvYCTkv7GtPlpa3jY7BJfsxFqtX2e9fy71o02PThq1fgicKLe005lO
yjwvmlJJDSBybWProuhI12pVyHXLyu4eZzUdJqOJ4j4lkpgyLi2701YhuhS8Y1fp
lScSM4QonRsar3zbV5mYfL6Isg2ncTtDeUHrFao+9F8mEnuyXJVv3dH54DmpnGqN
RS1rW/NDkE7CZXwZ6Y/Kw0v3ujQz/RokJCud16qqmVUaSwm9epzlgNeNy0Q2kVeM
x268sfL7nxyH5BLP5kNlVrqabUxQaLND7+FITb81DHHk3WBPzNViqDO8OrNC7poR
7bw+00+QlmHqseo0Giz6FJhP68ifsAgJNAXNoA3TWUsTyY3+rblM7QsbQqU/F13C
U5LD+1JbJOHhrSDo/sRte7q3gCXPNL6w1JfI2lELLmJub54mcDJaQRsX3eGBRQpj
XYizx+pXLjV+k4MZhCUvGdTzuzkVGzV8ecjap9xiElZ88DCEnmmT60AkK+YRGnkW
35H9kOUAcj6WM18Q6lBqlEFvVXhI5JC5ClkxeUbb+MIoqdmdTsubV/sv0MMjr1l0
l3BB+zJvR9IZXiyO259r/SEKPMDil/wTkDIleglA70Sq1u7GBtx7dInZnQsgcJkX
UBAF02W7bUp6XKxTwB22kWbvOCuLqImIUBrweCMr2ifcEwD4uNivu42Am7F+lzY8
mgpZUYdHTeXPzLY0789HRCStqFdUA7EBI/6fCgQL/u8/qmeGKTepywl1YtBkZX3x
Zfy01kS3dyFI+mZfpLas5X9c01qxA9oKt5s2YFRQfh7TS3RX1dKAsRi33dhXuApG
X3ljQAj0/BXcUG2LPAZ56RS0d0n5JZaXqGeFC7DG6Ozth/Wn2DP3RB6onj3nRwpU
bRFpkgqkcADjTK9Iajviwo8/NLOMoukD+wvDqNaaZWPmv2j0EV3YaVysX8PnUblh
8fFkUBUKtN7sp6fB7hM4ykDt41WhFBdVJgMbHSVrvq9FHYPQqOD2K/nncj+Lt5o2
LUPF/jJWXoJHThlLj3usZr7AqCD0W943E2Ijk6z1lNGqCy/sKgBv5T3HaVKleEJf
HsXsmRAsYw8RldTnjx8Y3lTM53PdlTt1HExb5fdoGRDTZOV5RsvXdinxGE+2fp3B
QdC2Fj6RPZ68HCCIeXaB80C2SeBegPpc/ftWJtrThAt/38PgEZ/GUjmYjiwAlPo2
I8BcOS+5Hwo+YhLoocz6hjyChjGYj4/CuqygZyGbANS9VrwO0RodFVMw1MT+t16m
ziGzn012V5xaM4Kc6uQE46C5cECfxdomK38ywhI6vtQMLfn8G9j4BUq2goJPrN0R
BtYRgjnrCTBXs1HzL3co/I97s7+JkKgK4Zwk0uS59EWrqCauYutkKg9HuVs08Ry2
35kyUaCFohf50eYwGkxLY3NheHWF9+cArxm7FMig/0tY+o2iUUk/dHwE0dVc2RzA
bjVKDye9pa+3LagO39BHYXxFRpcAshzL5Lgi9EKepKLZfDlmCWsYQm8w6esZttxJ
GgkcwXbuwT3SOkjF2/7aW252JCimwA30St5GyAZnyrEEHMgIvMFjBTNf82FBDrd2
5Q3rl7+gN+AlNOtmNsDxhLJcvjBCtplLZi/jq+TOWYey+n0l24ys/ZmGiNkkMaL3
ZQM88F0H1RCZrtHrpJ73Wp25P0KoiDnUw6ObvPCzUWUHwKd9XN4SJyal5PYRCjTy
Skv5XITrMrFKZMc6aOI8Ys+sxDlGKBQ3eAOnZZizk1N99p84KYY5H5Tcv26EE7c6
hg8rH135ZQLzYfGkIvbBZnJAQZf0xIpdu59SCgmK0Ws/82wbSHmI30wKZwBs8mVF
X9s/I5gwH3TlGwJQaB0NDLxyj1ql/MWILvzUAtFDv9mzEfMiO9QWYLrfyph7gzVv
Emcm2uDWwlnjSuZjcsWpSF+luEeyCA3PI6XvkvdEQV+O4I6gbiWv9xJnfj8jwadO
tSRD/s5GX/YY+gQ6CQ0ATj7iJIftkVJZQQy/wK2uxHNagflumQJyT+kuVDph6Q0X
KJI/eBNLFj5Qu8ihFDlJdMgiUYx5Y4eBs1UWrOpdj1kTaHw9cksRCiGi20qn8aFX
9ev69b5iOaCyv29uW1k5LUVy9Su+TAQKJ0WZmZFl6uz/nvgU9G/911ewFIH/ap3K
RMByRtxaVTFd+J//lLTq9DtRRZYeAYGnEIPZevuNxRl115DS4sp6a1g45Xz3ZGwr
472kbYCMv9diOJNxBNmf8eiQNItgpsESgjEQ7gg8SzOcjuzkkinyTSyd+xVmTY/m
knyGRhSeaLFsn+P1zG4h+klA4PiKOVPNKfILrKAFj2xtrojjMMAQ5eSE7VqEPipR
/gUYh8hmc0dh73RAEwwDpDSsmfAQU31ewDXQXx3LZI6rvHs6z7lX6kj1oU14Tjdq
d5ieHWFtUbYBvulIAXblR/oWJ5YSR/0pWkDtNlt04oHL5riex3a91/TmvOhvl/5r
C4A+Fsd3lrfg8VPwhtEScTCSeqdkwKYrgbvecCjR87GnC4MhQbISXth/zoPqRFvv
MHbh0xTZ9WlRjnBLLqImf+7Y9GVYU+9lX1b4HJQsn0ZitG1QQbNWHusUplSinpEL
HAWIfLu3VHqmk+8AYsVR3yCdBDxjKBrsqrqsuVDmM6fSGW5W0eU/51sVIM6g0qBO
UiOl2gn+D17luB/vXfuyvOVxabOdVeeUjfumnSaeziwjejhnEMr3+73KjaNqXPRw
HRAH0C1ppH+eYAAcpYKKkZDeWGjsrLXvvrrklsNOKsJTS3mCL/or+ikQ0wim/Dzb
jdWxrwNXNAVEA/YjtcH4njBwTqHulLK+5xOP4ZsczqmMXaEUxBVLovR0KJGQZ6nU
uXCxjRBlazvTldrB4IAGJnjFUHytKiAyEMk4UAzothh6f/2YtDufOzU+4sM3Ja4g
F54HOiOHnLJod3QUJ5aVCARgMlNcV0QhRTX18U9nV9+MbDHH1c7kwm3sdfqwh7p5
KiFKYwOPr/RkIbSwZNU4mVIMsCA/mm/Jxamm7YFHP9ZNjM5OpPTCoe0IW/3cpydf
N6KecMPFO249Fl5DrGP9y8WqWXWNKSgQLp9hr5bnqLqnYxgNftTfC5hvlf0r0Fv8
cUVN3nJzRe9ofrVdAQ5Kw8tqrp9oo5gfb059vCyIBIF/z5yUFJ37RR4HlMYbDEIw
N4BG9Y0uoyFmdhuRtisWMRU9FGpgDUUub6JZW7mc31mUT5Ispkl6dlu9YmrSFg47
0XRvDGVc9SZYAsFCE56mpkbNLgEiQNnNJz60XN9bslcmbX1l6ofhfCjV89G6ZMMM
P0To4YtwrwTuVdigRs5kAcZyoUnUTvPJbnUoOLV/5fT2VS1P2z2a+Ymk+Z4n5sm6
SThEH1ePjFuOuao6B9y6lEhvhkDBPg49gwTRct5YvF0Y5SC1mdPTGo0EFg+p5uhx
22c5UEIRQzLTVk4Zrz5mesnpdjii1A1fzV5wEV6WFeLlm6dAAZoQvkmw3TSyQgKU
2y8moIltFJTYPuuiWWWCGo0VG+1Z3TPVMhBGs0v2vH2dq9mmWxaA98QBnVIMHKbV
lWdy3YCkmltIAdlD4xqSwgKrHNEKr0RlgYjRBTuZGECx0ShlygBvOKkIhVWwCxM7
Hyu/+K/WqVZSCCILE96v+rexiIGO12kJSYoXqhKXghrQSgVB24Qoi73YdhvRX/7A
+ZB1IDjzaeDXzZwwlM9tkWyl1JebuuFz7VBseUu2s+cevEZd3FCk0ZPabsRlJKdo
7hb+jaegkVOeR52QLCYpPG5QyOsX2cDYWcXMRGgz0kFCBsLB4JmPEUdXfcZNsQg/
mRI3Gs9HmvW4SPKIfcw38IhEvmNmP/0/YU8kJknwGqoCFFZrnMQYbng83ix/0wx4
I0d9ixskbyi8gVRDtrNAH9blidyQnPL+cplHFGAuJSvgAu5yMT4mybqez1gOoJT3
9WT84TQVKvODTxz5r1t/2CxIX8NChyNk0Hjp5+J1q1rdzPCfG7weQyid65+zRiZQ
ami8n6OzkjPIGJ0PtRD8kYtBb4U+1ilGloEG6751qyM4cOksDSgRQR1ZoIdsyMOH
dM7fu3iFXcx+F2lJJNaGwACno1TORK5hJVXl7EYSD3gNbExL1OAJWzDGiRaLXW+h
sfCl5Sv/xpWxpOvnVpnOd2/P8IWY+FJqi4K7dWYe1AGgzNzbx1JBKgXeFoMi9sGM
MZCeJmgqJALdh6sSosLt/2/hHYBgw4UTZPEGRBE2i0dULlvQtiHcaSHhBVskJMWP
sfwjJdfOPbORFkxBNnPm5RsEwAd7D8hfrcT7MhoZzq5Hs5RKD5haLBckRzcPRk18
teg4sFXCisR3vrGgVcaDvJmoTn6kMiNVEZg5QdHtbtezysljN7amXZlRL1mFq9CL
hf+Y1wHIK86zOweBZk/vJYbsil9/0YFxOcY7Xb0q8n33khWFRgGWUAhip3Frj8Af
/a2Qv3yEv8/WA3gdYqc8KMNjdzui435lHEU7DVNoPjkVxIVnhsEDqzuaOvyYg7zy
CNdSqlLlKdg381y6s3TFahFMioZD+vI3urNRcM1OaID+UrE82Jb3I4CCjwPKnjnN
9Mjn0JyYj0yqfedvQkyMfoTuSWnEtiCuxwpi9TXp3rfued8iVSwha4T5FM2CK7gK
XAPulp9gnIW6eOeFEO3DjbBcwnPe/H8pi+jxaVoZTnGw8Saf3hHrBzEaw9cgZ26i
6fh+hGOlw4z0YURTwOxoQzthBDCsNuig8Kuwgy534QIpOMkKg3wfEyzcCGv7m+1Z
tHlEAaeUt22XPZIhDCnsv7Uav9RfsuvjVJVjAslgW3p5KC0Sv3sNeU8Q2svily88
InI9tNizp3QCIA9jhs/jrmnSRO15K8W79UAgCJtVpgIJxrhKYwF4Rx5P+oKN+Gxi
d8ul4HgNqtb32yXb0WXXX/TPQAH1sCUwqwcrBBJF4xxaLdb5Hbj48Jy9+/tyxLzZ
pUDq7NWWFKeO4sbvGgsZDJt57s3CQxBOPu5hHrIvctZmz/PeHY3Rvqxa8ia5k3hr
jeG7K5STrPo0AfmH524XSHS3N0T01J+3deRxhtx5JgLDFRKwQEz531jNT4GxaZZN
BrOq79jY8ycY5stscD8whpJT267u0vRW7FB3slDqA/0aKav8n/SyhNMQBpGSr+Vr
oTqpHvOyhvGTqtU7ay5DN6ZhLpLS/jLKPUZQMz4VAn/o/qqxeB2pKUsRP1NAy+Hx
5j6C3OfY3HDuBbTClshnEe2GwhGJW6KgPuBi1jN44/Bm/B6JjTlSlXAJxkJaTFqy
LqjVa7cnK1caDm6/3cWeCVdoQgegTXR6K8Kkx+Df4lEfWi+gV65coj/yroJdJANS
izoPfp5NeE8c3rm7wkAeghu77pi5lJ7wSEiprh6rJ4LWIUEplG9gnzYMiPEoEL0Z
AncakWCtZd8lfFIahx9bhaX606gfiStg4Uhc9vDsgvxv2Gauki9JVlIxd8II5trK
Zede7ql58Dd3hZr+qPdvzR3D5+BYTbh72Cn7nZR56ZlRbB2AdB3y64QFbkVYMKcD
/35LFMLheTifGw+JsHN0mgReekbK1k6KG1z6iV37WyFWYH3WJL7yDnDetRLvVx5w
dZh9wTSS/qWTU7Teril1tpAqiQD7f18x2UCouVJK+XBLVP6CJrvy3lgkgFs/SsFz
OKY8MzWk4J/Ot5y/iB6aMZXopq7Q733mGg0o71DAYVyXAkeRt+DK8fFYFOGAnUdD
HTUlxtHfIyTVkEj5YeV47vor7d5R9PSaYdTk8L3XeAz9sw2EvpquY7DtCQpr2944
xAQ5nqF0bWtnAsnrqwoJw2D1y4JSDzkVIMpan6CGX6uwitreNZjiqViao5WvR0cd
kZYKzdAvJO5a1fK6GAU2bgHnSXmpEVtFs3f1uPDkjWYR6zrLxC2N+QJ8s2WenOmO
nycbFieqR/DiQBA+K6HZKKjknMkz2gwD5ppexBu1MaaUKAIJSKAUkCNvxfQTdkTd
sytLG3DyFLaRJISAM0g3fo7wIr69fXzu3BYAJ5U0axyqD0+6Ax82Z6rbcxVQsHiU
zwPpAUNajFvhrB4l0AzeWNXRqv+8Qa3pU2AOObUM9muy00uh/9XbwbTVdl8qMGuy
ts+0xA0ts3tuzIAytH617Lqe5hgWx84AzsroOFuxRAE8xLok59t7InabBCqa3ILi
tCrnKmqHJ23CbgOpiMHdyUbhh+yWFdbhKGxLtTfLjcJXwMViopGHV9W5LztX9o5O
npFyb8rqTnDMHH8FZYK5OXERPz8xXBxa1BQspW/SilQQi6ssHc1ht7K4ud+IiVX6
hnLjI08Qu509jAlu29eXzBLMVUSP1xodoAbQeVi4gu9l4VVaq7UW9QgHlDBoRbNN
sqd9daqFK/s0ItRN5BT5qU9q4nbbBEpvwlZ1NQpbRZ/fXzUwV2rcDNbgQ/HGhPYc
KUQ6QwIwRIj+/naxd2C9utfsmCml1sSQTXpf93DCiYr1YgionUBlOkmm9rtcU+xd
KrHVz8iw4Ib9DW0SjYVHTHrRIjXwwMx8jKgFtT6lUmbPv8uzMvTeFnUL29vqjoz8
urKwncVgWS1w1+/KRhUPwS7UPNt4SPjYyjbikBPZH/6uNFd2EwQEghcbIdv4Bzu5
n8+AZbh8JUtNogPSTqDtvViuD7T2vDvSb9QC0qS+5shkLK5iZvAXdfXyNyDuhIXq
2LRF6ggpG47bUESyxxCZtyXazjiqkxeYuWBZahWCBq8UnmzEPk0Sd67iBpyV2qcJ
lI2GJ/bLbrUPIQpewtfH/4u+Gkgl7Gw3ObFHmg8mVSLDakFMjn1gloLTJ+jiqdPG
EjlYbPD4Qh41s5cWd8sxzOdGz/rg41tq3tPxxSLV3GiRfYKV6bUlxh1j3TxEaZbl
rV1R7krJ9M8LV9QMpi2oTIntbw5g3g2W78vQhRbfM/vL3WgpmTWlnYKsfgyyz+hZ
Vdkm7EE7oA69jjMVCEyLUu+hUm6pbkHq/7cg4JV+kSiRi7TbLMKVH9bpwRv332Vu
9ITdUbvz++OPI/hxR5+ttIrSbt568ORJbd/WlXU55UjoHqkOs6IRINCQ0LFWqCWP
R60lZmLP1/hEILxId04qHbn6yI3E4RtornCiwXG1SU1DTi9eWaM0R93qig+INIl8
xrBUUyEYYs4iq9mIH13qwS8Xfjn8gXDrYHu31kDGr4BeySkPtbkeJepo3ubFy/NE
tJHgE/IqKzJalTwtXIxdvbdYu3YxweZfT/ImCyTsdv/r6cuqWFEavzXhrL+2pprt
sfUG6A3fLlctg02OWQ4aQXgvVYI/RsRZUgUFgvSSuLMmWiGrqkk2QrhT/XrxsItj
QLPRgWsR4zQTdZZSUvFrXu06CMz2IrCIEGFa0Eb+tdxgsa8FNzxGHcw6+Tw9Ite4
tNctqt0h2LNX/alrQl23h+d39Hzk4DeBz2RdbgC1J0HvPJVq3nSP/jrylVYTTCW+
di5LeK6U865Dy8vPxYu06ObKVxa0Z/zkU7chH+0aApGZBVJF9LRtyKm/TSjzuNZc
N91lqwKgwdNnPMerjarfP4TurP2jEVvcZ51Eehjae1ePjk3h/ZtS56ik6zcACZ0O
mD9fY2cQBHdb8tGZ030WcZ8OPNWFoeDsIvV1psHGdII7Eaf9Du4cjESE8gUKAGJt
j6Np6OF6J3wpavteroU2UlIaUcWrlunwKqIEDnl+khgvA9h4qfe2JLm7SNkPObuz
U75k3o5w4GFHeLPyg7gCGeHmDdTvpkv1ZMb4c8n6M6Z3GEoyqdo6EAyZX+agUzuE
5QYKIhAh+tOZz4Dn3ZtbOfIUg05JF+U+9zszgN6w0ORLIXJ3zLOot5Kz6T7DysyG
DfQZMv8jDTrURuO9mXEzfVg0y8oES3oKcGQmI9UU9rujCsQG/yKUqfY6wk+QORVO
kHuZthRXAkUBHHWWJINtsDLWa9vev7sNX5+mt9AaAnzq4HQXZRFP7rbVTzAK7pEw
uaIh7aYEqUs2KcCwmbpHPI/gDrk1kKGWg+t8GhCusAOqU9TFvcHhoCEOwMXRcj/V
4gZcr8mHMIJG6x/gLj5MWINhRThwW+cHcAxD2i/tMl2BvixDjDxvVBPRNYEKMe5b
X2NLfI5zc7pZFAyEmP++NHXOalO0IQu6UBp0bVxzzbSMCshERhYH79intl3WzINq
zPulMODEtEFP7lxS5H50uvE9CcBYJrFRDJE3x7DJ+NGy0Dg7WRfvFPf8aIzXode5
5QvrhyyS4t2fjm+M96l2tEXhFAN++2EXkd8BSsakOaCN7IeC74g/pxpDTehIm1iG
afqP85lInooOYSOsC2hN+p33FrW3YdwpkyyLjDS2L8U5JoLND39XtM5XeEMnKJKn
uUFfqSzbnsAAs1aNAwzl5jTIq0GY8P4vLIRHt9KzK6b/6VeVZK8BHc5PPRpJpM2e
SKyzUul6ken8w8qHclOaeZyuzco+TLFuOU/BZRR500MiY2D/FSEUDaCykv3vSxmi
SwE1iZy/qoTsDZ6PjT4OL+6/6KhBNlrDRcomJfkoD2nZYneOrqb/FNUDx44ed7VC
Q+USDuMFqSc1m5iQUA8qnsEHeJy2iR8Eg3VcE8p4yft0cKyY0HRQAxzPBMROHJzh
aFsX8nW7akZE0FkLfGdcVO3c86KmsHTuYoHm9uQ5QGixygLZT/eum51RK9YscFCJ
et7I6hBXxo6p1+YtZyKt0IqxGiCt6lbJt1bb9194ovmea1O42x6/j8L7qoQJCC8c
unuNwD2ATirO7crofim5TblrrIg2oXoEslgTiWjagxyTr8nHmqNO+v4ckdDzLB+X
fQkZbbvb2ANmwu4X7VfPu7YINXs4qiNFARbi0X7C4CRUVwthHUhnKCjc9QbhbQav
gJ4JrkTDdtZ5OYIX4M1OzjKXd9uUZEiDxjjvzFLrtgUir+7gaCXHnfEbuoq+LPGa
Ic1Ol9S1MQ37MJ3j6dbFfqeGF4bI0CBNyMR/xVAY4OkjL/JR9ByKl3mBqvpX/KcP
Pn1t4t6FMCC5u7wUWmDHRObGHj6WGgPW2HGgSuiQL+xdP2wXwknN+ZVojHSyLglO
LGjN4vexmMQAl5OmKb6axUycfYSN/+MjYLlQdXgVpiopjGNHPTSpPYO4rAljUpY2
smIXiEetgQS3RwPbYrtDqLfX2j5eCb/6TBK7nByFpvrbSswVnZNeDWXRMNLgLipY
+ZPH3HqSghRy4y6Be+k4tJ18xgpoSo8e+/QwlsR+L+O3A8Ylt24L7WFxjGBikVAl
cCNW4+Phh9BHjP0A2FMKxKivWRyI2wqIQU49MFNGsKKV2RQoxEKyMdVsL41Mv1ry
mGzYx1lz4h4IvEx8tveHVfirMMspOT2R9NrDnJT8ZY0WssvaS0mdGDp8nsfqZxKg
kkm7CRHHPqK3SV4M12zYEjbjDrIFHzcCPCAtAUWdMwavXTWSkLiTl4iMFaP/iwrS
Ah5XbKjEO/wgQvFBrOunYNyfEcidpmeQqN5+U5MDvkqtcNSThf6nl3i7kXBWNsi2
h3sBsz/6kazWuy3wXOaBGnrP15dlllhv21dj2mNAfxS2OfcZHSW0K8n7N4EQkxnC
4BjbfFDN86is7nlWk5OMNfkFb2C1/N/Yg/guL5Veazs4T+ymrePSpkJIQXfrMmbz
biDzL7B/TpZqUX5XkjedGUHzUwJErgSf65Oh6SOmhPickm+jfgcdd8FRzueW93tx
f2rJuWDHwnGzs6Qja67YsPf6gR2PM3RNJ33hJG5Ceg2jFP3K9sDuS7I7M7JIkEOC
Fh7tBurqR2sXPP5T05UMdjdXH9Pf2Q8Zc+tmNVjLgE0FdjDwbfIt3uJCY73MGmgh
26tfNfE3lf/iUPvxXiR+Sff10pZZApyZKVPFldlqh8Qo/9hV0mpGEhX2Qz+h49rU
w0MpF8fFwhmwQ5z9r4rO9zzkNMia7ecSqFH4IndAVkjFgwdR1QnhKhg+coveBEFz
qiF+24lFYButothHr9mF3+KKwPNdA0Qvoh91Q7vT9r+ARo8H2C0R58v+8xPeqvEJ
9dG7Jhe8j9eemhOW3vg+GcE1jQo/b8XyQZqYaWl9tgI8cTG97vGN+QkmYw9P2nhZ
3E4Zw499/ABjTOH1I0dw5Aqnss3TphsjqfADPYRTR3vdD8DvyZqc1uNewVUEzkAl
A6qEL+U8TlblnkkrVuN9GaKdFX2TnHFUzhFejMHozpmcbgwP92trlbjiu2QzOvjv
7lgvTYXXo6xtJVH6rZ4YlWwbSzJIrCuK1HKtNU2DQzqOE2w9ZgT3SKKe/dO4Ki+P
TTMmu0T5fY8Li00EPUEKo0ao7hKFuiLJqrTT4Sxg7UZNA7BWQocFBYa+RZUP8roW
6knhcZKDFcJtr1JkkviHECWkAhkxq8wNvcCAET0JPPjkFjahlazO8RH8KIrctH1r
DIwdUlRj8apDaEDxIP1u+U+RnJ/aMPN0/WJWakB0fgyY8GARObtyUjm/a6J6/A/5
U9LeWxK6/Y+fyYKgLexqKjNKlsZLI5Rvz3AquvBSLbaj51gLgrWiqswLM5OkeXTC
uH53VwYaG3fuw6cWmTW6Wmniarmfw5XBOSztLxbGpWbXZYAzJxnB9zT+H2ZjYMIr
jZe2MYhgRb7AsPG3NNMUeAC+JbXspEKee+oyOgnMl+eLCBiLcfS0aA0GP8kp5mqE
pJ/IHF497Y9MneMQZCDtrzn0JS7e20OVnVgo9itzjESJXZI4IRelPtYOcjU5tRcb
CUwsnqjdQDseblftgiLyfIM7ltHd/Qj5lBnWFAHwxzHVRuM4c+0FIwcuWIc8+2GZ
SvlczGkygIzSDoUKUtnHPhFKn1itxakvbpDV3N35XjujR02xynOqzevDuRrvuHHv
QIW8BOBMshP9/iy1AJqGj97mTAEtbKnxgz9+wX0GJyiL4E0jbAVQqssPKywmq7XO
gFt6JkphTKyGNFFzM6mO0SOUCRYXPMyRInM56+3ugZZ0p0TeJi53tye+fPcJS8KF
YNM+dP+Iygm0p2lko66KH6/33MH5JrmgNIvPQk2JYZWIZMEqhAPvDegAH/Bdxctb
HayV//TcaKNL59SO7CtbfPphyghx9QfDO82hEJurp107vWq6Rz3oGF2X/z6puxJt
WTn/Vpl6SuT/uQht7hWNNouEKqkibvl39aSTjZSIdlys/FDeN9ySsZBZkBA8QL8w
dvgFMh/kLM3IXH6/4Rss5k98orGPJz17G0hbMy3EABtIfGNLbkbxicHds9/Et0St
aQFcaSNItd3CRYY2SXi5WCt1qNVvLc1dnFlNGw37XWOgFeH8g5VgsgIMQjr/Q657
Zh3g5ca2/6otdfUV07i2sc4GL81cERF5q62kO2FN24SV4k59MDikS6jSsRsLNqFt
VCN4jBHI6UMbZq9LTQ+pM7jZudfzO7CaeSvpo1HI9zrNICB8WOgFvI7z4v7NnQCn
eOLcP3qlnshFBrQFq/y7TsMb+07duO5rLD6+ipJf1qTl6RGi1wCjft/T59ee6fI2
8g8XjtaEI9vOB+MlSBZ2oPRWcb2tsB1TPnL0gaZUDtBSrPs52N9NOJ0o05QCzpzw
eJsH291Y+8Y7EiB6mDR0Yo93uO+8JbNcbPc/ubOK3MlhQksVg3kgNwyRt5AZOv/c
TwsNjwtza+fx6TJexIwB9ltru0hTi5df3Od1l6YShL2zQ9lRYH0sh3HaLsVkJdqZ
rZVvM+PtcweNgQETDMFTl/LtCgM8/swqraIJ+S354QaBJ9/kT4T+LJR2RmhRnqH4
W6rETaseeruAWiKiQcxm1bfRhsvekVoxnd5AlfrMFe2QLxqr3MRA93fOcHz3VVkj
HCEPMhDjGTdONENuUphdoJQIqmRDCkbBbf6oQOBihBSoZ4azCvKKBwUsRfakmvGb
o+jMzA6vZJrn8HKf+rm+Vo7uk97sxFeupgOn8eAzNqiMUsw26xpfhWAjWOIgLW2r
+3VFke6HsqgNvToTz1LD3redeUxtAl09X63LiTeb9IllDfekBAVsKdmo1sm6aLHt
PRhUiVjpw1FdSQy1iqWWYIQmaoUrm7qWWvggGUsxMYvG+ncF9oJuNYZu3oulo/JH
0a+Tk/auFk1ZbQSYUfwbo9RzMYk+r4xfHTlW2UApWr51c+39n0qPYVI2e9x7EdcW
fcTsosm+/hnVVjt6YQBmVV+I+YmJ5bamqB9Gyz3wP86xzmlredYrD0UGUipfwtCv
KPxb10uOk8IWDRoQlVB+iASUj5sQFleQpP4WhzeYhjuvcKEeCfWjolGyLS8S4mRx
lDFZzd3WHwfccm3RSYqsEoJ9AW9EUsg3WXvN2P7QlLQiDYoi7lvLA5HCbBrRL6ws
MlMYYO2dBmszgLmoECHUGx9xqQAT+tYX/k1FdFvCG4vQCW5ct0bIihf5jdQC1gFA
ekG6YkKdGDVQg9q2jNWwUC38Otgx79H5S/pL3Bce4SeJs7gjO2sPkmN8yhG1edVQ
t09dNz7f7eA8WL9Cnh6CuW+2byboq7jTOyzGXANc+t5pXZVcglUf9ZMx20uFaZo3
v7dvIKrYLLbp3GBkkEYu1gCxsSdQv8SWQTUP7yJzX7sqVm1cFz13CO4E7xqTW0cg
dN224GvRXfKKbIS6imo79h9qwbjaltjZFk5/yxYMPaPmF7PtsSM3JTDQswz+gZJc
ZEs7mdkVsHYKckSgz3M+OmHEvroJtN/hJu6x9ZkclAf1Px0CL3Kj01+5FvPf7Uza
wrQdugd/+GbkFpdWDjsa8vH05eXu+RB8OqwmEEe1axJD3sy6KsB+JejSP39dTMsw
4OIx3ODZyKAqdvNZ8dk6iF90Xk/nCv13IvLzOgKVCdQIUUgQXpCPW9tjM9V69mIw
FrbIFwtGsQKQaAfmhx4Ty2IRvxXXk0ovFOM8k1Yki7ap6daG+sWnbwespmAm45AC
x8YpevuTfM6C3hpRezTA3Vyf98/luYux95bSPSMVbp4lVpHos/gsb19ngWe3uN6o
HDLAgJyxaWG0Mp+6nrPI9MP/ViG4staAvDLUPLgDBJA4PxH7jYLsgiXcQtBnPnLF
F2HmmqTHT61d3GWCVIHzXm3uQGb4H4LwOozE9l9XXlYYY568n7xPt4E9uS4kKIiH
vWZ35nbLwRC8ItKrEHmo67im+cKiu8iSCwp0jnv7EslgEpHqma/JJZbQcNoNfANk
40XHtjaGsb+lyDnzpW5fGyKfdBB3An5q6xBLl2A2wEgKtctOKprbCV1q0W18s/gR
3RRVHgABt4VmH60wmyFqUUnrR8AbreoePz5V9IP6Q2RjlSvvlWcuKn/kO5zN3AaR
mQ+/yfPNCgXDgvWQaTJr3V/b8hEnnPF9+zu69RrokvRUp6OCxnJPpyyCMsT7u7JJ
541Ied4/KeoKZuvwoiR6/b4KrmSpIGLcm6cxhpgz7bP8+h99uh5QsZ9L2XyrH87Q
j09A7oWNMisKCLkmAnlmlyA9CkH6c3+0Jx2+N4OqUOMVtnHXq/ywp+PAiok7qVEY
91UVkZYQ3r5DcZ7uQAe8MEnOJi2++48oBU38ZBJpGllX82m1ZY2+PZW5Et1dNByM
JfI1vKa3xmeDk/dRJ+zHRdrFJnxbqqu79rNDB1mEh+TndIBn+q41V6FiHqERJtbJ
M2Dz1vgupk2XLjyJrhtBwE2PpbpGAC49gFdXkbocU1bDQ2kPxiiY8D4PtFiirlba
8aNT0AuIu2M8C+RJN7OaMNpFyzTC1zQh4BgOMJxCSVOTzM/cqsUmQjPNunlpBTC8
UgqWVUL178Acs0bokEVgGR4zCQ0L1Olv0LxB8pDxlmLG7TERAcMmcNx264uT4rAO
GJP4M3ixv5TEBhwuKcozYT9LC9Y9OripAUP81aBN9iJN+McN3YsdRla1wqlGVjns
jOgD2cHrXbP3BzrGaaxhKApCieTLc2NElVtAlak2X5L+VNm/Xw+CIoS8kSZhTg5b
IazYag5WhRuY5MHarlnuZ9Bj7myRNqps1V89DVOdv1f16oLG49tM+pc+Fd1Pi493
PNgWRhuhAtXIB5yNovhEbzInJ8qSKjB9uDn+gA9tTjSbUon/47oYIckv752UZcys
fKHxlmPdXS9TaQmf52RoiHfYYr129SZurbBectHGkggzTtOGOY+aanAddY8bfV7C
njUphZm7QbfCpXfnG0t2vgL7DMu7zAMDMe5I8zE9a9OG4jxmXj+ExUH6aTBSsQy6
5rN/fS3qTUXrIlBUHZrwq1pk9fmClspWKvJuljPekbgXhDFCXkhajPI1caNh659T
JSiBWLhMI0DpDSMglL3cqpNiurgjWZtngPtAf7ODEhmyLizmD637jGFgu3qNI7oK
SsJnDbT/Co+5URlkoaHwlH8P2eBb1fJcwV28kXMrrqXBUZ9x6d4p30X9IidqssXT
MEGf7mtRl5xJC/8mr8ZMF++iRn5+dzNbgysVvewPlZ9a+nKS5FZSu1B+I5NaAC/e
3KmQXyI5MgGCN/4l/bJVCjaPZE/zLvsjGngPCAtjMyAJ89tmzQrNVjps3s+C5Ray
TbEnX70X3bO8xUVWkdEGtz89nrKUwIc/a5yveouz9dX1++YB6G6MmawY8PBJlh52
osMwQzJyJ2NJyc0FbrFjDpyXaWhllRi6Kef8HMZHrHzu9fyW0hbz0zjVON4TsAFg
m+xXs8Mx8iV7UAD4fS+v+atQ8jAHSJOQtKpoq81PoyaemlDhAdKOhvRE4qiG607g
oBokcai8WjoW+M9YUxfDjjY0KSrwMMZjUi32gnM5tEFmNX6pX271vMcC1XeEHrjR
RNOibpnVLoLro/OT45VwF7no+VlqxdBZrbTDsDRWPs+bz9xgKREGT9a2pQPha/bl
01hvGSJSkxUFN3H067XHBDD+IIH9mNc9TPlGOHHk0YdqZb0s0hmm+seeU7SuYDvp
lsZw/ycethadOheaudwjIMhu1kM94yxMWyhE2eK/NHpLIRSggdkvTqzJnIJJAAes
Z2Sj7T2ElhMUYm5KWW+2+JhnHETr9EgEafpTnrp5mxOiRoWtnH6DgIm3AjLgaWjm
44Ps1iMvv++Qa6ZrXU2lSM3yCqPZnrZtsTzr3PadxCO8QsFmtGGxpqT6JVrlvc78
c4FK3Sdgd5Nsmi1dEe6H+liRwgTbRq9pHBarMxiLlKo8PYxrPG/D32ALTrr1le/u
yuRG71Tr8FgWLRvx+daJJQRWSPPy2bJRWmzj+eOdzJJwahvCNwCTYNVB3sfltcSB
d2/0TfpvJNA+vCmomVHxpHlQlf0mQq03fxVxqjHL3iokt626rAhbJRgZQBW3XJ1o
AP1kzeZPLwFlRgvzAU9r0gJqtJTBibqMualOZ4bF9VxaeWkZcA6+jiLwSCVw+KLp
eMciruDSNOM6W86u7ACuuP1xybB3pGVexRzlweCVQj3yaOe8l94jfobvx4fdqQY0
31w9zbkfVBKf2XlGUjOWR48lG6E13C9pPRqYN11ZGME8ic4zlBrt8lRS+BSIAFeF
pJI5aPscfC0eZYIBCrJ8oC+BFuCwQgGrXsNzGTGxtq82k4v+mykdVV+wOkB/bmGi
TkbtzlBThJDqxjdQNv8DAHkqWpu+7rpAqLwDb6rH9Ny7hqcbYCE7PJlP+vfqy0ib
xFV0K12+1IWZl1woPAaUMUFPEn/8vM93xtn2SCBNa8JV5JlPbAiTIgh4CvzU77Oe
arRHeVrUALRyQBTknFdTXd/HkyOrYpp9qbOAn+8dbIhSue1aUApvtTN5x18y0BVT
D17LMR2bckPK1ZETIAH05Pm6C7FO7MEA3tnSHRa9YJR3p057Q9vjLJ2wMpAkGbXA
QtIju53t5umNshw+o/PoGKJFBXxw9SeYFeNZFHdGQBWC1gUWR30GyPteHlIbxMAk
6zDaBsjdNYKFJshz44lEFgJH1FXnghcAM1S6VJpMEl3za4SsXs0vu/JYBQW//5ew
P9uVyCIWz+5a5YcUGkv5KeDasLRpcmTqnpLhiGJCQ/ByMR5tG1vwUDQkpgDEwDuc
KV06jwQdD69Kad/N+JSgNcczzypKwPGKavU1UKFgpuQkXLAeklhcTe8zwuAKWQbI
dm+t6OJ5H4awOTo+uYGIkLEHizPct8JgcGMg+ZEt9lnLZ6zvgp2J87zcXk6AQNc8
h4TapMuVwXw/mBG6oCvRR0h7EiP3mhZrxA2TO4Em5Vg/HK72odL4cCzXpWvhJxx2
5gzVVL3aRXJLFrJUolJcVLcJGjSFekC2ewDncGkbfuMlbUhpCXfDK6hugGBtx0fz
mfIUbG+RxlLxP0pozNFIkgQqarFQqRqr2md3Y3/JJWhpkxzAgtAL3htqZCkrnA7n
KS/49os5C7TGshCAhO0dbb2lxwDDoVjGR1UduHiED0/b9lx3KCVmpTRY1P9f3Exn
I1+a7jUrmJvxaa4kSpvOf49HBxPw6PRjQ41Wnl9kOO+1HhWezovzUYxI8fhGQRU5
ATKarLH6sbahiKwqxP2/wOQ+UVpmH/8DzcLEZUmYdqsMRrIyzWoJKA2WQpVa2Am4
yFh58g3KCNTwhatsFTnEkAonXB7TV0dQuCyBNP6lwUDxKMUhBR7Boz3YGSGaEqnA
8MWth7JueF4xVyBiGwrFrXh0hq2l2gjVQQV2KwwG6P8NvWVwR3YdDethI+C/nt5K
6/e1cqE71tvCSWM6kGtLD7t1z2IeYD8g57GmSxHT8Q0uyvt13S2WVTQ3LJ2ncKpa
AVDm3PdVRHW0p7cUicx7fBNI/Fm774lklMwgHksar2CmFIbQUUzg3WhbaHrpYZdN
2hnAX3rw4Yb/kpVnbMq0pHhuc/04ugO7N+tKiAnKnW5XluLgiKUb6fuj9L0zgbFX
biVPj+PHCC89XmyO3sT1jxVjC22Sb2uJ8ynDBvz3jB0aPxyT2fLVqakmuGDi38ct
CTqEOUGiXSMhd0yugC0GOmxPXaL2s48axi7T+NKkqggUC4f9X3LHlMoUrrrkPy2a
oAjIKAN/m6Vfbf2o6DQPr81FdT0dJRMReb0D66zJ7jzDnujI0cXdO/pmfNJr4VV1
e6QQ4WpHELBCRexVL3aO5EEyn6tyF6BSRKRV2yu9Y6/opxuoJ22PI5d+8wC/b5qL
qnxXiWDVsG+xEpBscwQmDeoFpQ8jAuiBGbNKf32p8R+VkMBGYKtadN3BUPSVyW9j
LygVQ2JXpfR4wc+GBjvXcalS8t/LsyaXj8trU0VWF2pmyAGxJaOKavHV4hXZ2XN9
pHeHfyBbtX7WX3+kzU3RMZg7x24SPuqaYd53Baugq2XS23jyJxneJrTY/EZVJMgL
WJ8q6q1jtoQtSR33R7tGgMgma+fljL0/KGztGP7NMvzRbPtrzDYkMHM785URCx0Z
G12/dmoQh627jEH2yuZ7ASXCIJxdu+Tdl4neEFMhE9Rfy4BAmn8Mv1emjUeMXybs
c/y0ATnARSWu8Ib22Keh1kkoMY0ZyMkO0OSNNUvZKuvdNSnhXOoN4aQvWVs281ac
7pltb7HP+vrYyilIE7OWlwbJqXto5GFJFJlJOc/l6USJjavJxQMF0w133RnfVI+i
16RPMWjuujo+QfSO7HPoU9EMIWEJi18CiP5LT9qbqUcj9Ksm73ALkt5l6U75f1ws
CKQYQi6k3AYd0JwVN8E6VSZu/oH2f6VD3mb0Xobqvmvszpwc1qaQ99SYiAXkla9y
1T4REXn89M2mwi7EuH4YUb7tHAKjmRJV7Kh6oIzrzEoz66Rxro7cqAh7/m0vwBZF
foUe/d9nzy2yLa2ia2L9jpFU6c7CK6QvFf0mZULzkzZ3VsXvZsZT6aZKZz5E0IQH
6+tggQ0Kn01a0bLkgctOVRdyE9ozS19xEvcvdH+Ol4bJ6Ri9qBMQrrs8kM3ilImP
dSDG8sgslkDGojD4XDExV35KK43FqarF+DZrk1BmK826uRjPo71h2jZU5HzQ5QIm
TyEQ/clIhhoKwy5lZY8hCQdGmCagcIalZTBidylyv7CK6YYSyjwkRdBqoY3Xk+LW
hR6sx1bWERrZDDV4LND1uyNcDptPBtiXvZi3Ram0WdKsn0+3kUKVLQG0cpi81hfU
xibDtpyDKctjYqdDMx24cVKNQvKoeKNzU/06ATWbMAf/I9WIi7s1kf6UlpzsuA3n
wLPVrxFTIxIVp+N5Hpa38TgelfprN1JIrb7tsM/BwERdny937P+n0Sh0HZys15R9
/ScTd0ymsfzIQneGhdduDtKeca215lJb+eU1cwSXp8IRgeuWJ7s315Q3N/FkHiQm
90habQ2AhRtBTNOFyQYkoZt8LADR+R27Fxa9TzI4+uWpcJT8UdpN5eJ7fVOrDtH+
XwItQNWUQQ2uYWI0xiDlEBHGskjFp6AZXCt0Yrxlc9j3gtXEMqhV+vqNl4MMRS13
woaViu8qiiKgcCynunYJapJ1sHpCSP7zLfqzFPrUEhh07v48G4YAX0DIY/775IT5
O8E983brDho8081DJ/uzq+Jtt/CCz3kpq12OdHRk72BKW4nKcM3xXMxEru9aOnFj
+ByTluRHDEYCPWHEhU0d0YvA/6SeMRNwudLxfx2ZsKcs0IpCBR6vwHis2YBm2Bd8
RYzmwqbvw1I/7zuTB6Q2Hlwyw5W7KuQLvGqsn8+InkAB++1vQyVgHS/rzWRXDHwL
TZ2y57WRJXpywPz839qnvTROGSsPOAE6RiD+0ZQ00Z4ToRpqSS2TDxZV9KG5MSTI
zPD2a9ILH7nYOoXpbYmJad/HPANpBvKS/5Y3wmg4SOCa5Hj/SV0kNpu72H4CAKpO
YhXRU7B1PxMvlcO+CuYtTe8ZjAFLqTigTbD1O3uYxuB5RnxoiLH2OJvlrMQbwhk8
KfcmGsIAaZ4rq7L0A7Jo9QMD1vskiEu2y02+ycCAcRp3tdBJYjEf/SLfqr8h1vt5
4IwEzP6XqRtHKIUgTHe3nKWFs24sa6IrzkH/q/yMfXpJdzWAfc4+Uw6vQ6Gtwi0M
Rhde6rbQocR32kZ3SQJ6LRuw4GYdIeKcEEahmv8TYOlUeDRvDiNAYLkybm6VnLBR
wfFzihc/t4awGu8Gsn2TQuzZIFiYLj8mOvLwV5KwnUmkeRmK6sW8qlETf/Lq5MVq
xVsziCzpcH0EIReMQv8OkW+GtmYXvR0c104v83wg3JHPXodngCoDgIDX1a+iiXNd
8nmbGQrwuffdGawq3adoRSBB1hhA1OCcCT/9K85klc+opLC2btGf7V75Hlhj936B
NzgV/2eqjwHRQLW3IZNYWrMLp6X+whzfDkmQtU5sSds+IfFD2sAzHJS6JdQ6SU5E
KvFc2IqHTJv/VN6aH5hn4OJ8iVD3bJ6bufLdEN96xzoAEIVb+4/tM+chVWjMIO1P
B81fXKZ20VH31mmLLtECUdFSnK1QKPVQssunlTpOvi6nIB1vrgOH0a4H8e4Wgssl
lg37Qh/KvgUmg3rmW5TcaxEHWy3/6FeHWqKBuBmXrLDH0XXj41hcXeuK834GmYWF
IidE42VNEo41ZkYnUATFXF1q5OsXY17FHi7eIU7GMl2PIzJ8T0t3QM7n2hkcqrpY
4a9RZX4+4wCd7fcJq8tijfsmPLgZ1mKJAS3w00faghwY1956ygsP6ll0QhzXcfz/
ozGgGzFf4Ajgvo9i4khqociQN1tGVbgoVKET3RV1QMgS20srvTgxsHPXo+miAWVO
XLyydEEqsZ/WZR3uaAJkbx70VYctNcQknKBD+bCbQAE2LfS3zQcZaF+ryrR08bvJ
Cm8IN2Vr7ekkkNpa8jfKH025YyN/SrR57Oh9+RPc9ryny1ANg80q7XboR0jYs9bx
fIxjn6+FZkUChU30Y9W5+JlZGw1PfHOP7q9a9tVSBrd1YEXDf7nBntDRrOcF4K7L
aa90YG8qUENQtfcg/BVG9JygjYwxO8P8SXvPmjX3Rd3FbvUR/gCptYfe223mQmxa
ZkHkvVt4HmbGOYw0Vk90iQkxJAyKbGJKxqeeRjbpkknf/p1xXHXa1WjVCsJuPsg2
p21NY3vwMCXG9pkQIGjnrjZTunff9xdTOCxpA2Zk5xER5+thhMwmTMEL4SgOGeqb
++sN4xxIZbo8lJe3sd/F7TMUZpY15Brju2dFg7Zt9ygSzFVqAZYxyD8GoJAXnjR0
+pi0rEPOHAQ8IKlW9FmJPI+McNrGm+3nljkaTkzfd3TGNVNFTZSZCrHsHTpuUF/B
0jSjpBJ0FbkxHisI+BrdfHpc4niSYHhdL5Tsc8hfUOgliySpCLIixBC89m/K3K3U
N8ZHjFy/ZwpyP5oCXcoKNo/KVim3vrXl2tK4189vV3FiVgqOYFyUP+RgChZKA4P0
4ojST87YIyIoaYbO1+NqVN9mxYsmSWZ+q5FyQ206O2xgkud4m4EAUalpTR6VyKZ8
LUu0/zvoaESH6eG2fZXj6b0pDA3S+k7GaQ+hMAYnthMtJOrx9tT9dXtxBNohAX1i
mvOl7xFOrbaWuvRd4YtGt+9VHEOGGRRbVBg6q3LlSkhOPjW1yus3zTl5Mi2uI/ao
Td6xSRGYRUgL8VmYa0U7irITPGVRwrHWnE+yUSq3NsnvMpfuOp96KksCeFGfLOeD
cfHLfV3Ok1TAXnIxZfXvjCCkSW1GANQnlQ0VCEviTG4fyrQl2Rm32CQ+Sp9xoqLG
/S2Y3DaRFLXvfVVsAYvn0a/lAfaPafRnKR5smS0L3850aJD9DMDqMFpmShmkTkuC
fJTnDHXP/zprc5J1T7oiUJ3UEmvPsvAjRGc8rZEDIP/YSwr+fF21jVB1xTKr1ezL
xhkhG7qDYSgn2ApcI5dYPRc3VAdv0rob2/Dgz360XaP5dk+MJ/4C/OuLixsuT7Gh
1BiBK/l9UVVhYQf5PmHs50ZsvPF6Sa6fbAU9GudHnYp3yYuEnG779LQDesuenyBd
VXXS3aINqKRHj4+DdJQEqX+2gyPnlyImfMB9z47YpX5JIm8QXjaEXwRzXYtUP5Oc
2+dOXTSa+YGoW+9v08suM5Cy2KExXlJVRSSK73sKPnzuoruWQmyWGCFQLpHDax5r
gc+/b3jHLfhkUiPAHeZ+If6kp37wX2Uxzf0erZO1YIv4e02JSE/GWhq+7P6dtJ35
lquDMjLAeKH9OMlYkVdw5ZTmge4ChwznLfeZS0FXhenMNhc07d7wcsd0qOtpj+Uq
cRIlseAp4CT8fWfaQuVPQT9uRMAn4QMnb3/6JN1ojf01esw4ksv1ykl+NzQA/pdS
HWIzv5E9oap1KYgMY+7OMHgHGjldy0Ra5caqzHy1ed/2s7xO5WZmyd9ACO8YfbfE
e/Z9rQI3uTazJZLCKCffDNx0z0Sje+MYcpkQZztzgVvhMt9neDQ4WT4HKN1bLdXz
J3vMK6CIyDOK6eGD+Ael50Y+FJi1ppVkkhdL/K1lWfBzFuxhpbIsqGmuiUANbSTX
QiGL4COG0xuZXLfZjxKxn3f8MYcodWPOIY7tCw7o5r+Wi031en4lWuaJbg5GkOi1
9CD0QCiCZ/OebBWLo6zYa4ZqwUa6kPmE2xxo0sd+tbl84c2gN4t9PmdqRVoKOKRO
pnJaYOYdMOM0NBSwh8O0w2c9QUaGXxhahdNngoNb9qmwvIp0qkx+tHRR1PAhHAQy
TnObmyA7JrNKThiYVd/ngrKOpGSiXKD4CoMd1zf5MtYNsWk5QojfcogkDBEsyT6o
AbRq7XjTUCzBOWZBDxyGvrswrNLNmMs6jp0rYTy9vgZQoX7X0lb0Au8anva85Cai
dHKJDemE+b+uIOJkvkjHOYQ8hsrR2QIFjvXqMlfcAg6BCx5OfBHdtTKdt/KfVWsJ
DPY0BH7tois1YzMT2pcRokZMCvAgYs47crkM8BAE8uBcrkU2I93HnQsGbSHc3lDH
fsaZ4E4KvYHK5nRnJLof8yiXuu8LC2MjX1zIT1GY4MVH+GUKV3rSIX09rBEZ56oU
JE/QjNMqOr9bX27Nfj8EcPJi7obeXFHiAlXl89DVONZQ2exu1kwGMm2ebo84we/K
TbJJfNNKhaywUPbnJJBatk8fU36ONM3pWC7QcKhngkCPthjIH7XgJUPgLQt5AbGc
WM63C0rLpw/SjWDMa5jbxSgEvqs4mlozc2bqGfI6hsSgaRjFTcq+hh+91EGNLo6N
/O+4JOQDWoUrMDfJPI25YImIuj+0PYjmuygT9Pl/LNmkmkydSL37zI/34URd+xLq
yPi87FS+E0oCZgwsgJ5zszy4JzKAe/iayRmM3NN+kW+VXKmKAyclIdRcnWkJfFaA
EjP5wzI2rImMHyKiGoQmNquqIo+5roz5DNhPfmh6+zK+Po7qNv6O8rc88DQidYnb
71K4V8QIcBtIzrlRCGKR/Sn0QYhxfVCfKV/zwR4/QXTYKu4zTTqYiiE3wPpIQsO9
A4BteTeqJYNA/ZwwtWB6kJ55df2Iygq1tocszgU2ia5O3Ev5x2DQQTr0hY9uqZgg
4Y0BSxrIpXfOa/UN1PcMMfc9ieNBF+dnHsQPmJ1mQ3U4NtphBg6CGqpcFRDWepKA
S8R+b3iF/X0WUB7swwnfX6T8FJD0lE9SBTgEiia6IM5vtmf5rXBhrqar3bdeYxyA
GE1fU4f/L1Gm6ItxUWpyjZx7PJJP68Cnujwm+YYzK/usDt8B/kXYVeABd2r2xOd0
Fb1P7rsJfoH/kMYtia3PL54ABT12t/Nco8SwLhtDWW19EhuIP3jmOmCr4nsU+msx
jRGK4bAIbA06wxtZVG/TUC59hH3THWr0/6JeB+jsMcFr5hTN7s8oM8jkto8LOjOk
sBr4Fw+x+Ifo6BzvqQi1w9pIFVgQAT6qtmeCkxqAWHOi8JuxT1kabFIKfVlgG2Y6
KKxRNyY85xCQoq16NItsePEAp0xu7POu7GOF3H+saURRPLkVQ60M47afoLmQyyTx
fBvUzWiWFcceJmORHS6vygkebEtPPI9Iz7xmvTxizAwM0wQLvAksOtGFzsW5roVY
XWFN7aSxgWsnDNilVQ9O5j5Gv7iJVJVP54ie7xmP9IO/QiY138d5L84ZYbYXKfT3
ep5FhyArWenCVblOd3TF4i6vxv90lUVUPKhCiGOr34yXheUFKx9MvqoCbMyI+ajq
oI/1n1822eNFtNHbPQJDiI2mL0BO2mAqd5AVARgBSGKEp660TnVhJyB9/Xqm9LEX
N7l2A+BLF/cQbHVXAG0rnUPC/dJqYaM1qWbxzyE6TaqxcCP+a7fgRB5yc5fr1yHQ
LYRZ2FFR75ey+rxEfbSZUTSDCECChzCuhPghJx0I/MsKyPdhVbjberkp3Livoz0L
yVnVT7PDn4iKGNJgiuuulEVPQD/KgKW54Lhc2pddpv/PRLcnx0qeSgPx1H+KiJ9n
Aa10Fzcxh/hxTr0Qt6lSqt7I0NEmYETPPyHd8DUrN2rjaMd6XGKLLwH+EDwTincc
9p8KpEiPDKpHpr/qQ3MG50oloyxLQoyXEBhV8QW5zCU3hvGCrWDfmVrhv9mglnFT
bpDdK2ABVCdn8qwefDA0fX4hOpILqDTb9MXQIBEwJ/yAIk6X6JiLDpcPIItiTyvU
1KtMzhk2PAtafQkkYsM/tvFqIVWUSLYLuTzAUeaasglNqJqXEPx5wAXu+PwJ2g67
UZMLKS09IHbRZ+aO4UzYdn5yG6lnf0smJkdGL3d/VlKpffZ/+xgB1xJG/zZglO/x
kynt91ZPk7+ADE/6JbrloPmSNGwa/eCtFjBPWmq8fgi9t7J7UMEY2OCJF2ZBv10y
pnrKCjL+9eENMwmzcWM+8ZB6o/lmeX/mLmYeNdXDgxjQYI1ATgpgEp1/lbuglVlk
KbzUFVv7OEsl/DAD9LFkMLKqzo1eASFzm8oKdcq4iyagyMhuXNlP8HL5Ec7Nskba
n5qSqzzMR7kLkDumejwcOzk9J8MFnMiLufVdWEXBPjm4/pomp29/5wsdBXTsv9iY
vEHTE+Og9SdVNZdjqtfdPDM1hIG4lwS7iIHrPKtQmyAzq3oB++7PoGuAIFeVIoct
TYL47GNJftxGAkhqSs/kYHAi8Q2eaQ9ZR1RskeZ6pqu3HRaDsjTOQHHBgNv4HX0a
GED51pSJSXxeHmJsnWAh3G8wcANGqLYQU36ACSc7ilH5O67wPzgdgZAFybg71HjD
ey9bZj/JJT42TrpZuI7RsMfTnVdUuWxNTvscXTBEEAPYGmDCjP829cpfU/15zxaC
DI17NE74+SMabyB385ECDue2j1TTJb1UQGBtnQLHIlsAe4JnrwiOZbvm/Uy7WNnR
+2S2ebfrM/4s3fSy9gwke9okLiNC8zQmwz2n5y3F0p7q5afF9ojTqkWk6JfrwvKg
L+ef/zZek09j0UtwadxSJNM8cHdHv9Z0pLNdwxryuzHSWhyV6XH2ngEIjCv0/R5s
ke+pi+2pnzVaWVtvZXckSY3KzCKTScGOPFWWtMwewW1CF35FmPaN6XEF0LF+ji1n
uaevyFd+ybGFGzrlmMKVuTDxUyc/6fQ9rk5cdBd9Nt0M5nQif/bziyOjoOnK1CcK
fTCayLMeDrBkdNRlQbBGxS2r16T9GPmr+7A1ubT3Q9GPAjH1IyoIbikNyEFfvpkd
PEN1hCqdTU8bvWCYCkqGMlzoTWERkeQOn3KhTU4Z3m+v8ODCwgZ0H92ocNSytQN3
mXjuxg9QVsG7DDKgJZwGjyXB85OiMbIf5l1LLzbg8sx/DiniD2OnhNvW+RB2EJH8
18vqm8mjvquEdd04sFd13hPYkhyKqf3/GlmY1Way7vEucLUVa2si07oTUfUWccG8
K9H+O/vIPexPGPqE6WR5KiTQMQSRdyfW9tv1D3edBVpVfevlvxJVJe2PpgMQNqrH
E78MTvZw1mdhqIDM9s3CnuTmasY/2qK9RforfISEnpFnrsJbc/sNQnCM8OpLncH4
Z2KLxCYBtaR6d5OGHhu6Kxog8taYD0tmyz1T8ICfDZ1gqvuca+8wdAOxcwXej1IZ
XbgqS0yT53FuMD/CW1NSinII6HM39QpX7YB8kgsl0ZZ5i8W4DBpTMqFYGGnuOn6f
S2sI0s56AvC6T3kyn7WJ6YvymVfDgbKccrnafD1XMFKqmvRxhnpAh3m7UNNQtH+M
7XHMybemG71ob0hULC7sQV952fLN75peV+NnIbRkj6hTrRZ35rYBdS/zEFRQok6p
NwnJxs4fQt/+7ZdtuW3aNYbo8IS9jSphFdlwI/1xPaF7CVuv8U5Q+5ROmURWy5Og
OOyFvyX0/YHfmc98FfgTl+O+ep3FU4n6O0lDAmjWMg6QcFD87ksGUdxlE5ZwyBun
mJeSXZ5xF/VUuhEiJE9wt43vqtDPuU1ief/PJNlJnRMC1/e7IsTZ+rx2rLILa2Qq
3wkmx+Kq5zEH4B5BH+hIKiyq8HeDnKCl6TIAuXF0gDHt++kbbopwD8U7ghYXJjAC
V29r54otLqtSUHx9Cs20YslkVxDmKaahNZSwJ58syB6TAtmrlxl2jsOO8tAGZeWv
dZJPAYtdX6ggwkSCxPTZcBxsKSGCaMJT6eVCjkOTrtIwWGAM86a7+cZmSP/yI2OV
SiYRUgRunPewBcrab3LtGO1CcNg/EJdBnC3m3b+gWiEXSuFvAH3W++/FHUoKy3Y9
B9RCaEc7jKnA8eNIX/SCYtBxGQABzjA/vn9mLTsKuqvhovnWMpfCu1jwEAwetdPX
qz3WZe0RfjC+GkTzrWaaK3EnO4ZAeHYjMioxMPAt8mtJ/0CuAwjSlUMiLgVD900W
dsXa652NboWd4hiObyFtAmJxXFgplxVrN2sxLTsflUoBCBONOzGM9aw5GNL2dDCW
ydORAwl3ONwJLgmjsTmQL/xiNpAAj+TRfvPps3KrltcukQCPzqfbX5/LF5IT+Olj
5amQ4B4syKhSdPB9tvS5q9FqqPSo5B/udLXPssYw0Yq5RkBAcP6CmGAh5LDvJf8V
wTQRiYG6Oqiwx+4V+YpASn5pTZoZt43B3Bx0Apc44QWnhnqhggHDV5E5N9qLzH2J
cy8RkEpLuPsDajBvqyEvxgpExsuCgM1XEX/A3hOU7GBlZyhgAyNsKXOWYCEeM7NP
ba2/Vu2EEXZZ5X0+UzoeteZvMcq8uCCyA0pqYU2Ywv76sgUAGf8efk85RwfIIYNz
9HIB03BuwqyWXDoD25J05tnaKveys3HyUfw33csneTerjVh2vYC3F2v6hmvvxldZ
7Y9p76FMUE9MyVEd6mWQFO3mdjE3HCbTtzeijy2f+QyRwzbEAv454dm+6lCcmbnY
fp4Y9Egr7+Pb8lR2hc0g7MFnEoy/3NSnBjCm2i4ecujguVIoZOKekkjiY8JFJdrL
oqOjEb6LyZGJMFEHJvJ/2xCuS0Gi6Glfh0AL1oxz3dT36wUF4arWWiiOoE0mQxTh
/km0gVIAhhx/FawjAgLF0y90P+StqxWPL+JjsmkHioSeQ40enJy7pMLcyjesE7LH
JiMqhmYiK0z5ApAae2CaEk4KgwMyhjHoERZfz+iDPqY+4r6u50Drgf0WYxaW0xvz
+yOPqqwwGeAfDoW9Z+PrrbhBW85gzvyHTDtGrQ6j8FDdHSYWeaK7ZRDAdVXYr/cA
TOiC+vSvGUc1Xt6GYCcT9QMNy3E/U5+LAwirKuV955/+zpsMnpONIwzmm4aTX6YQ
E0seMDKVs+o8ui9XE1uNCWYTJlAaFgdJ5/3bCyjOJrxvxSCwfckAZzGos3XoNfC6
z1oXfPgSTXVgSuQ2DOl9tBKs1yM6KodVbm5WBRosc8Ka4XytYAHOqKUfCWtTgRnp
pbxFGC5QlQyhBItab7xRzP0z0G0su9/VZmHDkF/ZpY6UcwRdPmuDFl7crBct0UG+
E0SWMnuw79oymzKjCjCF46Mw5V3bkHRcYwMSsEOJPYCc7EnaUs+5YD+oP+WoXi5M
flEdEShuSIc4Kgpt6EgpLSZaqKWhlpBYL+5GFS1OsK4AYR9Yo2U8j+pSUMDiBFYf
4HIyMua0DqVnEe3pPK3vPNCoRhLErM8RNd7UEH3LoKVlGl5YCMiT2VwSLh51f2hH
QUmZ16tg+bVT+ZEOsE9eXn6kkxOOrPWhw73Ga3Kf7tUEnDhAyTL5d3NhdAdl35WZ
h99SBR84/Z/ftHil+h20x8B7hUaIUD0nnRqAeQzIEQsuyX9PbX21VFNlUesB4Ifb
LNzIifskj7J8iA9TFpjtqVMPUuvlCVvPmx2FjH6Iwm6T/MclYiV+iVDun4l/eDPj
PUDGiE7Mnw5X4D6+jqvJ0v8WFDAGlfwkBfE0+8gp0HeQY8Xkoq9QvmduopjNBMp6
iOJiAWpvWtGoU/s29okMLZglzxCmFNCH+xpCVez1ChfL55+hjShQmN/N1nAaUll6
tL7tDUkD93HrLOxr3b8gJpfcrIu2M3TgM9c3cvR/huLSM7WZIWX6WFwRnBFSIFfN
uWV78BZKZ97rZ6+owD6Q+nXmQo2accWervx8xuFQ6lmmuv+Sgp4qSNj664kLapMW
Im9nvyRdPScY8NnSlG1CxXob9x5QJCU3b1nbPYhNlKQmfLrDijP81KznlThhRN6L
+O7u1g6nwPeKJBVgMYzwaVrHzckmqmlNz01m9SwwbhHbzHnRk+6qy6aJpBSvu5DH
de5Mxxpe387D/VBgBrrl0e/+8herK0x2pTaW2WbMPI9cRtEksGiNjkv3wgnqwSi4
+Oy10T7azfn4bS4MwdxtaoBHBZl3beD3im87KzV8elCNWYCibtwu5tCc2UC3p0Z4
I/KD17ACEXTvrlISkJpeNhwlm71nDw5AOep6/tZqFrAWeh7x7idjsGXAvxv+boei
VEeDQ+e2eTA7lL1/+TfroUW2Opm6Zm35vd9fqwOqRKnBbi71kOSg11tA10ajxULc
I6Qr7dcZ/Qm+HV7LLyRn5f69mNJ9J7+JxwUf2/75SHcN4PDH+Kbacm0pHxo16CMu
9u8j6ATs8bI0FvujmC6+5L42+ueMVnoIuUJu9fR2iroFAmHJmridxnSaN0du4/IA
yn7HNVkYJkNKOoXavs7NSY+WopOCOqmDH5zeALHTYyyusJwDR6ISduS22lnU8Po3
af1l4XnVzRz0R3QIRXz3a9Lxt/v+XKwOeNwvFx9UGDUxgvkfJyJ9VGvy5QEkrzPh
wr5CMLxADuiGqOg+gxT4aqItJHxmb3OG8KAvmd4b4KpEmjER3DdqCcfmwbibiDhT
AYJcNakwx2IfzZW2hWtXIudVihgc9YiIm+/sa/f9elOvPv4r3JrZFpB5sUF35NJn
1vtx1UXED1tEI/UL/3BkW7sy/muvHWcTPgls8ozUaFguaHN0YjTuVN7CigGz7Tex
5Z7JU4qrhgHS3nQ3LGh/Q7oWJpQcNOxwrz+/SYlM3AVgYaBUvUE1iLwmqOAV3Pd0
y5/R/kOCPUaVgwOJ5LWGwrdQ6wczwh+fkfL2GCJw3giaKpoLfMhPh3QK3YvZHE93
YmzYnEuYzi5IQLX+zWpZLKuG8VY0HeXQ0c5fXbdOLU1FAkJEUrvbQzjHEjmd9CDZ
evZFpc6tao6DvOnn3nFL0V7f288HCTqy1p5W4TuRKRt7j5WAciLmTIsYxTQaq+FQ
jn5pIrTFxPOfPhWTpGpAm6ppcA7FXF3JzqkhD0YQJMFCgtxzMXP73YCkQ6ONqZwT
6W+aHOeG1XRAS03uI1gZ6xLpW+m1NdgJsqK3wAok4vtQPMbcJb04jsEcMvLsKSS4
i92hFtkZgX2JO/P1SywiHkXeZxQOX4KZMVYeZwzHTpPFi9RGThpGsYO8zobA4lUu
09d5jrWzJpOqt6RxH4PD6kLEXLfyGB8sb41tCvJZ4jVJm3Vrvwttqht5+VmUXvxo
JRhY0PikI1ig91EhaxokTtDo/g/BJG22SDO2FmMXdJpuHhyX+2cMCxZWYev/YgAN
Y2Djln3z4pj8Bo0Vx+dNORskIxxbH0wMrLdPSjcTZAS5GktlOPqRxnq29E7qP9Da
d6tiZmad924Yk/B+afeQjqxCPeSbzNDd2aGviQ83yH7z7dF8vlmNPtlMPAeXHnyW
sZlfmtOumMrPVnWPf78QYFIysgcA8nNgytxxgLPVNUToo8qTVGo90vErpq38U7pz
/+R0UsQ8asjt3A+wdsbVeT9ihBJh68wF3TrWo0tlESqA6BhLezB/WXeiAvrKIxWb
1tftgEIIq5c890BAGcAAG7PGzmapAfQIvR+oaVU9kTlaru+yUdtfkqtvs6IovgUU
VOIoH1hsfw73klHX/c9+LsUQvARWJj6PLlmN7d1DtcvWnJCTV/t8ozl+LBOufED6
ffDQ+Rx6jrIcgJJ6KNuW/8zFIZv4y2B/P8GKehylai3CHsQ8bRGE4Gp2icoDRi1N
yFuigG8ke8G5wofhE2aoV5DiM4bv7f2OxjJ+Y+aaCb/93a72Gr8hAzEJ93Cv8mHG
AsvYvhqAKUnCz9is+tb8QA510A1m9/FRLyU1H+Y/aYKIQ4m3Yz1k/TdX+kJvZxde
GMu9Oh9VIn2eY2NlVgvz8FWouZaKAqjdRhxk8NSeb13ApmbKqhRhJeDGOWGQSJQP
FhHzmGkvnpg/2PVn1UZ5+C0p2DTd4GMuhoPUaKiEQPebz8FvABJmbQbVgqtI1zfx
0IKd+ab1WPcKExxdPMDHlsU5MOdFXu/WpBInkxXWr66KEpVGp6wskfldpRGYdR8S
r6Mk1KCVWKVMedJlzODlevEb9HDUAlVqpfhWLL9lqNnQlSPLgvoVHnoeGqOBhlxE
T2xYUnNcTy+jxyjzR2dekTomRXpOeyH/p7PrDWPPHYcnO5404vK4RCQ4gmohLf+5
DIpXPEFQMYnMg1edAd0OCOEPQ2cj99bCwM4ro/xzX5k4pduUpdTY4za/siULN+jq
Gg6is/UnRq/QzfPWVC7nZs+hHxXmoa/6JtqP5Fo5VZL66bOVGjoaJvNvvYnK15kc
W4fZ8Femx7hS/9DMKaXYSosIAjPxdMHt7OuqDu0FAWAFcya30UaMqCh59qNgb8u1
YMXGDAxJntobY589xOCJnPBdAfsVCnEZ5t1vOLE/S0rZHRzcMpb/4eacDiUqle+h
qQP36ppGWe/9usUxXOTTweS6g6d6vcTIh9Li1boCahnJu8+lGhfJBASG/JSIwTyz
LaJlfDwGbPEklA3qIFNoud3CY/1UDXYa8wXcHsW27t/wgPFpDSvHE0YhI57BL/M1
wfr+l8GOmOk9rd39Y40M7WRcXbEauzGdeZtTgjG9qURkaGUu4IuOl5M1BKJsBBxQ
8h8cAO62jRi+oeFBdUO5IL6eIksuEjQ726W4wtgtvH1SBQ/ykg4vLH5L7mC4Aq12
7y2t10M5JlRXADKXnMVMsWskrSXKMoipiREFtuui9i+Z64zLD6sJ5iQkkAYoB2V2
Im+c94AlhyspZvEG9Yms2eXJuG/zgJDiz4YSCI722U/dAhgCf8RPuWAvALe42/77
G9WzRc84tKZxgf5B3Zb1IoPuIGEoU6yZK9yimlI7ELMiuuo+tdAo1YaoZvXIeWFY
UwBM424iHY+gffZHGIAD/uupF+6t3be5EQQcwpbo1Ace5d2zgwYUvCf0D+9TQLAD
Q+K07WTBHo4auDzCUjjxsIGx4QnaRmiQEWoqVl+h8EM+JR8q8/vMSd1P9e3Na6Yw
UnPGLrzbv4M+/tzaALHMLg8joaVS4PlUEFATLepF1aOdPrGNFZIfj6pLOo6xJJaS
AR23CdxulkwZv1hpTsCFG4pa0r6EQq2lTDK7bsUQh9QeDZLTSFzb9YZiSyEdAXUB
MbREA3OZnoZNHDHzu9y/4g9U+8NxljIzWZFcjrhBq+OcoUI94mqv66VM7K5o+IiC
Q/jvPMzg9z3mdqgdl4KlNHljh1h2fakkVMtq+BjqEcKnuemjXN7oCxL5EbxD9yg6
FJAZf6FeM1Be1vui3ssmjtHzebmyLy0iT10jv5JxvNjUQn+NX1KX+Ek5rObIfidk
7oSdJRVn6JoeITcqmOVCEtDa9qqXy9sSX+piSm7lauSvVHxDxg6PxCpg88usSQNk
4gvJVr87I15i187qL1IFtZlCIwdzLq1Ax+3s7Iq0ni60ee0bCr3834/5Qf27FOmE
xBgPLZf1USh8OhZsZqcea28Q40rkkUhwX7U1pwg5ubHs8POrK0W//Bp/ZQgXywGS
eR8S9SIEVDGcNYwQM9UzV8JKR50UMTKZbcIPVxBFyFUKOP3dzaeSJNnvbftSdm7e
1sY5doj/TzkOJY/6MWV+h1F93X8i0xBAcFCgCPDEOmoFytQIhR9qswHEI5z2+O9J
LQU2EY5yjT6YkSZO4fr+/WoyaDg+FnK5ARdtXS7C+9zxThO5ebwkxhU0U+OqNJ49
PRMQtd0qudCt1L0I403Z7RJk4bUj32SopjoBT/q6tdwoAMgsAQoHNper6PmlNSnu
whqtUr2jP+akxrBMSr0k0dX3LFgXIz9xoI+5Xc9p8T6wVB80sLx55XvsOh817kv+
QSNahS2t1BxFGukL/sZBBrmYOabE6i+oZpU+lFxoCdrsWfNi8JsIXuSdasF/iiIi
83ML+Hw+oKreznb8GxlcMDwQo9wMWlYl5hO8BS1qut609IEeOxcrcmR70LoRnBNt
grkorkUmnefM8Fh8KOpDsdNjr/nXoDLN3wNlFr77hTQqWSBgCZA1d/7p/SyXdQin
Lj+SjaR8avqqNOEURlF3wxtTuiN2v2ah4xXvgXHnk/FosXU0q/vgsK42KjAJ9wyh
kOPzpbkPRjRqib00oOf1/HjINz8e9Vq9waigU8dLCYimjSARaLY2kuzUGAjMIM1L
V9miNkqI324cGthvhvReK7p/uKyi46zPHq4SI5eecKV7QOaozhvl2N4PG3KMFwM0
vJeKIs1v9gzNoSTFRLyF2CEovQ8j7twWNz61NM6q7Fsfhch8CNDqUGkeOcABC6wo
u754INZQ81JXEYM/VIwcrH4dl+k57rQzl9a14zR9iT7VC5U2e62zKgaG5wg9qm8H
CLv9n5/+we55+cdON3FOi79zxyfJsZh/vJ9xjp44HEg4nr/NlWFkCMRIUgubR37a
ueBG1eiY+I6tcOa8qU82RnlNBHvGTvNObndDAZ0WLBuxGsaoaZrkqqShT6Qv/N4C
q2CnGJRQF6C2p4PNEjltf2W1Eq6cPTPd0kZMsuW2Dz11rWBG4bTvCoV//VRk2ULv
O2qmzowEXUGkOjrKQfXdUg0PHoXuKfc1oW7BQ5BDCGiKNSRwR9Rxe+LL/xPSxfmh
XozgC4rdnmf48JeNbvBIv/85BCCY5s0r45fscMgDKhEqI4tNsefUW8QGX+l/5VFR
3itbJYHT1c6crrIkPRuwRGVmxe46JMPTiyZaC4sVMQk3qAa7si51hNEF7QCVAK80
iNeGmW2eiMU2+kqlmvrIQyzUpUlZycpiIMj70/dCfAExZxDnnEoooHuTfX82RfDm
gnH/nJVXEON3wOvNFJSZ0owTF5175b3zqcMEoAUttXiINC0HsNSqcEzOhEinpYyy
ZvIndkLHFOoPtr74hCVX+2wfzvFPGj6B85ZUQa4jNI9FDUqGqb5id+/2sdhqZXEV
VJWAjk8yU/uExSZ3/5qrQdrlMFQRzmRWCm+cAg7f0TpXRXu8On+eX26FVtboBSJi
oEDHYA54ORzmV1W0ByKNvRYpg5FSgxWbhqHIU2pVHXT9PkB5Cu6VXcQEsTvPp5rA
r72eyhivGUfhFrfhjW83HI5G/lqskbPrVtWlgrza3ydz6xZyj6w3NWd/L9ybMH+m
yi8qHYHPw1Nww9l/Jj6xvw1bwq4HssMl409do9eOz2lsjhiQkFCHKfIs5whOxm0g
5kJtZNrQE5FX3zBhPF0J0pYSRK/7cO2qvO7hyqFzLrce/3iDKkhCmCVT61U+obA6
M7ndWrM1Py0EL3t/v+8+5kpxWmxR5w4QlUlAYBq15T5bmbnu9ObOOjwoBGPiC5EX
oUhOxrlvaLPIdkXXXk+olQx/KJtU0InwZFDCULffCSPGSCGKsAv+6Ymd5kEWNSIf
2dfmB1BE8yqwvJXQzmi5F39sIVuriWgg2MwE9pNeK9wzxuztrkpGNQJQ0S+yHD/v
O86k1aTwDtqhJLLy9Xu2Hd0CkWEHW6kmU2kyKv4npdMTOEMBy0oGGz9diflqzr7G
6A9a1d1pEtakfX91TigiaCPrBtL0d7DE5FCV4q8Ct3e0GEAC5g/j6RfXOAFsB9Z+
MutIdaJPAggOULYGeeTU+Tg4nGpJY/Mad4CnnTYATm4TkYtAIF/qwpdRArOhbs1D
IzCYz0hgzzHpwBkbBCzS4cycrExKp2Yv7Z4RjsQVXArXlGwl1CetHP+sWQ4c4TsR
bPORXQYCvafVC87eGg1fMz17GST76xzFUbZ9Ke/udPK6qq6SmRsSGVGr/V8RwGwM
fGyz0N4739uTQA3UpPKpmzLmtA+K2wFjTfi7VZZ/VFxrAj12Ga3JGMA8c+nbUeLC
0LSCC3QAHn2b/qhidIZD4FQtTYEmYJhV1u2yrSLC1xDugGkkXJnyURDeH6TUjKG4
c97TMUIWp3a2X4OMOySUPWNJlbc0l/osbZQjlpzp0X5Vm9HxeK6siQ8Kur2cV189
sj/O24KY6F2ut8sQxht3Gy+09M3etPZ8hV36Q2nFqrSwXiPxno0VQDQHulKGvHzT
PTE6eYruSXQnUHoAYCm6knBNTNpBhqHsQaazX1aV81vx76/G7ogBJYZsPd2XbWmI
XnMAAirOqekcZvN3tK8vUaaf6rz6KmJWNNRsnvjpQWvWrk1ACW1dstFckvw6Vj30
pxA3kKoWCnqzXUxCZlu0hbgGCfoyO9zEjffLMA4z+YeasMe7bmrsKP1vdKTIeZ8i
6B22XpKufExyiS0qZTS7+ZejyZoTj+gMQLsZI4qdeg5QQE7wF8UftPIEDt6j2F7b
7SzST7DeUEb0wVhpKme4C7fLBkqBbaLZBndz8+XF/ZEkQy8doJ9FXdOkcUyV878P
uWSxGNJFV7etphC2r3ivX112qvY5u4uJ+tY+uO85G+mwrRiYa1KbwIP7WeDyBbq0
DDO5IAW1RX7k+2GStR4Gdb1V/POlpjH+GmsjdcoMEhMHaQJNcUF4TZcN6bwLCWmG
IhqqO/+yZJVAQOJOM6EhJDAaaMBwdvyLmwiXfPfhb/eqMSlQI5QDOl0ytOLlTufJ
kIM42V+Ro1fV/cZXzluYxnQRKt8PklvQkpSppUo99F6Sf9RylkTTnu678uyNDfhW
+zNLPefaXNrpWpf9JEVGzHLhM1+BP9egZ753YYVIaoOzKoYfzy+AY2IRxDV6DRwf
/SxKTg1W8Ml02IB/nnboCnM2HDN4NscuSDvNmeyguMrdmP45LzVWoQS5obhzNsY+
sJzeg2Z1NX5gzFOvOc9z0vgy1umlmtfPDv+brfSThQlaRf4FM3YStV6gd7owh32c
6MgUxuH53REOiXTyYFUJrHT8sZFQjjJfaeFysY3XxujdjlyHFmvmFNy1CofzT4rf
ToHtkH+QHB5ko38/+9l/P81GPBvfnI3cat3iDuH47bjuuoZJ8bSnB7NdJOMODj61
mXEdaTCcLHb5l2IXUgARgJGrQImVJcJIQbl8cET3H+U0IqAp2M5TFBuvC7Ltgxs3
Biv6HuAg0upZxYOSGQzonwLnJ7fKpDfbLt1KcmK9ndoHLW395ktJUgBOZntmzw9O
/8bAQp5EFw0FHwa6Zrp8gzF0SVoEW7qpk9/OBhfzmCZ2Vdhnm3ENbu0dc/N0/tP7
cvYdpi9gSL+BCdMXbhAS1As3cHsKxesYeoCrDtYOqIA854hcJ5gio/LkQaJMZoU2
JCFDsmou4HrXvvV+C0qXGDYX9n4111Ivlz6g469VJ/li83udGcEcoFLP5ZCaHmXl
ifEmzeamfiZM13XZ4EP+FBodsEB8LEjoiEGFiEcCEswrq5+yBBOw8tZofGYOO9qy
XL+HBSc8yWKht+IQdY9vfbjlhMJoKChd5as10u812b3o6l8T0HT9ZomWAyqnRGqG
U5JpSDcOeUMl1dU5q/OlzrPTGPqlXRWrWYe+epleUUXKZd2k6KtW4IAkvTHgIJAj
9t0Qf0z7KmSJidpy0inZS1Yz7h+m+dcst604319rvFT9cJF25f+C1wsbC9ER2MaT
lCMIOxEfv9C2aIij9LGI2+9miF4opDzXyVRDzHzveMYDcJUBhNFarBftF8QYdj/r
qmPF3Zga9gN/Mdai7C4NlHNEaxSKRxYpaiKIGeuNFtxG1yoAItUMa0jcgdGnq78Q
P2wiAiAi1TZ+oEtsM/vTTGXpUYzLlCgdTvGP3QHkcCitZkxv92oGWaOKNUU6x3Dr
f4y6DdADMkq0tWaREmTWlejs4PcmQ0v2OdVE2mxNjRez6miPWSjXQMS2riqTcqfK
SEZZoiujYYeKOzhRL7C2Q9mFaC5HOwKXZQVDuwcKxShU17aYiRBEF3KTO4gjBFHX
yK2MFw7hAl3Kq1P8wUYiUZecsLVfbMexvnNxnAR814I+TRSdYN7HE0X0mwDGPRb/
ZHnSyiNo+rbTV0OeAgncp2HCama4IqLx/kc3Mnu7KgnguFFs3n+lJMyCEM+zhbcp
4G7NX3a8r1MuxA/GSKctd2MXNQSBEEntitgn6/LjAoxebfY/20p8fIh7cx7Fzayr
k9W2NMXCpxiWaS9O03TEtkuKmXW9JffEPAv4Z9mSBWE0yokwBop6g87z7yHhjuMU
Q/fqhkI+rNE6lqzMZ8k53mWIQONa16MPPT/OVjlRrt2qpK2+lLewKkNJy4cgwmRM
Luz+ZRWNaMsKkFxUua9OBoyNAOVcVhLIuo0Fi08pCm1TQtlzd1jRdMI9Fs8+/z/P
fR9ZLuRBgB5MCNz3NgiJYLzd5d8bhzHbpSum0eY5rGJqkpaxdGHMG+N+WYb1lo2M
P/W8NLPW6PxyWJrr2PqdOSzjF+6X03pAAIlB8ciIDyltqqw8HSqXupvRjCw7OQlU
G3TGH//Hy4BPNjUvqzXFmHub58vmEj32bgclGuk08KBINH930yVyM6wDxzUqOAwl
ZsJJ4cib1OLDW9QOKuyu5pe7RPTCBaAyOxnIkyQMqSOvXa0wmf9maF6hG91ExANa
HyQlXv2bVRC9m4MivH/shWZXb65TvFxROrESO5KJnec6V8J7Z+hQPQA6ddyeoFBo
pKubH2BIHxTz8EHzWdx2Yeg2uEzPGLHLEzU7/eXeTsM3rmVBf89M9N6xmsicYYER
7qW/lLtYBKzIWgN8lONDmz/cV+iGE/sDggjZjoyz/6Wtf5K/f6Dm+iVUUB8t/roS
vYJ1m5whuQXMWK2jv2j3+HdkjbsnBIMJTBufnXV4h3sy+oWNnCSBnBw1teaTrJfd
dzxd9IwXCe5RO1EfGoJpZIG18OjVWa9cm5nusxHmPJ12MrXnxGciZQ++jfOwPfO6
M/qJZpxrBufmI8Z3Ju31g9TOs+d1aPrTCXhuk5QrE2CpuQsAUZ9xfPB84avRkO93
DXNPXEvSpdoxAx53LVuQWKws9A7k63kKV/Xb0pdIj85VDO0dF8tUntLmIB5sMxWt
IcKrnz3+okTr/9BBR0E4wZRNVs31ub4z+1gsrLmsne2Mc+ziwEvwjqscLkFxcLY6
p2nS32BYVmBaSI4wEd0pGEaUrmCzNKCOz/iaFSMbaJ9IgyESJ5aBBC6vdIdCuVXf
cGIXIpsGOLWrEbucj9BVy9T14VLjh5d+qcmcEv/uiMjHUNzQ5D+4Rs5SprNtT7Kh
SjZSbY6uV4H3yIZmih/x9EMmgbA7xx7CgtrtTdWbVFGxCR0f1dmz6HPthvm7RmVN
gRYvPVuMGkwrCuzIYrU+PL33JLlsOsfg+W0NBxgpcB5d+rXDoYGYyYoEqobjxYms
uzfclq3uwckgtAivnQD2YfCsUDml1Yd/DKzT1S7BZQViRVNguqKnDgZiMeaJvtKf
bbiQOHlWNtt8xNF7vU9SUEpH3AtsIGSlnRS8SxHYmz+dOzfNvQmN3cxtwe0LSkxq
vQayPm8H4Z/GS7FaPciOihKz4LTSNxQwCZ9EGI4+y5fCe6e9rd1xXjVHG0In8pc9
an+4MJLEApLYD1FLXGv3dnWUhAxX+gIFScf105Jik4TxC02l1yj6j5OUoG5Zm/4L
Z4KvZ9gBdTFx3ZgrCzEeryNDQsqYzOsHsYai1PsRVBQkXVHowQHeL7tspuiuRMti
raUluArvrwTAYpfuErKlig+LqKXTW+sWR6HCuf+NiuyC4Pj2EiIRhwMRWQH/Nvue
yTpYb8GCIJtAQ5JOX6iWxdRRgmMsbhdn7A0IIRSlt7kaLSYKLqlaQtVaVgCY5x4o
uw/d1t1UqcHjkH6Zusu08mYBKSeOxYacb2UiS8mlD2rmGORMvac6cTsQr+0sn5Xu
AG2Gy1G08pS2SKr1aCN+LrN5VHDwrv6+tKrzBTmnOi7o3M4sxt9ivEAQxrd7ssCV
d4IPxpu1i5w95lFBe8YURkdj9b4QkGx/2gyOaZad5FuavoGUFA75fIgfaBqFCWXu
ZTPsjEklRsD3UY0OF+UUjF9PacXviY1eH5ED4rJRelP06g8edg+tDn960x+Fr5sP
2uwwWbYMjiG3/oNC4xnDxP3sOho5d4vIU98Yz9cuB8tPcSPBT65boFFYDRisXdOy
R9qfR4I/cbx15f7MARhSuwKwXLnfBu2YOO4s0Oyr78M2q3nndLTZgkNcPs9k8lpA
sS4Yv0LNAzF7AslukGHus2WR2XvzPg+jJrmcVsuQYplAvskTWjIrv1joi7rPRaY+
lTLPd4vu8LgUCdeF86bFXk6Gd7zUsUqYnebbLtz0v2AudGWi/TiHyH4mpVMzb0O1
J57yCdWKJoScswUWzY2cWkqE0iMCmzPNurAuZQmvrMLkxDs3nkejzBPCxsjqMjcj
NIWsdUAbmcYh9Hp8SHJP5UclVTznoBRIoGK8Nq6MjlFwxzCfXI2nBzpNMQpZ79JZ
i5/iMYO/QHeGGReYDxRPqvaFkZCELl2TMmYm4VFiKPgn629yYnJUVvBNXAThzMvG
V8amYPcOoGtaMhvWLfL94ymKI3mMj+djqIUgm/F/fJ296F6tDemjx0xi+gka1uOJ
Dh99/A3eTliRi/W6G7v3SlvmyWZgnSPEJknJzV7JmCEvw3SQcQz75SaBKtoHvUhl
vN0UNoSwuPVVh53N+IEK+npsCUBbDe/sjRisiUFNx4yO9DAuavLKux6TEM/PWBz1
AC2U8JKLtgIhDZAz57IIowtcsXEmeQYdyNqNPyzwiSo4D0kX8B4fN5vLw8dA/fmj
tP/WDnwFTxmvjHg+uB/iXQVlJ6VaVLtem8BsQCFGp4gazw++KTteaws1r4X+QZaH
E2mZsIajfKlPGhZX4nu4GToyPGx8WaBFaJPmIzkwcObxEWAJ3ndVEK9efDOfjDUD
G+OPYmjyMTc0I7z9jfTRmP2gaQwSzNW8i6BKk4p+leb558zbpTnBHbSJexn5yfhb
ndgi5dMwbOK/kYHbsDgPRfdfDjDAq7eubrjqeeVCQYSvNaN/f71o3N5Hnp4RBbPy
CziOoewyIri3m6rsmX/ZcliNhJgGnUZz5VfOLD7fwGysddLVPXLA2ts2dCteY0s8
2zvlew5N7DS+QpSU7KtMR3w4/VIjU0MkW21qHrtugVGs7pgmJcgqKsSChWyZcqsP
sFOolORydYaw8pzJO/I++jgabkMWbBrrK97QUlt/flsnKcrxgHpsEolPibmkA9yd
Nj7W4Vs+Sa+mgFCTqFQcdG1w7SiWHjtNKcethBM/NFysqymRdBwP//Lh4/R/ULRl
XWLJW71Xoq+76QIxbnJIkKvh+WuMOGXUE4ELhBPXXhQV0KZ6mbMcuvfW3FveIJIA
rDL1rb67RcUlpfLVqut103T046oneQHSW4Z97a5WeB71oQRcfF8lcNuNCu5johEd
g/6g5ld+ceurifPwSuXVvQopDHqehf2C35tt93aqMnGbMrXOGUd8R8/VbEB9iW4U
S043heZJzTh+AV4mE+wW4HJug08DBK0uJYtj3WQBOro5jz2UZE2DrPns8f1cSatS
N2CDjVR0YePheqd/HpdPvutYMwoVqHBW8sxhY8T57AHihxlZ7Gpd3+1TkXmuHkIE
KinKFMX3vKEzzP228DFWKEstVftyh/ShJcyoi2hL6oeoyK99NAn8Ip2b40etmP4V
rHJRG4H8af+A6to5vwImyeYAP55vcnMxSqu+L/nunnR6jar4ZFmB68NI13Nzi/H9
SQYpViWvmEJW9oUvNyqRCNrnON/AqFdPNUzL/SFBs9cDhuOqhcBooR1190/PNgEB
gAg2CQCDLJavESWCczsTctuclf2W3dYw/rXV8p9uTGzOkkShMlcwMrGIpK8gPkDq
MZi8CBpDUzMxoX7bZHnxspOzGVSEU5GiCQ6obtQhQaDguMGqqBh8GVT/h10/p9HB
q3HGmZ2sNKWu1a+8nZLoZIlAYFr5n6Z7KUDSJORT+BHY3B8R3pn3iBe6kebpuF2Y
z7yTKdsN4rIueZM46Aun3BZx+AmwdIpCUNoTg/573PK2+USjSP3K0QlNf1Xs++8A
9ZyXJCuMl/igE/74sFV+eFxhBRkyy5hAlZpEsp36NCJ+ptjZX9mczT8BtyhtLWX9
sigmopvnmYhrI7qCh5rU/sqrW+zMqzLorL/T+YGxlSIHRLMq38b7W0NYm5zjQAhF
jaxuZ3bIcvJ65QwwVRrcSrI3Cq5S+0/OxPRd3t7k2CbztdU86emctL85mplvPvfN
tCQ832OHEbBlReRzAiRJJ1HN+U2E82a3PKjlUYMWEQ0g56rZYnopIHDBvLWEsMAV
3ni2yKMXbWNPCfTUykLdcFvaAFbpyg3GH0OBueZDac+ha+1vyYJAC+GLluMH+QCI
Uy2XfmNiV0h3rW46YL7bzxb4BcTktbouKyNyszHBCh19Raa7c0iHtdqZvkaN3XaN
+CanO0uP1F6eN1pQd7UU+RF/KKQ31k9Ia1vGIeYMdia7GCDdg+BdUqyLGxiYRzkQ
5RrUXwPn7L1OczHGya0Coa1MLOZ0mzKDD24htMF7e6sqTEP8J9ThwTf7cJhdCCzv
FcqGAJZ5EPPVbYrjpmmk36chPdzmFhOMYMXKyatWeQ9Nf7VU7VUhtAP5gVTh3UPU
7xPh0oxIcD459Fvyk0ZeL/2DabAOqHnPmE+VXazELgsmLFkOs85NBF1gDfhxZlSV
tfbNkGJ0almkSPGep/wD2bLW2i9kdMB76CpqWqorssXQlBlVudK0qMJI7wJK9knb
y+/GADtHVjlP9WFnvkL+8PpLOwcTMtFhDmrUlZxVRoA0SAZGjLtRXpm6T69X1HI7
h7ujAcqD/bMLvZQRHTDgkbYRvPS1RLlcMRF1sA3BArLAQ/zPVEjPX7D2cM1Nli3p
OoNoIhTmBFTpHgBMoCL6xA80cfWSWF9fDP6am0PLPpEsi5Fz8KwdaWtZKGP18YgY
vl1iL6n3C4bcvPXZY7CoCqd/4WqDWXik4ImdDDjYQGWhQss0A9EiW8t8gKBjej3K
u3bT69X+a7Go+kJKhen53XehFO3Kj20hvepAmG5Mq4b5MPefCw6zZjsEs6yRwawg
uB3wwWKJgDkZIaqA5s2WEXtE97mIRZqfnEqPm0Bv3k8a7+teRX9Mujp/BFZ/Insl
y6QVpM3qJ28mKKXIVsYIOMhEvxoooysBgKwfYGaM/zt4SN1B85TatBmoS8IQku57
ftv3daMX5d0iJRx/uIQjiJOI9WZowkg7/QBa4Bl9r//gpxhEMaWSnmdch1OI43vl
GfTrEvV491kfw5R3c0QGzC9KUYEq39vk2RgCgqx+IWoGZ22m1iVg3RWPlwYi3geW
pgjODoK6BbYdcO7mDUSM2zp8p+mrCVwBrqxIJXD5RqAkr80AAINIVW7IDkxy/go+
WgcMz3gg9m3QWWSQ4VNRRZukYBsKmdIHnnTFsaIv7ES2ZVtR5spUYF1WuZWcqZ0Z
+4fvHlUQ7c+PP85mbqo4tNDII3smO/JbRUMhK7jp8zl6XbV1Xe1HEUVmaepLObs2
0woHNzizSklN5gamca7u6nbVoKqDNLLIas28zFrQKFGwF8C5XZNWbYQgYtX/9gr3
YzFswXajC6DmLQPFHgo3ik7xuhiwe6ku//IdTH4zldxvwUz/w+Rh3PHKuppreSPN
2erbrUVvPXZCsHQHKpSMq4gnvk1CXhmazdIaCy+DGBCEsJdB4q/2dEewed0DNfgb
oJn0Z0CGHV34rTJg8UANbnbXDugRlx24CvgWauurc9CNpJowcPh7qiv+bzWA26Ge
PDHmUGtMX6mwUZ8f/5NgUEWhaEogULqiBuYy71FOJQxClmy5U3ZZCDCTw3kfyjjF
sptjVu8l3GTpUYrD1fNHFw2jVYKSRu4uLKdg8E6nw7BxqASosrUAcBvf5MMbCe8c
QVhIbU8aQ1892dI4kywRzP/zowZrJbU0mh8dKBgEWDHU0XWAcaGf2NlFgcN3zl2+
3MjYFAAicCAQAKMRpsOxcB8rfxB5NqYtT8EjXe3vAhZBLUmg9ZTStybYyDRyuyjo
g+w7AmicsCAF5MsTrn4ob2fdLV1oTyZjY+fcDI+o+MRVBjLP4KUE+rtv++D3D6rk
fY52+UCThTky6yN0nzpGfoFtUO9JO4CIyvJD5TcAhAqrJCpNMUMHZiXLhOBT48sq
4vOoGJprd6VSd2B1oVa+67Y9ULn5geetSMgZTHV8S7HeQALvnVD1YkeNCturTwZp
J7leBHOTvW8cqZ1mvahsF6z08/1Bk94doObRdl9VeCIqDAA78f6yhRGjhXH2yJnH
0KQ1CpgKEmTR9u9KxvP+yjG7FxPRM29IHUOhkbs0jFsqhU0H/b3BTRvqsYzKBCVK
TEtVNzvEK4dkU4eEXj+04a/2QhbeijcVkIr/2PvckX9ZvkTwSRoG7uWbP+MmqVyv
8HDxT96H3oa8HrFiwcWlXpkS3DUeW5h7EHLy35/6C8HOAkYZ5O4m8S5bM35pGw5i
BoklR59KRJ1S83gekyONfJwqMrm/p0GYn1SQcz+SDq3D6H0z8q48bKkeWps4Eoc2
mCVVZDGEJr4VsEco2pebq8IBIAOaiVN83+f+hgreVEZw/2hRAQOjcgCRXIuEbC5D
xKatvgigxy+7JpxRejlFPbOg+J6GCXLpLBpaO+CN8EPfHaBWpPSsKszbphUBMCe1
4Yhgq8GxmqZ9yzV+ODxZaRpugcx90p46aJdnJHNGbIC7NpGC+YAqe/fCwt5BSb7C
ImXqB3kvk93iheY2cdtvgQWm2U1ilSSPuVilC3ngBkl7wpfi0kAee1bcWy9oT3Ff
kNfbUNHSKdlRkT/Tcl/HdeNh2uHmy9lw/6yAANJl9Ausamr0zu3/aTk9w7ZV84GT
ZVTWDIIHDPs5YIbCpUoJZgZVo3t8CDnrFlQo0YY15k/HTnMZbmdSbTWqGRvDKuWY
KL+7e15n31ckYaemeOU0DHzjTBLihlxILPw609zJr+0JT1U0Z9Tnh66x1BuNppKK
4pCA3eW9CwVzwbERBhw/Dfc5JqEfHOGbDQP7tmtHDs/jk9Kg0qQVIqXPib81c6j7
zKDCBu9QvsOPGV0GL4ta3gSJZuCE/OgmvKmLjkUK/MH5fQzeZ2xFqYk7X8xojEH7
tGdqqSRdlU2gzSGyDOmn7qCWtfZOgHR8d2945uFBGEJ7J1ofv6s2+L1eMqKxGcie
/mkJlMYs2B/36pF3ehY6v0CReyKKeYOZ/gjYhKoJaIoqn9ZB6wwiUHEjFHSwFr3/
7a1Ccc3Ri5JFjQiQodoV+Mmlm0eF8Kx+XBzueIQqKLj6VSBYmtKvzFyVtPUNZrnn
tsJDDX8Dw6G1L4wR+pTVQlnGBFzn5F5wBzKkf8OO/FLP+SqeE4aVA+LPUgUIQhCE
92Gu2QLfqwkZtc/hQiHg5X/Z3WAWwVbNBOOlzDCNbmvdpeH2CO9xkDXuEYh65OSj
wTs1ihAsnh1G9gxkeXCMpjzHCYL9mkFMI6Ikfe/4GbRtTRVhgfj4Vy2d7oRnev+T
fqFzwk8c0o6FlAA2swy9bn/Oi9vme29B92AY5bSU8yw7kXfkzGw6FeHE8MQc92HL
hXLsaPtqavplX0soI47elc2unCuBSGRRQ3aQlgGs5woX/+pXOyWNspxzg2tz6Pv8
BTfnOlh7hATpmExQuldvOJdSa/h+XSVLXz+YaAdNBc2BRbZ7g1lYTWe38PbRNB0l
T1n0oDyrXOsRQMg+L0khXgZ37/0CwYI5WiK/KKo0aIQVHhFqZmrzyhXUOdUWEP3e
awA/sWegNkbyx9Sm0oJBP0Vn/2t0BfuSRvshCO/FCx25aOyP65WezK2v+QtHKpWF
EBvEK5rh1lQsxxEB3H50ZbsE9AZj9OSNZeCqYYjj2xlx+oTaaTTGMqJff4wfkGkI
ylFe7ybRb3a2/9Vy+iUBNOEUMMFVWX764seIPZo7CccU000LKsn/ifhzVKzBmF1d
lq8ivwDb+nyimLXZpUOUXvFXO1b7b+kJwr8m8satnc881g2PLjYQ87yT3DHwammO
HTvVYoNd2MgZz5tCViZc8bWa7qhEAm4j/Xev8jqRFdAaJa0DkR3DE49kr5OJlEgc
0Ql/Ov/LHfpDjXwnViRUh1yw5bwbNsFisixvo8e+FKfcttM9kY5v10E1Cnkgk6yr
ulwbjkCWVjIaUz7/ZHwZ5hZBRkghpzVUgAnXYXIBvJ2EWHj/R/XoNnKEaPWYLmvv
X6LzbPbvLrNj8Bbeo6vtL90A57qD7VB+CQMaOjsHDx1d9N/C0Y35W1xWf1cTozP8
XADbg/nqEewWeHuo8V1xux/UxWFmKFe6F850DbwJ/pEz41tBX/VrgulqhmkWKCFz
EUqmpI1Bbr/hij1vQ0hc1Tbp9LWc40xmRlQBzeldX9S1hmnnMh12BAK7egE3JDxD
LWxKlZalFgI9oqLeGUkkB17eq3Mecji0zA/OKkfTfiXyLEPbY/vi9SqwO01n2nYU
n9XeeR6conSyFgBmnxxP/sdnVsqc6CDwBXRv4RDa66L22rk9e+vQFTc9NYrShjz0
02yuj4Ue1KYH9k0oMWFhu7zS1Tb67c+amwGsFVdGQnzX2+R7UTZHiBo1s2KgCKl6
QhKMRUoPRpv5JvSfAsFjC3jWijkqEYo62MMJpCciVmrz/gmRj2JulhWN0IKyI00i
60kiwkD5ySVCJ9XeynRP0/iS7beT0SDlKiKRFWExAc5gNPGHpvwfWGoYgVeo/OpN
lYA6AFlGodOvqfHVpSSUhkL1xr+pbosoW224bl2mthA2lXOCrFiCbOU8/9msnsYo
FR8MDK7S3OLGtaWIHg8ekEHv92JC+zyCMFwXBX+KyW2myv+baIa6y2PoGI+o8JWt
CKsq2Vx2q2ZsGpXqXTohgpt9Ba5GfznWjIB7MXIrVKfz0yvIQwMfucAI2KaM3Z6W
GFEcCV726hc+eA2kMhVF2eDIPDEtifVPE5fuAuIazgQbXyUGTjN6Fjzig7BavRBQ
gKjcFsPTTZvLftSCio/bqoHAj0pwlm2bJLKullFFuyloBC50mve1fqDo6FrFC8/O
LtNS5UP6OBwYOKKWk0cgpCicF/V6McNHBpizNvNyectr/ssvOOHlJewRBM+oSyAP
rg8IXOarfC0BbbExJdeq7Wa2X0O6QdExjYvgprGT7ZQVKVziIXJjM5zkF1oNQOCq
/uLZWPbltJT0leT+u0fXEuSUxe5io1P5OupF/nBDZkFVYhRT+2wWLYgsbfkg9ry2
Maq46OLU0mzVbnWb4XjaTlxJLIvcyWabO3XEyo0s7udEpHCKxDAgqx4IOH00TBzD
gj67gWPKjJD4V+oKzbFRMsBY9HFbeRLYBnAwDKrRD2CfjpzicP+ZilJWYuACsqd+
bvNzG+fZtulmTySVsA0YZqoMXjzwJYzquhQ6lcjB4xPUDZe00GTDJ8Lq4SHoWYgH
8qHzM4eP1F7Q7G9O1hCqsbRh20FTeIa7mvRep1OzeUvc6bg0zG8MGLVzlBjIXpyz
648j9Ct/jZCvqezejlb/1SHoEF0K8Vzc45rJaCLzBhnZvZi+BwU9jKXm9OIdA/DC
7hev511EXHzFnMO565eIHYvOcV1Xq4lGrg/oIwNogtvSSElchdvrvwfW0R2nbSPz
ImBF2j/+oKN7giHW3/WVUCcMu8UHTtno0joq8hfz7B92ht0yRqS2tTNJmu6c5TXn
yhAaXzcICqfOVbWqxYHN3+k3Itikt1N+/Zsl9bIk2e7U75hhKhgL4+27IAuT1HAl
/OGWJwBEQ/gdTcL8qyk+yLpd2SQCI+PC43UA8ZmRuWzZPp6HXo3o5Yt0GLa308Xk
YqNJfCVw7GoVuFUIRTwbkm6lcYIl5Y0kzFHzCSu49D4RX5a6z7RBJz08Rs7pIEfa
r3Erh+MLqLesYduRJ/E0HBFf/V0wpV8jSNBPhu8kyPDskbT+LC37ssfXZuNf8NTM
0XlE6Znbyu8ar3uA9VRx+4hi5+oLioetTtEM7o7ESPd4JiutZ6L5TZ3r0hujAFDq
1J+MZOnt3C+L9W+cbVTgK1zpsFOuH65b11P23mK4sFpYHdWl/EX8Qp7PEJEHZ3qh
ylX1UCZ4wiCymkU49C6BfXP2Gwe1qB/yYX80CHLcHLVzlyIZyfA2gGF41KLJRNWX
roMP5aTIvu0nYqPA9fm54u0AR7/feJaRRxSPjspEp1HjD2I6XVHGr0cBnv0J9gL8
58x95NsCUd+knUPJAq+/nrCmcGBAMR4EzDHi9IL+UeV/t4pAb5zj9tOguqZQ33rD
HvJllkLhjxpLhITgAD5ulXAXm0KolRXPelPtbNmIbbja0EYwW/maqmnZUt92EtRB
mbZ1FGOg0E/2nUXiXO7dOB373x7pdF98lf6w6vERCvE2ACaPNLjMtmrWF/qJVjb/
dKmzlhxvUsj+xqJturPaDz9eB74ZTYvcqouv+boVuCAcGyrAUVk8OPzsrO2ZORAn
/by3mUGeVFuu1YcAKBa4MKVrR3BwFjUWXIa3efg5D7A3wlFTL6WCwTOk1lzIfPR+
arYAZtVErJFwSiAqoLvvB05hYcGMmsaB6nUmGjxpMd52obhOBW5wD+CYKMlQAliV
rCCzfSC4dUCISuMeGIcK3aAPQov69ymIsUXU7T/MCXs/gwKV+nPo5PKRj9odm9wj
LayTHn7sJaSJLkkZt46T80fCW0VbT6unKoZdVXxsiurlNGhQ3+9mbEiaxVGSxacG
/yQ69ZW9eij3dGgxZ13W2jW3g2AotlYuG/m8+3t4pcqN6JLiNERsT/CzlZbtntT5
KP3gUB8jmzXXW4Sqd6R+C4ZABf7iPTvP72h43UT7NJXDc+K0GL/YRRvpc6D5cwT1
4h8/1c6s1+taG7bSY00eRu5anK8yT49y9DjMcW0+9ThcQM7qVR+rYU5ecoXliitx
rqLrAqsJqSVSbVhiuM0TWRbhk3tlQjdWuOf+0Sxvcw805Y+ZyMNSpzlXEKPCY/HV
iDDNt0y3WbAGJYLJrK2xtuTzpGjsmEH8pQs5aSaPf/4kfhnZmQvWd4JVt+6KVC6C
LfZNWCBHrEdClg39dE6QUfDZvVilZuLa4PkdkH2jNvx2gUCoBp47W9XcyWbiqHiJ
cbozrPkQokHu0ndqtDKw/J3neTruiWkMf1U2snvCHVR6LM+R3Un759oRbtIBDH9g
6iVHnuhzrxujxUrBfvxkRpCn+vapZhR4iWa+tyWqjNNOtGx4+RVz6Y54SEptD19C
LUVQIvFeMXBobar90gz/VkmBWUGaHvVO7IrdYIYMsc/oHc8RspLMH9O+cbseq2rK
3kTkQnt1z36XhMDF7YjX7wE4FJRTP/biQyXHv1jkKNtj5Nsio8Y2aENLqem4SSaT
ZFhurO++niuAGQf1ZHS4C3P20WEvqwih21qGttLykpwzBFL2J5QSzXO4IKgoPARq
Snz3aW4PKqGxQB4Sm+UOb0RahXRua7sBD0gSU50i+1d8xPkl1pDkkuAf6eOftnbM
lCCT0fAMivGE6vnUO1YpdHDwR90nFSNc3O3/+7vFnEKo8AkiIDPUhPsyEC1QF7eH
awIsiCm0/hJee0JNQC/MJfmogjsjnBfzzMMqbo8eJX6+uRYCNAtUHlk6cD9nghUi
93XGtWc61y1NbZZk3+2o91Xpd4vPJnRK8/gb8qsrbtfypu6jAWjd8MO51RnU/Mq+
94IqB4erWcCLnBwXDZ4IkgjQz0rDUEXN22ZrDbsaTyr7/jOunIteLgu6wa1BOLxB
hKO3Vmhbe2KyMDIof5IjYtQO7DPexOyC62vpfV1x/Q1lHfrr4udenLw+jXWqbjT4
BPBjUVwAeY4be7xb6/rEEr3SOF58YfN3oPUYSYS34PuXg4NQixq/gxHGw4Vwt3sG
SKL+ZmmY0Tww2FZQFkNQCfb/wbYRCNnCi9yt63gkoVGasBuqCq6HmgYbW5m9k+vZ
8upfGYlTC1lHcwm1TAkJ1bhyXOPc4U8bJ5t/6LIMnvIYqxLsigCHsxWCx1Fk0UX9
gXToVSkPYUEAa/UXXY772uEiDjnn5kS/9tEHWrGb+5r/mNv9f+2f8u5ulsDGOS0j
roNkJR99+eJXsp69ghu4Hj3oStUhtyRb1iTPKSHiNuv+n6GYvj1X1nllGLn7n3KR
js067JXzZG7GaVM8nXeHUUekC0olDRpL8Oz5AzbR0zU/MBBosG0UTJaOAmh8/J0b
cs40LpHkju79Q+e4eXTuyg6wQsEyDHt7f92V71+vE0j/tBs+aLOusVWQZ5/JsR1t
eKFUocKXqZ5XjBEb3VKnrkA4U4L9uE3y5rJSQqM51TAeM4xlBwiKQrEmArslMHbO
1svyczXkwvN2ZKVc58WZbgeVulg92jV4rCbkG0abtFaeGwYv7wzzAt8hIC6zfSTF
ESmwKRlEe2StfP6mJIF8YraVYol6gOEGREVDIwvbAg4xGm9JVP4xaIGz/kS/KoPu
SblqrMedWPkRGup9EVaDzq1rcGolNlDD3UNxjTKUEeBRGFUKXKAC5Qh/KBGD0crv
nMx3UqBK0+thwasTTR7vbD4okXF+ct5+TiMXG4hVzCj2+N2iA6aV5FOAxhA8mZCh
jzBJ/49R2xz64XTmCtRwyZabvlm+bm2rOt6dIKtDF0zLyFpq059FRVpbEHllB9m9
fTkt28VK1igiaCb5RPLohFV7RBFEARqm2tcQ7W/wgRbLewlbjcZVVlpQmk69mz33
xsha310vkZ0AbMaulYeOUQ7HYW+So3zbQ6Z4tLbyWjf52ftgSE4VFpm8U4xtrk9l
LiABXfjositgowu2/VFg9DHuWFXoISXCybECjxWpAGTWCRMJC7hfq57BeBjpLJeJ
zAe3+4CxShiG1kxjsROj40g9BxKYbt45p6fbIh+VGGil1JqJexx039xYciZd+Wm1
Wdejg2Hb2+JfwOFDsqYGtWirGuYQOefNKUXA4MwlKKToNSGpfBOMhW4qljwpQwq5
poqWIYab2vufb4JIn6iAdJAL/kHjropTY9s3FjuOPJi0Fw7ES24CMtgGmw8w8cgF
Do8wXlDaVGu9juXxhQgWL2oQkqVrjmYEox5c1HQHEhbxfXYFE/aK5GKzuOIByXBR
/ixiXCM0KW6hYwN2hF2DBwitKxUL7gx+UBGAlu8plnSoBsI56g6HGh0Cn4l3gko8
1q80LSfqFlu3CmUm9eclnHS3JlSpvqTxqJf2gTf1kRAJhOE9cxmt9nac57I7VAFT
PhC7T9MIuA2v0p32ZaQ4nitF8L9KoUHBZlGFjSUCnoa3XeZvzj4QC4cFdiLFuwXs
PvB6AAKk/m64oFbKDk5oS4NL4WbwuNR6qsXMm35skwGcaHu/SlGEEbY+HdjU3Cst
ezBQQxDDGboob+LQnj4It04dRfWl+PtbcIVfYgKNvPGNII7/C1FycCm45Wo/fcM1
zQsgF/s5lPw3Nljf+EvU3Y1e05WST1mJlsrZNm1P91sYd+wilZnJAi1GeznOtme6
oQrazDUTeZ1h3NheeMghy3tUNyvanTYRRPMMnoLyPpIn2p6L9tzlp5cUR0AWS6V1
QdYYSzZJ3cTgE6fHy7itrPeJ2V5xwJeGb31SLgcyK4G0SHw/hHZUQmBn7LMLIV9o
8zrK9tGp8pS2CUIH5YO59VIlkf/N2ok1IYH5tf+Xx/Bf9kAit+aJXP36ddwp9BmY
LIBfxmUgbXQK5W/GXcsJtdDQLnvxyBkcfOcCcsVS5gEqYbj7PMgS+m1JZLqSio0V
hsBIYgKRoXSGZ8nL2lHLsOKrA82ViKJB8c61TVB9Ifipl6LYgL0oVXUtG1fu9hbX
vG1o9EvVXY5dW5fLyJa0BqC7L02PMdaZ9d5XjResdGxDiIi9OzhpaZbl/Z+siOcz
QrWglNaKy7pTGS4dttrOIcFoGlhkT2LhAlNHV25PKtCOkjuLfaHAErrz95dxqnHM
SQIV7bq9k1+F6zZw8HDNhK+zY87yHZf5xAXHr7oGzIhYUQHUoOWXovKREEyQLGHJ
fM5moYjvqECfIAsxT2xoSTS+6KEq4Rj0bDAKPhf2aKMysm/Y07VThOer7YZiuyXc
hsphRgieJe8s8BklmKHywE2Qi2vP16AJlEUwPJzbYTPXvZSHAofVUuRmal7IcdM1
oXSuKkQaMlQJbqhfv0Y5W8+jKeHrcGyt54ZAshRXC+PbthiI0JyqZqkjjZPe1KpW
AfMY28IDhCOiEwNum+W7fKGlCMU6igjvZX1pyIN6mCkL+UnOi2R/zGnKaA9mPcGp
XdW7Cxo4Ou4nIciCoZBFRM4KNSgWwu0ofNUeNhfmk6+Y9c8mSvPm54UDhok7dzc/
H9QYPhE0BiV+HwfAJTa3EGiCtoYwX1/RscKIr3Tm5nVx6vElx+ckQnpaoNmPypeL
9elBguKqEgi/wbZU2cG0lKk3wRw8BQQVEdmHm+9EI+HrU7Z+vWq8sCb/3cakNfMe
HIlq53ryFoktCMfIcTXV7b6JIu/HdF333mbGYdQpPbnViWXY+AwxOi3txbh0+jaI
WbaV96F4n/rcEtvnNYUbfwNPtmxSMS9wauCpBIvOXiTz1pCAXQ0PHZgOgHebLGiv
914X1yPzL0INw62FGcaLcNkIic1K2G8jLyfGCQaomq89MNbr94yUQ3SvNXJ2kgBm
BbJbsl1XV4TOZlKOdi5AROOtK1+YIrkmj3AohhMr9dUsJiYNUrePTesu9ZwgbbXe
4Qwr+yWKSuxTspD858v27Ra6Go/q9/J/rBZuSc0rJ7BzYPLjj2rAoe/imKfQmNd0
2rqFyI9FNuS2eGw29kz5RapVK4T9lhNg/I3kfq8cqu2t5R5D8+VuCt9JTvpRg/0H
2ays2aayMnLyiSfOzcGHORVCihlVMxhURz8qfTnJgYloaVSrjjLN6EGt5J7Btjie
d1mKMsxeY0k0Ar5dTNHzPFoJQOtyOt4hRqJeIwWIcOWmsMMEw9X5xFd8W+6Q5RWv
AzG/ypSfVjkBux/gGME38NUtq9zvjVlTwJpjNnszEdtTkMLbDZucWetOypLWV+Fg
3G+Gc7HLxh6I4PNRHzb8ykl96f8HUc4h3QgZGbpWDio+glbeU3Maakq5WwtANdNx
Rr6N1CEM6WpPsfJvqBizmRa9jyWozxbNdfBeTWn61NEzL5AKgrcltj4edPZp/mCv
hXhDpJJ9OCQQkem437Im4nxTDlshc81pH1C6KwAW+7qzT2M2yy/KeqlKsUrWoN0V
hGbdxZ/trArnxPRaGip0bdh9cOwTBoT5/TF1cAvbm1RxtbTh5IQlJNP6FssXwhA5
CkG7RZv+YUwp1ILIVI2HOK7OzCGq1Su0veX+VyprcfpP/BgUf8my31TiTOff10xn
+/9qeLR4b4xRMIuQpZQylqlOhk8kUwM3ezDzH7CgrvzgJIteflzX+G2aQitB57rd
gUh/Z0gyU2lchaUzk116Iy7qGsxcQh7cvy4hiUVmJjHvTcSS1VMXeLMZyn8Sn1h5
/u4NebJ64crNNbUW7QtPREuXqbmU1h9sy3WSgNxd1dggEmYGmYy1NHwB+/K6CalJ
WHhPtlOLjBuT3y7DbzUoMTNF/z3CkE2klDtO1/oLK7v/WwgO03mbX5iAJDt52bON
wnCDcxSAxGTOk0OauCIqtai+7GmUqdoFxcWEOnmopuTrl19nGITwTvah9tzYAiC9
vZx8Z+5A5oHmOiQdbGc7XYr9SqAMDuxSkbWzqUOcxT58Rah0XiavwrrhnByzRLHJ
1FSE00TJrTYghL8ZJBXxfocinJYMpZvFQAYMKTJ7xGxk+6x5fRM4wfwGZeP3c+mR
1tze+dGNatTenTul5yzomKzNxirGomCG/NwESQBdQSIGIgFttZkuoJ4ZqVb5U0GC
P/k5nCQVbxkKU4P+A+ma+AjaLjiwypZYNatCxOaffCD7njHzQ/kk/Rugjuk5RPsU
vQnbEsGVMhp58WqntPbI6AtFvl+2S55X8Z2bHSy9HicQHImWBxAEA62hWsfImRz9
pURCLz26kIICvUsKKUKVRZ66GKtopn1ffdd5mVH/qwxFs+HonzbJObQmhoDea64w
CyOw9hKuK6LAYjBpuVO+l2aHJq6Sax57vLkVSG0wHBJmAIvOlWMjxHV+mAFwggtL
uYe6D2PFon/6sw44eFUiDH/UyFWMR4KmopIHKjLStUdPVAe96B5SISvhDvGcCorU
ODNyscF/uXjA/PkCUt9lw05Agw30H9V8tKvZ3AOiaVnAVTW0Ek9ET0U7oHvLnuFU
WGQAPGMg0+CCF3N69Mjaf0I42cSWpAyEK+LINNgMK5BgFLQhpETzjODWxuD8+Kqx
QzkPxUycX3d35Mk/raWjA2TpB5DlSG/aZZQaoixovqR55fvudMIkWPw8TWBsX2qz
dQa3ytSluzzY6bBVIJkHD2FFCtymaUFwQ+NFbaqNkzSqkn3oX/eIOzczve5T2giF
jEt5MPiWwG4LKaUrkR8LDVODZOgfUxLntmJoa31S4Wlx7dsdb+uJIqRkWMC3McoR
H93Blw50CLVNKCc8qDl0vJAvlu/LYKGV49CgYIEI9nl+naPP9Ed9sGQr1WL3Im1b
UaM3j1ObPXPev38ORweHR0CAwEm8BI+/waGEYJVHu+0uXbpcHFCssGU6XvyhT+iH
hqsGtJ+sZEzXTj+U8uflqIf2rE9vA1C/RIGIG5/+5CBnnHun0Qkn5X+Rg4A3IWm4
Dnz2hatbY1QskAEOaSJCSHcE30758i9meXhkxn0V0W/2fx82+fQywtN8BtR/TyvQ
4N3CGF8Oyr33JlyDgupPsZW2V3NrNIqsuoXvo0oRDeywpM+uzNtI/Yr8mKZPP1q2
8Y7fJOmBnXOShxLNIOSUmyuk498kOVTUcnx/GbvWBM3BmH8wx9ixeXZwQTU0biLe
lRXTH3ZhMDgSAPLmdIJRtTNN9L+eb7RGIoEaWItNvU3MH+vswNpn+rwXsYLKLdXW
RDxZ/3DthveRFcgLXcn2DWEMwBrQWgC7+rJNLEkyXXQtTp/5ukRt9ywKJZQ82Voz
jnFyhjtKnPDRH1zOp8Rnj8oZzH4LdPHFcLkgRozMYiknE82ozG6llK8OkPDAAMLm
zZQ4Fm0qVH02shYDs2hmkVJTHZZcSZOuHCQoSQNt4jUHBqxOKSj1+5XP9G2AUHcP
qSU7gAfdMGvsfxQaZXw9La02GHhPKrZQyzYD4WgxPZwKhYuHjb7GcAszrxK3xfvg
/4VqvUlgWbi0nZPmUOS8BMJ2hApDEqt67MWrx8qI8KjlLRvFP9dUSEDwgB82IBOw
o9TdNRNhRY9QApjU0v0dBket48b0p3H/ADRyz7x1VNld1kD8/4IV+upDOXm2oT6l
4QKcTlfIT825A8n12y2lEEI7lcFXW7HMkFp74yIODwDiPebMf+srlmb9+dJMFlLG
kY+5HFmGXf+p2oj9s/3mgOBjFa2Y8HeaAWLy4tH4HPKl94prtlKUxGTmV2e1huyT
Y+YngF5owZAJ+kPb/dCwvUdmLKoyrwAVSjp7pq8dVO1vRW6yPkE7gYDnkZ6BYgrs
q673mab/iUVtbg3Fv830TmIy1jw8quhpmmyd46RbegjaZbn9W4VkUjjVSIMWZEGs
R83vHKJ5mhmj1k2GKZjN/Zx042MRv85Hx19+tydXVF87JBExaiVQUGUiWLfrIqMP
QvVQHNBHQef8MeVf7669aVNsDXdzQMmTi4Pu8JrlCsEaDdQCThzGa3AkmrBnQaGT
uViEs/vg3q8vnlq+kqTgT2TwdrZ6fR1jqsegxybExogoBP8qvkJl6Tf7pWsaTmae
DINd08LgXSromOmzckVhsarwowqdkbVX9GeOA6Aivg+jSAtYeJr3LUgUkq+oeM1C
3/vXfjKAwm7TN+JekAYmTuH7115wXrZaaDU+tQz/XHRQ6hIggp3aHW6LRdxV1f+2
J+tXlNaWJpScWvXG69vmLC7UOJ4jUVMKeZtOGUL0oT7KcbTTO2XW4hdq28bWNKvP
/BA0j9dapOvDcQXt3bJ78BV+zA1Kw1xQXycGQPVDWOiUiCZZJ/HEe+fXtV10eL8h
yWhlcmt1W4IX5B3F5ZUhDP4JVOifhXuoWnuSutZpvE5MeE2IZRiVTLXnJHp++oZc
QCaVO1jSq5+nIxWPbWJ3A5bkaik98Oywb2QX5Hr7NU/k/ssP+5Ze/xzgooApYVJw
n0NlduWF4+ARsgpy2cQHf2WZSDch+4rpdBBLb3mcFiHXxXr1n9d3Ie3WfMHuX6Pe
LZWSB0vPdEjrds24YCU/bpIMkyMpNPJuQrAKDipIXeFLZZ27f3XF+leA2kbVC9iK
SHhcwXvz1wxnIO/66df30Ez9C0lpAvFxLxdzzL8GQWHAE3SRRMQHw5XJfVwW6Xb0
nlCI+n5yEsvlAniYEgnYmbmVWyKHNmznyWbhKa1SvVXTAmixijHCcCwA/kJ54IUa
/xJbbxf0T3M8tgUNgOCz3Kw3bqm4OMu2vEzfTNEgYGQrD5D2PI2g/fuKzZj5K/Ab
BeEwLSV9gGXqeEgi+a61P2bgUZ67xzD+8vLEyM88kWq2TTqDqOJ5HI5Moo5OxT/c
+LCzxYeZq5WcS+6XygPQ6+550LoaNbB/PWP0yGta1uyJR5ULJcjMs+VhL8Qqt59t
JRrSnX8ZOSiYpOsTTJYcVRK5U6ueTZVlyuQryOvma4eHHnYD/UVp8V+FyV+RKhzA
RurZ6G6ji6hLGTWBRe7HUow9itJ2Cp9LoPKV+kl56OQY9JoiIlAjJHprTsZg252d
bsJvQqchVgxec01vlKECwMeb4Uoq50T9SvI2+PYh6u/dzhVa4t3ihNLTv7Y6LFwj
dKvOvH/tAopSJ72Sif2NuMxq1ftAj+X5W/Gw3eDZN62QnqPiTfj1gG2Y5lR4ddYT
VKO4F2VfRNb3s6yzWJxBvhILPbSutCby6xcL9dJGYccGFefa4QMZvfXZKGbV19Jc
mY40VbnhUhxMc240dLPFhx5dQbbwRmkquA2+vgy6/s/pR+u9MN8bilw0p1EzaW3P
W21+pSPdJvhYmhA+xxQKikRj5RVjV7gdNWGrmibCx2sfklz0IyHDzJtUb6CGatWs
MGM96wpP3sSfLOHF71IXXVykshZyk1PfRWSluaNx71/eNpKDreY9OUU2n15COQrn
qERr4uH1hDWk1F1SfNzz2H0WzrC0MbP2cVoQjcpVCzQhdfZ561U87tCFLgVCriL1
bYkTBCxrlPubnEQ8QSXMQKZykM9BuCmEujznYrrt/n8iAWbtXhsWT+6hinCdN5Ay
CqWoBnInO4TduLVwrtE0FXPJj6StBq28Mh92lk+JGZPP3zSV/2MlBsBnwGP0kAe6
LzPFXVXHArwnSMyHmgqmCf6icbg+Z9doMamiEfQ7crGnsXt/d0vvbUqqpyYthiUe
AKShSaSkAiMrSVt8UmgoyGtpqbFg3O3jvNZ2vleLcptdyiqVERxPPT/dU6QnaNYr
LqbWekJbDAMsvRETqVhMor1ruhq+DNw2EgJ6CPbHQQxfqLzTBmDexghnmW/jRFsV
JHO3oewsla58GdvaRgwkmagrKcfnJUIJKMEig/+PG+qBkqlq6/EMHGsFPMNaEdVh
lRWV3v0A4THN+Wl8dgXjMl5v6kDKzCb7kL7+f+FEWy1AfBohwCxcr9DVV8TbWcWA
f6Im6MnVNQW81kbRSRowRzRWLe+ny60z4Znomeyj7RiagRc74CbzHoZq9CeQ1lZ9
54By2MY/z4TOlOPsoQbBs6g/nU2f8NVdFgPBouwKrMX0PP1VWfy1W/U9rjGGglPZ
lU3MhHt7rGnb56sASaG6z4cluA8nZ8FbkAf/mPYSo4DH6pP8/9LgAQ0DyQca2kxS
gwoW8+A+26OUVd7Ap2sWc9suErG81e4yosuWz69iIBWXguGkhp1Gj4tEVtm/K5p4
7zo7nhdQNaNrLmPBjQBfr9wNf6WyZF0a9jyVf52jZFPW+ZRQACWwc8Q813Fn1qRk
xZm6KaiV4DIZdZtFcpclg0DDyfBv51o0Qi8ncihxFwbvswO3sT+THSegS3CedWG0
2tsnj8SG6ALksIw16srk0vFxl4Ku84T9aM4ZX3e03tgMjBusBSSy0/q5Tc1TXuYy
cG66fqMaB85BsYeZnP0esnouTg+60rsjvtm0gW6N0PjtTBS4Logg+y0cAds1eW0V
77/mZim9bEj6sZl/pxg2yf5F4EoPU273hAlUZhSlsKVVQ+0TCjPIOae7+P61JmUd
zDr/pljrBLoKpyzcMSgnOtlbtatzNxd5Q06qZm+OspRYb8DYKA/thkd/da6XiLg0
Ntd8BzkC3hKiuKGqDd5z+sGDNjIqxCa8PSBUE2vI1bZ9vmg6ofongfwz82q/Yp1E
2XSPwNkofWUI/LoRwqlN+PiZ5idEN4kT2Y7xZoZCFMShzn0kfHpMN+uQltoa0dqF
T8kQBXgB5ylybiN45juSrneDM6uWClpZip0M8as+d/+hu9Dw2Gdl8OhLnmcCfgEn
RA4RYxdMA1JAZ3xabGNT7vzNmjanqq0FZxFe1lsnhtVhG9MsEDM1sw0iffpU4i55
fMc0iukbwQRWjuffYGTyOtCFUArtU21i4kH+IUrYd9NNzUYH8xfS3nR+cvjlOOlc
L2cyGwP3FvVFI7PgXBY5B+zkgtOMHhZuzFGVoNuzso3U5D/lPGSHRVIQ4gc8WGNr
E8uXo8Exr9MaF7lv1+k42+EMJ+YdS0rIFTJ4P/vbHYcUH+GRtxHJndg9rw75NfsY
d7qLQlc6fchbfLbG4OgsZRQY/kwqNPX1idY29wyE7W+hkStJZ+ADdUxFbETdqvZ2
r14mS/7lezCGp8fSgCpo1tLnsYzrlvcOVWYoIp2MxxcBj/R7847LGwhbFX5cpSne
E6QMhbjs2r1uSUo3+aM2mld8e+jSEzjzF+wpg9qloZRYBIxYyAKEvGQR9qHoRbax
uYsGxVPAX3qtH2uX6/OjEqNC/4C/j4ZLMg3onwcWwXsoQJS95aIQCsOEvLpg8wxm
8aIM0cM576ZbqHC3uLwiTZ6DzTJ+qA2otQ2qnDBY44BNffWl3zqxfY87/DGhRhkn
GtnL1fZ4QdXNJoet0pH4zrMpgzXwy+kJ3QeEwgpOmmin/ULXkrj/WQhIP5sAe5Xd
SL+3o014nfVvkRqSnMh0Fq/2itC0PPS3NTo4jNR6tKdOYkVBb8rdQfAju2qDUnR9
5X1kXlTXoxZV854R5jTAC3nY9o2ME2B5MOYThBHaoQdEgrNQZrFKNA56pTfp0qAz
WPcj/rJTgAA/F2Jtz+yx/TTtDDWK9jVIR5Y/znb1/Xn3xxEtgd3+80qbGWCXlDuO
w8Iz51PZk8rmdCbnIlX/roLbr/5Fq6e8Oa5lNfzvCtaxG7UjFBzXOcYdiro+Gwej
PL23dWdweFyLRo2nXCZtgZ5KHgCWcIfaY1jdRs4venJXwdi6gWSyBeN9rikrjLZT
luUiELBOx+SjgDejkxUIUqaP/NeYKIQ4rhPPdvvvqb62FtMVA7lpMwP7ZN2Avdbj
vfafhRI+tmhCQXdnbMImi7K+s4+Sb0EmuZPC6rPO7HbedGDsDJ+4YucRPfFIGMng
6drWSDDKeFqiAM61/fvuTMO14faHlIOPV0JlUrBfsWNPvxTM3adOy3HVBcVDwUsy
Mx8d6h3RcLXnUDw+ECT92XXGQmcXj2r8CxSJxpFQrght1Xm/8BaNHEXbjarmJTOw
H4fCBSorHZrJ6jKdVkxuYr8VXasSoBLx8lf1O2YyNq6rNSRKQjvwp6Ux8Z4msRoh
coteX3+rniqXxpmM7jAVH8Av41olJJjmsIyNmTE6zUzqm8N0VfFhX3yd6qzGnAEE
dyv65tDAuKMzyHjpMlSSqWPIPeswCDij6leN0EwodCLfBcvZmBO+ZUntTKray0sL
yU0fLXPi4dR3nhEzJfn8jeHGjsat/R80rrUREMRmK3vkOZOe+1yBRspYUHbuz0El
UMcMuXCzeW2XGt0SpXB5pnTjYxQxGBeRXM7Q3Ux7vF1TYdyKC18TogWLACZ7GDNj
O9R5r5VSKmtiOL5FZn+2FxNyv6KZeUPVqKHOj1pUXIdN6mJ+Fdn9Q6oChhxXWZRs
x/diJ1Gz5/5Z4bp0otMfa7Cy4izR3fmW9z9fPSoyXG1MAQWpeaKbtyneYYe7vj39
uUwPHhhvCQ/UuAfx02YlqYeznijJ4VFlU8XCkiC3273E8JaHEfVyWZB7MLZF8UA9
7+oySIDLv8QulvyF0gw171AT1uLJxcCl/hBB7Rd9gWHfTx8qLYRRivuv3wyf+wfJ
2Kh2TCfVhVKVITNv0AcxLv0TjCXlfDgy9sJKtQ9yM8vMD5EJW/Yv5njE960XaIi8
Udt3/0/ECm2ReMqriNffg5RABG9rMxEc/xT1boII4+NDGY3OyPMwGcGzkIJ47j3F
+twp7t5evkkA8H2IP5NK9/5theiMyRb9CjVYGpD+nGhQUiz0w1fgnQSZR+OgvZ9A
ErydlDB5/jbChcRLWj1S7Abfs7TXx94NpWOUw4ca0KVcL8QkeNL0XNyFHZRUwCyz
ZNKmTwAPG87GxtsqoY8y6o7WsOmsxexO5uxAgwbztpe3ko0v2DCAylwdOPxAWdEb
Eg8l1oCHqGIyjZCRbWVwOKzM65YQBz0LPJZRz9uyQU6g6cYPZ7aIdiLJukUGjblp
PqytLGDNL9XdsOG3j/hH11Ybuv1GvmWoSUhhMmmLeN54v0BteEBgAu//a8qCwYeG
jQUUW/pzDtA95R99C3x5BNQBJRS3YG162+mBEbQDBtWvI4Bs568uvOl9BjvhS4Pn
VslU4AhFeX9Euz6KNKRNcHRsfQ+TSzmdetjymmLLD9UO9EgQcC7JKx/X1DwxEbCo
1aKJie9l3iae3l1sawUsQ6HmCXyqUm1jKu3HXZgw4sCnX+vQFkVLX5zIb8hbBozq
XTxTraySLma+sdGAb3gkjl+Hf3RnWM724SMkV0fJ1+x/PCZCX9kw+jCd+STGdEyY
W3i4BF35yjOrabWz2/DzDE3zqwbvlHGcm3Q2s+fNYYYOaMda09HIswjn4Q5F/t9/
+o1cGtEzTVZ48YQIqvlCXQHNIeYiXvyb8XUkUS5s6To6HGXgP8hkwlXnUl3L1OVD
vN6MiP0L4uX/8aaJOI8mraylYlgXxIBgZsJw9dxEaNn9sAi8iUniejvDFW7cDE5U
W62p9qgKr4+yJqTx9HUnpRnl8i5MjeYfdQCGa1tljTQvie0lmmKfkaaQJFzolOJY
tx4y61INpaKx1oGi/EYFjB5BjOhk44+gcNfjzti0QuYAvD0lHbpn+7JJHOAxzqRk
C3UgckbhtHVRpphQUYsWSt6f5u2I7qsTMKsa+2zGnGZl4rCoMzdci49viATQENUA
WyGc4+lWD8grWbMubfVucPR7chfq+2wfN6ORbNbnZ9UwcYvrkVH1o/TdjA+m6yD+
e0OamZu3xKZvdwg7bsTX+pNU79YnmlxK42ccrNzsKqXuJ+S7135XB/VLcJ2Ht8Lj
1/9QG1owz6yAlwbMdAvAmUGYZcEVw0R7nd9Yu2W9iqzTNUjlihFPjP5lSXW6h8KE
vkc63EY15Y7qfW/6a361/8XD8bACp9W7C4CFg/NMXx+sF1luKIqvoi72TjSogImE
C8X12373wjQO0bkz6jD/x3PHJ8YV0ZXK83zr4X6qQldZ0Ogs6Gvpj0qo0g75665O
sZgXIjdc7oFt2H56rdXkThlDBE9iFHKoFmgdK67IneDxqk6pKy4ifVf1H1bpSGpt
lhetmWIJSoBkifwmfkZkXtsvRT0mBxCmvjxywCUrm4jP1Qp2v724IuAPeTw4wg5l
p/6XWFxrH9z3z044XEaHzh6ujozthQbob/aBiYaOVVvgsaj63uH51dEXbeIqq9iC
yO2z3oj+RNTMmM8yLxgee1ogY8x1nQhiAfMY7Mqieq/KlVZWaSwk27u28cbg7g3w
UwTKrMHAfzI+MGiez3YiMual+yMviWqpQ6fz0CiSc3vZ2iIvpqodJc5Ef2QuC1I/
E4W4JjCCqnRze+HaC9gmIxihqy/FxA9jAevqqLZaiqzuSOQbLH1evShdjmb0m7NY
X3J65TRsUAJkzhjvZTB7Vnc1s0CggRsqfiEOuxnpsUWDdUQDr0n9JKM735DIGxRn
c3nQRkubyz7DDgfol97yRy1AfdyUqXViNx73Z760J+5V2V56Hq0kQI7ng0B2MF6L
iYx803C6sxOdUGu2v89xTMF+En6e6Z/6+cywFBGhw4dMrLFsHkVKo5dSmQ7XdSPP
WV4UBhKwD7cxTPM6uZJebXX11zyu7elNHVgJ1mULfwplk4WAMOmDsf0eVTyf2ssK
Al8fbiuYldEV0pjwVdNy1TlfSVCDEkmIK5RUuC/ondBpS/7EWamjWJcooNlSOPCo
w4qF/GcJ/YqdRh78nZEQqsM8fk2hA5rlKtNghM7NEo6Y1a6xO2ypJ2wK08WCAIA2
aO2i2avlM6ucq5A6UqTWab8K9pUOxSszThaYacRk53TSKskB+RhugTnrRf7/jca8
Cw+DwavtAbIiLAVLp4uxfBXB3+gYWufWyI9nrRnyMnPqDqBXSuXjFWi61DCfG9Bk
pfNeOAVID5W+Y8gwsnQC0iIM83I0kQeQD9jc9oX5H8oBP9SN6s0Xg01JX4fazoqi
vPrTMFUaOhFx0lL3OfwPVSZfkkmP4qJNUBZEZs3R1/ve4uJ9yR3DzCFK7bigywBY
A3Gh0IB+pUfJqEfj8dKKs9BCopAQ5BsGhSTOFynODD0rSFUcwRCKoGGcSH+ppD7B
78jtsHrSFqCS7Dl249XiY3C2Iczs4RlN2ySe3tC2uiV3TCN+NLVAZiTwGpddfmm3
EYvioGjAoLYLdMTRnSNn0hQI6z8jitiLDMV8PEpnrZ4o1OClAfPLa5EJTAJVzm01
g7dUViZIq7e5W0N/rFbAcEtGGNCpnfAZcaesnrjoxzazR0NYXjV2UhMZNM8YiCq+
CzVJPhd+zA4MFeOAhkGBysD3yzhjxgW41l6YgUYdSw27I+UnLw/nYveQIbYAN0pp
+5Nzmw75cs1b4UH7gOiVNGXMMDj/x6o4Zf2u65jRzjre8o6qT/e81YF1IiB65eZR
ZTBR62K2odUgxK58ElVJ1AMYqtSxrzXdzMsbQslYiKAhh4f4Cv+t/aznsjSyRdJm
MJ9k7Umqoc3fWXVhnvWJMPpUWRFU2A6UbFJNcwQ8G8Sz51FVpdg6GBNxN/Xb3LRO
0v6AFUvVeWA1VfbBdowHwwV12816e5OSphHOyz4PVrGQqRYOmAdikSLhPTo3QQZ0
6BBcTPV9yNf+p2iyNLDuPRRj0Zg1CKKgh+6PpO+3bB9XcDtbVjDBJ8yj5fmOv2M+
CA85ABrtk2QCEynP+aqgmbTSm0KKmhxvLm7eQXLq9xLt5fBfotFg+Ud7n73K/1Rk
YRnPmjFEgwaj1qnBlz7hbjsOiouKRGcA/E8wmGvJpZ1rlXCnRMq68x0UA2m6/wDN
fbYKCIk2xN/U7fMxY932KgqsypwSg2Owj5zbPtWvzLtbExIW5STjQFrSYKQouXkA
utMIHxKdMHa6sN5x6YlzQbYGolDjlihFG20ZC8XLUY9FpC5qYrYfasuXMpny9rLK
zjaUwGTD+qz3kZyexs14iemVBsqJYpfwC8ip3BOf2j03pnnVhLv0QVlqDwcArOev
C7DHAyHHayPxoncFy5dPCMEA2wQUh5+egW9Ibi/iasitEV20vRGO5VXHgFzgFXP2
eFUFmJF6KOIo2EsIw6GIs+tOlsotmRm6Fe8bVYwIaxuqLvGuIJCYqlDCv67/sUi2
0yjsTnKfaJXOp+c9sE93UOaUdCxYVY2MjJqe5KZFARu2V710Pkzi1LoAcyxn2Ccu
CWxwJy4CGIvgPp5jQVF+3tXbPX3Lh8EyAqFgDtB50JjUzVvwJuB2luXX1CcmWEw6
NwD3jJL9QVBynCsdROcqM0JhKPBCyBCpqoq1sizp4R30doB7Lg4vzLMJtGZFRmlM
PINjN5/G8/UNuxuhnNMxnAc0r63qaWb33vK7R/MSyK5pg+/+DaTmDgRN7TFI+2ts
Qzc0wIguVr0jVkHEpkSbRWWGiqayne6MjdcHjMHqp92SBbWCs9y8R81mUgd7/W5c
NXd5i6kGkM5Qcpgr1oIYtEJAAgrxO5b9cJSGes1qNgklyw6hJG9VJFV2RZKpapkK
lXCsqpjI8yRvAGHt+jXpCuv+RFIbXozXoYr5k91lr/7PlugSr1TkPee5mht/CTZ1
XCmFNEJ+CLomkZuqMVwx/vgQRGkJEhNkV3wabe2zaRE/Sa2D2XMHQsqDTMmMT6xn
DyBU0ZI5NzXyWXH09k3SdwjgNngJqlDqWzwHWTPtmJCHGUKIYTvhl3/VTexmGXXC
unWlt/BiGUIpLhyVAoLRejSLsB9TbZ0jW35qmLCNCwVW1UFcAxSizbh+hwDqWjEF
m0IZPDXKlCDeKZ/5sz6WFYAr25dYMIZYqz1obcs0OGg2ImzONiX3JUBFQAvVKBO2
J0MG0o9ZBxWlPucS+Pe4TKJJb8llUrzhV1yotQpz2fSAylQHAZeQ/znKaJqgZD/r
f1KkcKxZPQ5MEx7bICDUErVgurVij/z7GNcPXPcb3sVU10KtzqPy6MoqMeYu3XTi
jW16K0cUaGOHTCbaB971URbbSxU6pGKUewLjYo0PpDinbKmG7MRmk77Dwg5ntPbH
Fc+lqUGA8aisyIQajsYsTl7CakkyedaYduzlR/nOXT5s+hAVrEy3HLO1NYKHF4pz
7JO6Dg4FzotvHI5uxleTaxXawKmwMV12d4W9egD/vEZR/5+0YYJfqX5atMYL8JKK
JqDsDc67sDNxhijVX2KMmiUCXRIOm20fclxK6WawwCsxkCrn3Ylyr2J89M+m90Gb
e1QsV3l2fMOd0fSRxBoD4C70n9BAH4qT0UaN92XyQP65H+HFpCr7r5cTylhwqW4a
sYz4IuQkoL+9y1wYqkB/CkgraLwtwYlBCJP8reFEMJIVs+01oaIp4r5IsGEjvPmj
MtBdd5arLkW01p69l69S4rWNDzdKNsNSbbg0KjPoQAm06WR3MrlVHzhTN9OzjrsZ
uO/ARNzpux8jYonKHvcBWq8+JCzrHxavYbByTC1HvT7yVdx6clnxLK0B+xPySByL
txU2gmDCXnc7ZgT2WImbKIjgEZd/Cg05fPWvVHMMKNMsOKdBS5MGkNIUUcqcRj/9
GYRE7/dBxdxTpAdq/M9oJLZTunZ6RGXN/bcw8hPwmeC20coO5AP8y6Y1aDb0Pb6H
GaF/2J8ofFPCFm6DPPWA40X1M1Z0UbYEyq8eHVwOQ2ZJSEnLtEpyoo65pq3WmiNd
syrGOmY3Czw6SPrL7lfJ8vU0VoMwgX4eDmv374h04hTsG4sN0yLgptxI7ZRoSSNI
cJGThM+ydBsY979O0rE6RRg0yKTCRHhyj8gBcmQ32h6en9oLne6uhOaQuqENyoAk
SXjbRsjTvNv3kTNB0j7DVzdH6ac3HUyB21KFMh/8TCOM0RZkcJJ6qYQEKHG99F3Z
xzv9Yskv5HfEw9Pb9IxYTAkRHwPdzlYQPLIaPSj2ozzlPRXQ29oa871073lH3Hj4
pCjc1smnfMwyYh4Ir7EnNgjUwT9einVC3pBg3ATQmr91DKcqnbARgRBLAA6fFPb/
N63pbQS39pbJ8TBiiLWRpY3g6YKY5BkTU9ElR5XQBCFwySyjWILsgt/q6YgSDfQ+
9B0sbJVCpxw95fIbSiKFRR2jyQiVYHhW4LwyHI3cWo/bKFQc2facCdBhvD2BBSOy
LYoBkFvsV4QPURG5vDoszXz72zR5jEauibhvx0mimxeSCdywgim3oVGH7N9HDyp+
b+T9r6h4oLF+U3AV2KzuibuEqNcR5aS9pehmhGux25FOCKMN3s2CWmfIy+TP3dKB
B5SwBc+k1r4oCkG9rb+Y+amJdVI1MFIZAion4l1/q+eLClzOLsNE5FVOxSqVU0p4
86syhcrAXEfP9Hcw0J9yeBCiWyb5kGdaSmLs5zK8j0csLPCnVTjzVZIbQdnK+kyj
XCFca5biNx+J/5MIzdidB6FGmX0iq8l+0SwTSWBkMFH5zsJmrpTe3Njdzj2NjkCf
4lWQM72VvOHq/wOu9vco0eCwILIiNFchZvsGnCHyRDBDNfe57XRGR9k92c5ZByZu
OFkPD7kxjl2/6DmsljvRlOKbVf9b48tikPD4HDoykJ5oo86fE1GwtEYZMj6Se74g
YTVLMfQoipYmziLEr70Zt4DE2v720GHVtR+tXUKsTUlFTGl9wQ5bajiQKOOT5lag
7F5WVSdvYn5hfgLWU8Ow7BaMVrn4tUCuzx6D02EQSnYUgL6PWlbz4O10mFxtmD9R
gQ/6EWSXRluohHqTK4EtvynMogWkpXQxXvxpI8w+4KOORADv8MaOLFirGrTi3OkZ
kqRx0c6pDz5fvahAX+JU3rQ+V8r942xXQCkUUZNqP4oxPnZNOgbYcnJfsBMV7+at
dlt//M5QeFX4LRgd7fiubrrAfNUjkPDrgZb3t7srnapaPy9PJL0wVon6cF45zRt+
FP3XJBnbqZJrLqcibSx3K62K3AE4WtQbBA0w2tNP1Gx6u8lxiOizlpao0/+O4l0X
o7OUUIPmdTQO4en9UIGbeJPWbV2sRJnMYOlicGpBKXnn8IDEwVfvRJtLZpcwdFYw
jSt/toAOUtZob2RR+EjdrvTS35JEeEg5zgA64lxlr+lB/GALlWMyoey//5MrFb+P
rowSuhN7WETwaNgX0kyhou6bebpNWzGsAjghW0qbXYWXqqRXQ3X9wVz4MR3Ag4Ib
8JHAD4BJwQCmkaCzVw9A1H3PSXv0IDMD7bCOIbYdh0c273o3WK3HtHSwLVB+UAX0
WMPjyLUhYi5+o2XQ7h5p1GFy3rOSnQx/+FI8RzlgIAEH8ulQXxmHBvSb9+sBuw1t
bAavmVlr7ELOmoDegGiNy3JqzM1cmtCiF+Nn5YXQisZcL4EyHmk6dtii15k9WgLa
B4337OyjZ+RGPKt70p6vrBc5aQcqnjMxDvDFOznGSqFE6lCLjOwY/q6J1dBYwtu2
Qub3r4Lw+3qRKHPSQFySpD2BzvyEu12fUf6+a57sFCbKFTURCqKBXWMRxc4KlS18
NaUxeqw/sUgUDAyVgljT3h0Iyco7jBN/yvYxW1MHORqbXI6zYwvCd9zbDjOVKEYl
rhv7K7KAlNbnlLwXAjR62uOiM7ClHv50Ck8WJo6bG3iIoV3biSFMDewtoE2nKIvh
fqRRPdvafY+qxDnkjXD7oI8irpxd9bmEt/YFG3L32bkP+vXrW58+f/GtHdlv04ze
Qq/ActhUEqzsbOf6DQjfWip2RaaiCpfQRNNFcfmwKhjDMelsMGePMPbFpyC0FBnN
z71QwxDYkR7gDcW/wqZL8mttoVRvNpYFW9L7vAI9xMqnNjZM4ErvB/h1SqEgnyys
efAl0flUw+dF1Xh34xltIxECNB0+N90NwUxXBjhD7W6hvW6hpxmi719j2PxRmp0X
3KH1v+ldQWikl+WK5Lny071yMwZpuy1xGshnifeBGxhyzacvDjjEleQUsJXjSIfE
ygOHG56qzf21rdixDvDYG19bwYUMTL11Q66Y0YZ0Qa/JouyVUPDvgzK5RXTujXFa
u+kzHT19z2KwS2CNi1FJDDFhSvf1ghuFjI8WJDOLc4lCLTMWxglhqzHOqOpKMFy4
ti+j1RqHs6PesIzWYdhhXboinB11IvlSoNRibxSYVTVtkHlbgXNUe5OUSdzabOJ7
FQCpMK0furVf592AelgasBtor7G0T7p8PNfB1dtuix4R+fYrCuT4mVZLGK0Wvu9y
Wg0Gj6CPDcr7wSaDLV2TdVwBd92/vr4OJ0mvlZa6aB+E9Rd1mcDL4AutOrHQm/Y3
6GzC4uYFdlxa/C/ruuWYU/J7pIYCA0FdSQfI69BU5TbaJaktijGGccBpG4vZbT23
sWgOdOycR+ZSvwc4+z4TiRTGdWADFl/gZBDkwOtXB3h1lWHccvI2Ku1TFsaFi3+M
pCeu6VB2Q23aTTgfQdXuRKEa17sF2cIP/0F11bIsTYX566NIcZHZVghXnxyaiZmO
nTYW+fU1YhaHCaFOIPfuqzkbVDrp+Ga2nWMHWODMWa0D96CkFqlRWaky3CWP14Fj
GpKzb+b5v9jCVWu3+ke1cDOZUZZlWbymlVXq55Mk/U5nzW++c+l8648b6fAoN+Uu
jCCD4d2yYw8aU4nKjOCCXqFOWAppe3uHAZfZnnSsX5r7FJWGu8d+TlnycCw4jSCn
N9zsuk8nMAFes07d2HQfAw9vArlig5c9j7C8Zi4woPVO0DUzmsAHbEXwuJKdOYW8
hnLaG+g5DWeQz1dCDASAbK21Xpl89Sc2HRB0RUfcQCtp1IVGXhRAGOL7erpnKvmH
ZK5QpXg7PPfzi34esbhvpFHWwQdhFyikI8+DXQ8neShdovy4r4bviRXv4zNKJIpW
lirDoWWmyNsRbsiaGTjbPnyVx4PrJAUn3TFN1OrENNWEkxfoL2TuA4Q/qPLY7nYi
D9syXTRclXgMRJP6vbfC8urr93q8XoMBBEww1F80CbdLB9Rj9iKH08qOtQ7WZ6gA
emy5x9HRU9N+ZUOs+9ye78Od7r6TDAZqVZgQfbZahNJL9t/Pa8ijRylzD6HdS6al
omfeOnLVwjqxDJHvAk6HarFQcTnmzSwJdUPMjKzoiYPrCPfbRC/uGfDxNxJGpVEP
dC9c9keYSq7dPJC0k3iJmPT5YN1iy63NhtrJEd8iN333LJ8J7jCy2i82pJJUW5U0
sF/gf50UK0u8JaeTvqjHWKVDHVt7BWm/2+yd2ylH9/7D7rpkJuVcfBRtQf4ea/h/
qK0YJ0CywB4FD8W2y4E1D/rPD7v+BYxr+sdpkvIzBpO6vgvfvgESS4R2l0ef2tXa
JH8Ya0PfX0MjfXqBRu1jKx6pQDYqdzzxVbtnOG2ZieXjq9toB90UHm3O6wT0tfsd
qPxxdvTaLq7QXYzHI0+b4hICTXrNIeclzA0ivHvULM2pz+Ez5pkxrDchZMrLqKg8
JWvzBmNjQL8rMi9nvV1GMwzzV3F0cQAIRMRQ4Z5z/6cc1N5DN+uAIeUjpSh5yRKy
PcPJ35pvZrm38EHjtNfaCGpFyJMmgi8RFMbgJ5NDlicUPEgm1ApbrFPrTLdwFPGP
4MajCZHf2ADe+wnnIiBbsORwrbkFOe9eSCqlEjVVuN5usfn/4JNH7T2rJsKa7VIo
guz8XFUzmaSWUbtmrQ9dz13bzo10bavw97/9mhlZ9RJ4GiFfyzYmfrKjFUlczEWy
3hXAm+xJ4zGlByRafbr+8ZVwwHi+fI4wysw2otpsTjiPYpZaZg2ch46uPF7qzyA9
oZw1gEJCYx8NYU+ImvS0VjpveZx6lroJgxsHBv4z6cF742BDwYe8/BOwJn0c5X8n
5Zi3QtPW/2IR5SlmXVGPOXwaGoPXBEL4/nwQtuQQl66lYMVbYU1q8wo0rIJSyIAe
7jamrcHvUKDP6/J4vOTiElNKye3rrkt2u0rk5jJ7RpEcjdKw3ED8Sj983xlJ65v+
/qiDCLMFSkI5g5ACBnaqR0XN1t/8LVdY3y2JOV9xKRGWcTZH3fBV7AxIIzhtzjn8
aIX4OHizBONx/WpOYs5iDUci2ioEfv4B54camUOfQfAgPXy7xMvFp/kup/EDPySu
R59lBEyM+DV2fHpNuS7vj72KBkkQNApXebopu6hfy2s9OpRwxfnYeiKdE1FiUgEp
O/VnZVMOLpecARylusthr+DKS1Njz7LCryPA3f5pwDsRIovBJkQQgzZ0Wd6JP+9L
gn6gOYHC65PwSjs861ZvD9dAQwWJ9fPtk5jU0pKyPQuRYr2hRnTu1ZJAqj8SdHD7
QCDbZ4Ix5gZ7ro+QGuDqZhiw0Jb6I31uvGvWudHlchetoZ2PFS2vBHhK/bcmPYwb
XAUD8X51dx0qEuwiic/rMnyeCHDHPxQkcEuIUUmut7jhXnuN1XYZfGF0hodJ74xz
hjX+CAXq6gYf5OWTwaHZG6hPnFlt+E3/HlnSqGVxSI+ILNUV4J9dx4etFSc3llsP
Pz62F2Nk7IHJAwdQq2OgrkYXnFrRnh6aocdKJekrwPyvj3Mxlfi51jetNhBOiaBF
vUAd5Ym3SY+RHK1y2eI0sjYLQUbLCyfxeQy9hZNlxy23FZC+EBkxqmQXyM9DAMaf
IOLhHnUHvxDScqGHh3AAsJPkFvD90ja612/18gT8oVPh0JnAkB+Y1Q2THP152zp4
sF/G1HcLoHExRqE2a8QBvVODwoZT5YMI3X/7hX1CsVpVk65oPkg53FWc32/Q1s7Z
yZfMarYbvSUSmBfea42TLyOffIBt4DBvJqcuy7ewFzcA0UxqwMOp4bDb4knGCH/+
dvWnABv21UcHZbdFPqo6AJaDWHXogAzqGbflFmvLgVgFk5feSTEdkkKe5zz3Qnb+
Qvb60wh4mjYUZVmBwb16GuAOmeZHgYHGEArIPbAMvrQotUy3a3mWsgdqCkBM46ce
VctDO+tO9X6O6FTg4wyptl0pu5OZTmyU7nQZxxWBfWRoR6F8CyTYeuc/ruBJOFOg
kBCTahUdppEb8YLO63LoLq6XPU4tG3XN34y7sGNPQsZ4OxCkjVG/hC8nndzzIayP
esDbd2JBx1ncC3klsWnW+WoWb6VB8thxjjvHOlmCZ0We6nZbVgKh+n7G6ctDNReb
fsBSactPelziAKDoi000JshZKZzPxeaEBDhGPjJqodcXam7kW+/OCNiVLFdIhrvK
NbDFPbIlkPWC33IiYbzZli2kKlY84KZzmijBL8G5mqi0F0oJcky0HopIO2sFVS6Z
sIFyBF0xQI6oGMeJ/7PDDi/PD9sXuF7jC8ZV/0nPwm4nxEgtkVmouWPCfxtSGS+p
hbjHcnvt3f3g86lMs4cZcYDllcWG/zVvkOsBMeS+B7Fp0Juvsw0ItrFmWlhxpgjH
xANapi6M3aUJZbIRYrA7ggA8GY5lq1MP/RhFU3SZXKJFk6pnCfqE3vPsEQ3+WsIb
9Muc5w7c5j2mKy2haDNzq9ORJhrLr2Mnb363nrq33EWSmWFDTRkaADdc4TROxzNG
a4/5gSCu8gI0i/Monjdx5SGlcPYJt4TMEyYAZExI+0LVM3FS81m8osEv2ujsi5Zj
Ec3vUxXlnZPIsVwGba/tlFvZXmnhiCVwOUO4kXImEPaPwXf4eIluB9kmYtFyT1f2
eyf/Zgse/a3Cc8xR0noeC2wHHtmFXkq/mcSaUfCogsG+S6ksUTIQ84e/OJjVMFFB
ziRPj4hRRl1N8yChTHjkoGeW6W6yMjS307st/SmgXU57jJQZolfCVcMQko88qJHi
dbf6UYaHK4eJyP0DvF+83G2xq0XEH9w84YR2czm9sVtNmzHfHp5w8qGWMeu+FLLw
CyegTG0Hqmhyd8EMWAOV1+a4YMfzktLBkoRBEidcVUaJ6fHWdqHHQHA8hA/WIzU3
p3Y4KBktIPiPKIVWpuBy6mmM36R5SfA+xCAxofaWv6ji5JET+vmvA34ebjENJoyG
7OeVgWxsAwwMf/k84+J1TOJYmgWp4H83UtjTFsKKahHR9Sy9r0W58AbXmDJi+ybG
teIe6sIZtlx5BodAGVfEqhsOhDIJ+TQxJVbk5mi2fGXaiIWmF0kDaT39QQ7qGZJJ
EZ+5S744ze57YKSfo4Zkd9fQ46Gff0zAGR7aJNzxLt8xjqxEaH7JPgboku6ovmVw
cpmLe5MEr4hy+HMIiXu8GLhXu333Tvdjng8Ai1S/Lyod5+vq6sHo1laKSI+/C6Po
HGnHIqLbxBGisobxQxOFATuJF8Ppa2rwOx9r486sGv+cGSKlAbkcIdQ8yKnhFDAG
Eg4hVUATLOC1vohvQc9dtPv1XAmJDxGUFSXXb23aVf0R7RqTeI8456Xsm6fvYC9G
AYBIyjvJqoyAYAJ4mg1w/5VZvYIFZFYyzaS/D524ZdN13+u9vpwHMu1vPQOvXW3X
C6beSez3wkCNfqro55mHM8gWXHx7Ob9CFAkCGokayuQMbfp2umkousydpTOQY/Rv
+BX6ymnwkQ7rNMjqG8YLMB59Od6ExHfPdP+tkEiOhIFwrTyq6jkvC2kXZiFpfH5x
1LeUze7mfhtaAKF9/FpXXbaORl4E8XHplek7YueWhwiWWWGwrk440pcYc0juheDu
neBB0ijEkW+7Aruyv6US742J+zSlFlwwc7jxm8H/jtTP3h7XHbnhrvxqICZ+j5Ca
AsWq2cApBf3OOU8zSt8KZNTC1Bmbhx3TzkFe5WLMhAU9PXQ5GkqPsxl/lF0nkJXK
mY5bRW3BpU/X3vpq6zDLrBmAjQDCH0cIwHLTcg5tQaRscYypXvOL1mv/fRVVgccq
Ny68MhZc1+tEk6CcL38KhTyU2xD0OeGEIqkyToFV9/hqEWNN/sfRD2NrcmKLxZYg
vzcEzmAKhmHrXN5r49oIHfpEdkQ2JQHcPaEuJmaFeVMayw2gnq2G/N2pK1lTCzkJ
tFRTbP1HlqUd2AB3QrNQhliN1cM0Zsy7bHtV0Di5NtcKXCJrnu1xEexKmCIenNdh
6xbxETAtWadxWbtqzEkSHnZUj4h1kIbPRFPpR3vWy/JErXfUrZzg9QwwMp599V5Q
T93sAqzsKUowVC4ejsApDfsi0Xf23HyJTgVPQhR8aW/JsYYnBpZE6W6UXveQmuOm
wvU9oUz/9vvW5VuFuvhKyQZQuFTmv1dd6l4M5aQ6eODKViJI/1hz3j3JRD0F/C21
mDtk3BuYDbsN9HAOSQcwrUOqNZbDxCXYDGr6dZs95/4Q2+Ea8oxzhemZUXRby/I0
htFG4gik9/MUp6cO7DuetrxHqX9r7ZeMcMRevg16MHX9zk3PsZ5U7Qe+i6al48ZT
P0lbFgV1hQoMIJRq/I9937LkijbxSGq8SJoyn+UAaGp4CGBdn+ZTOHApym0OC2Dq
pZmf2SPJwLSnjuEUGCJRosKWVNVSpeR83cw/lTzVzXBvquD5m1EbcJr+tAL0S1HZ
TocyTmpDlO1tlER/8x/vzclqWBGgXuuTHaQMzzDX1EhD387sysjnuRoih1Y5UbOc
GhrA2mvm/zSCXNK3sMtEPSwUjQcCfB8u8jVCACOHNhIGQjvBVQgh56Nt4iGf0JHK
VC75F+VOW8UxByJDDWMjFzgZs5QA+cGJU5IV5Rczt39j9KmnyM5koHxWmhucE5Bo
YteJjKWF5l/NfKsFy/g9oWFgxyDuHK1BWixYsFOO5It3f9KUqeTox2VgeM5D4AnM
q5PjYZTEYLaZTNcetnK/tIdJf6k9emXfjtAbYe3mJEzq9H8knLH354ZZjoQbUPMT
iemmAmNVvEslJxuKg/zDLH07iYxwnxirPmp3No3JPc6cz/Awn0HkzVrZzlN68bnP
IcBdR1R10jnbZU0BEB7Sqq9CaL83zAg/pRXyqM7NSCJH5QDzFOIXSelFFEYFxUN3
HUwm2MPy4IoElG+61rv/ygSvhemlHd7gjgroxt2sKEy56K4P6ObAg4sCzAWvcqjw
V2tWX4U0TxdwpWBFuoODm11G+ExhjouwConWpOMWXE5tyBfd7vdnVTgMZ++HWuLO
7xiAQSPYKkXxnVd/hbm5OJfQ6vcNbG6LOna2JL42xngWn71bpxfztKPqEl8fO57d
E+0GBxBOqsTpJs9RnvRhweo8Z1WbLZHWzdlxVHU5NWPFEKmszPEoTSGtO4CrSI3C
4616ZqByLO2Glxa98faushcf8IdglYYuYr1EeNG0cOB4Flnezal+2pd3TSeks3Re
Sf2RxVWJYEoSjAHdKdIVgUlTgY5p9RVFJsIbUJRCuWeSaSbk09jE1Bpxa5lyJdLK
A6DcKBX+aantwb2IWsrmxRh2VtFgrkjfQHDRgsDpIUJigVH5V0SFp+X908EXU71x
h+lpq3oP7lqGXJg1IEVWGG6s95UxzX/dzImRDqYg6wUSoZh3yIM8ui4uHPeSu0aw
Sh1HZwybzumy/IVa0wSWi1k/WnSoWdjfxPnTUFUrTrZ/ij95FCeZTnwduXgioaEI
pIoLxMCVYv3SMwg75Dmxqb6020T5QqFqRfw0zHwMsCiIZR50AHtJZUmB/8sW/fS9
RwNEIUNHRBfw+V1xfAGj4eLbp+Lncnqdg562HSnCp4D05l/O6csQGiJHf1un8SJC
BxoAf7cTrrX0OksgJ5alCKQTxjvMgxhSO04CaFhck1Q6VK6ZXQFJ18gpd0TNPyr6
zVm7P/GzaVwKDCP2VykMR5LSNpBfPdMT3Eh5TQNEn8Ocu0NM6M8JQHoMz/dMA1aO
1jj+2bWs97QnSCGfLKmNcaU3yUcqHux//HdXCILlErODqHV/a033MDv445Mpre5F
lzIWFEAm1AkF1Miy7KkKStqyXTxcogNzzf/fY1pIdGrOFNfLAMghHHxJHkZmfAWy
nilAU2JG2y56Rfkt1I0St/phPfAtVLT8Qxi+EvDlki3ExjswndFX9MhHy0J0B5qo
6JeXROExp8e21CnCNh6Ed3+R0lFNZ96xDF6+883rOKJKo89+do11dx5I8RqPfCcE
LbahHfFqJbgx8gfWljWLELpTf9dzAJPUDWZM7i47YzOlP+khiAbDuEuFbWkGSbpW
8A48nXqzsSIn8Ft7DjB/gAnxfogGGD+ekuuvAdagcUDD9M0jmERdPogUHDV2stAF
umdH9PEPfwOkDq+McD/6mYbXBLEobrfvIdkiM20ZyptzwgEmcjoHI+zpzDrvzeP0
eadJ71d1fP4ooxx1tS+UTbqBv2ETrTIthDgSvigaXDoiZA5EqSyutDHmlcGZzgdf
8phMCCh335I7r6OPuuphW8BtXbBIiUzowz4aUEz5ddieKVYdtOVTm2GITQBasdiz
ftTDuB/UlhXRxfGNZXuk2DPrsppcvQEHw2yiopvME7ULpWeAO27+XEuFyhtsfX2h
hNqqjWeqOneZezkhuHIIsveFOWUsnGeHnM4gBuRX7MY32F/I3XLpWd/8Lam+HlWx
60/jqY+0vzbw3OaS+1JKWirsu4A5awUuQy5w29ZhDjPe9EAGZwRsLg4lFrAgcXgR
FUhOsMfXF1s7wKSkgCNnShcFjpW0uXPYnZs45mS7rx+8zw++ZNbZEq9/la6tkoQN
RUb1ISP29EVSffyUU9SwabgZXZJO3bAW/PgvU+lWoOp9f3IxiobmTaSZng8mtNik
FS9GViMRMGMGMVLZBvxxe8eTbjaovtoHO7ZZ3D8qCWGYDqaAVWUS9W8bJ9ltKcmm
uz15mXu6H8hEHkeV1ouhqC6cYBQTBr30FXMNP/uINF/FSaKPVQPvhPqMj+hopqHq
kOY54bueDfpEy0dcaaK9QQOaG4mVmD3/kTvzuJy/nmndwWxihmwX5JjRuZ4k5fCP
7GH7XFFvyF2g4v8jDViwJb+olICRekWPQ16EPyd2pbsZ039sZxsSL4t4Jm4EY97B
T5F9lazSDiO4HfQCOjSSsn1oiyBlOL0SyrDAK++7gqgBkWUrbEnoFp8ZTKity1a7
eY1K6Bsq8xQ3el5uEMFJb7bK93azSFIWSoHI18vfPE6tA6XG8LPG0x3N26dDurpM
kfzmP8Xrauc6FSEHtMVVWsj0w4B3faladiok7lrJhw7ZcTudkkcoJ0OxuvL2pRjC
cfEqUOvGvLA9FNw7kifpF09765tPE/arGor54fm1b0CvvHOzjWxBHLJoIL0rWOVE
F5qCTmrJnTDAlEDm+qEoSeprvZ6AzJFLJ/9oFX+NKHx8HUBMmgWb4W+Dsl6hZe2b
jcVZDYoLlCcDLzCEyHV5yHmEGyBEMHTj0WDJhebdkIicjRpWZ+ofkIlPvDnjqoeC
9ypq+z4RZxb258pgbnDZ/u0UaPkl29TF2LrERaAkqKnA5jmtaFepeupPZ4QsTCw2
P9KFE2lBi3SdvlnqKh+5VcsGWqZxWKjUvGY3q0Njndq/TfcxMHcbSwmX2d7UAX8X
lObVKVmkjHVK7nYo+e7LWyWlIwRiKm8d2sfS/UOqrskPTjK5VByA4G+i5ZSuPSia
+/qB+gqr52gxIHctW7SFP5kxAgHCHTGTayzG0PAGxGj1/EPodATMK9Vh07WKhu4L
by12wDuWcNgVVQMmYRLg6fUs0rs2XefEprOoYiAPbks9TOVxWrpV6yJcF0xZBQ+x
lhSAvY7BeTnpCOYpoTG1qyUABFoHNnw3PsjRkXkThSQ/XsxGZlFxh9Rf2A8pLp4s
eRxY34Z6GVBIixb5tqcB/h0420GSJRQduVTOP51lxBNCaoPYYWjDsY1UEj61Cr33
jhL+oPKahXcZzTXO7GNo2jA5x8DUplsBKPj0y00AOjVNYeCZJMhKAJQ5s/G+UeLk
yreKJC8vt/yLOyTvYYQVzRl7DAPt2oteqQo5G63eotHLLmSq78/DAA+eHJhAr8o6
IWzuPr80TtahWt/iE740/YhgQHGzB8m+F1s7CtAeMMVkx4q5xIvmq5iiR7lCyqrs
j9LhO6DGIRzP/vjTtLF3Rc1Vf99NOXAHqQPke/XRfM4qo5m9alFG4FzN1aGdIj3L
llgF7+AashgjIxBFsE0wYL/uRtQczQ5WqcJrZPoNsedoz8qxkttrHC/qTk8UZ9W6
cS4KezqMEtatH/YchaHZfNWmCOfSeOKsl73cuGkgWcotfc9mghJRL/wt5PFF76XC
rOzY5BkagLc02uHmJD3fBGnUrvaHX0k9JXN0RSwYE/cZplxQ7j2tAV3fx7VU1qck
m6uRtSOEP12sqSkEeQ8EyQSKHipzMX/p9B2jxH2NyIeJxsaZ2g7RpKkQE6C9Mqhr
uxp1Tg16+itV1HPPsamuvYLSxPn+YmjfhX/du7JYkSzxHjO10K/+gJfLXbubmsO3
cRExFBe+Wb+i+1VUk/0c8a3okRZiZhZTuRS5WvZuIw80R7JbeIoUN3GtCz6xpIyU
kD3RIPkgDES8ozVQw39Q1uTrxUv7X3YxnpwnANIQZhT7FZk2rwb3c63FtL3KOpZM
2p306OcovjHavJ60yVYIH3lVfuJZbQ1pd04pNE1Kiuz6/4CoilZHgvNQFKMc+lBQ
CnlMrQIIi0LKksVDxaT6xO4AVm/5ArsR75COmC1zuf2J610J82OR/hY4YRoV70zv
KklxoxcYyMee3CaKjTPl9f43jQIuM5BqIIrHqyMob00mMi1x1ydjdYiUCUmxXLaW
sap124I5Y6CY9JD+297JQZiZYPX/95Ren4ZAT6TZmdj/iVG7bJtA9PTfdid3GTEt
DScp4Mm7zTxLr3E1QCMyphojSn7NGMgM9hAiz0gRw/m1UzOnhq3EleUTbMGiRqgc
ZOsJReS/2WyTFWsqoMNoz8mF0gMvBJQJGLvNVxnxbrczmPFF7TmmtbAS3aXW6xCg
TmaYupV6WikxTXmOOQtMe6FiptNzeA1OZMvC+71WxyXwblwAtZqnr95i0++tCo4D
RefYAlcz/ZIUcsvVCOgFqXTKGYBd0lox4pOMm3QRK1YFnCsXGlNLDdUiNaTap0tc
+EpdOLL+/AxMAdCOIglo7qDnVrK7zzChgWL/hngBIioDhuyH4AMjWQtaYLFjX454
DyBJYIpnxxu7SAyNpZoi+m8iO5OFCx6kFH8hj3YkRoi5D+F+zZ14TLjJL/JePgLv
zEIxNyxK360MksSb9AmXVP9aHZVjqFzu/pTKO1c3v9/x5D4wGpKOPiIlqP0Jaou9
igF2yedNdPvEx/NjlPW2yo6LUY+UFgYouVCH24y62IMqumXfIMegsAjgaHbhrSmd
uME4FzQSK4muKxu+6iksVdtVIKpWwGlhLjsaQ9NVOY0CJHasL1now4FMzdXcT/W6
E18sNg5R/TdDp0WoIm6boyU01YUsUStQttYDVkQbFjb3y+caXJSFY6Af3pn72FvO
xBPIGDVXShJV9VuVMYhbylJRnwCXlITfGUX+MlWGxeIoGzAdVRlos7O1Cfx4lK1I
60r0sNEcChhWwpjvmzO8Ox1M5aYtvBysLyCeF5OhUb22t0sOIIqM2q1vpB8iXQu0
hJIxG1ibnKCgN9KbpKi9u4+aoYKprWuXW3dBVvMCuTVbcGgec3WIrDpJRMlqYyor
Im5ZKJ8ncOvjLyj6mz3RxJ+kOj0xVneHFeczbTEiufCtdQ7Nw5n02jj+KwIwzDhO
Fk9eHcr+ajpz0S4TAp3iPl/Gx5Zxy590++iWtcyNN6oZKzhBfqUvfOu5YZAUVh5v
2o5xMkpi8F4TXCA7xzEXRlY86K8epxbBWf2cGYLLJQWzSYvNdqkRJqGNx+DHCjlr
s1q8WedAM0NZ9h9eXRGuVU0fvJzz+GCaYCu0SjjaHP3RInibHzeGckvLrPrFUfID
JAWwHH+Ghun2SRDBjujpFSmumSrodiLx1JIH4EIZBKg9SALXdODv89nT/pdqpX59
pwvtDBtwlwCigsaFFz0jh7g02b7TOZvWZRgK2SjpY1lOXPInvKSor3TE2X2vsr1C
POHqUaAkj0wD5t5PLA0MxULsIKKV9kuEeSmi/WVmiE35sNeLVC1RXfp0VFu8yUZm
SU7EQWysfqOtQ4QgkHuYQgkWIhu+OyytmN0oA8YFAymAF+3blH+yLhorxZOYTjrc
VKQWcVbhX3q5y5vIXa8oqbQ4iN50Jbe3NIwGbN2PG2iyWC0VvsuzVKBJYsji1t2P
VrNYufSFTJKBv3kC+tQg9hPxJ8gFTqI/l+HdPL8Q6PyRwyXjzcq4ntcL1CaUB5e+
jKrW72rl3O9IgylvpT5CYlK62fR+xubfnJOvNd+7lRNG3tCgX2l+IVzBX1HOQISv
dQqwiLeWQeo49sUS/aTspH5wttcQC4umEszn4dF7E9GG2I7glrtLjQrMs3CArv0A
6gje9Htrqo05jG1YcvKrQ8vmiwDEXTFQmSvbOESqMJ5lwhKHV1QJO26uCS3f7chE
jsYkaxbx4V4IP4gZKzuf6JU5+uOG7DVq/YKDfVHRsJWqGu6phbu2lC/7Nn9lyPkU
i1tXS8GVqRhtnGRPTODdGqsT0/ehKWIzJR4UBlkQX5tbgrIyyxc+HT+FHeUgU/PL
uD62z67a0VxwIH7q+MjqUpLFSO4c6AVFd3cLuQB0B+IExrLrYpiXkan1WfDCah2B
iK5GH1kqiekrzj0/qM6QGC57V8EIR94OgUAQXJiwt/ZSjeLnPOUSjlUDUtyxfeSW
dDQBgoZ8nhh46XnBfglyiTlJtcoHEFgEfnfNNkyInPm9m7L9vytQjHSAY2S3y7O0
9ophdjUiNNnJZDtjw6IKlXaxsXGyj8lWKZac1z0LeQ3RsG4cCBGCAkvKNr0bn5RC
80e4rxcFpfE7IJ/EF+Lfj/KQUj6uoMRQVKrm2sYutRowiY1LQoxXsC5Oumz7Um8R
95t191OuIOVck3S6GzBfz/4tqi9Z5kRbJ4J44HC08tSHaJxI2IXnyx/bA9q65PC7
pcS8WyvLN9+NiR3I+ArkSQlunuZLOP6HVWURdPM3luEYiGQ4r9y7CzrwQQTwuB4y
tpWKSgxbElCj61E/O99DHcrnwN4tIUd3DSKJ6dBd1YUfJXv9jQZlpEwxmblv8Ivv
rqqtbq87Pp0XUBYI2/G0pnWcvV7jUjE+UtzCW7kFaHna5AE5MgyUyM3e9qKR/8mb
x6oct3pOfchX7imBZKkHG8L8GjXHxTpj/vf4xupmxAdavArZ7l7tUrjaz26z9oC8
wrcosoly03QyPwXWT7mQbnREzKhPbC/zI1UZ3+Bttm8nA7lBuy53FTa+0IAeQSPu
FFGJM5HQyrlluXz16ncSQS2298KFIJHk6zRNGQdYlcLKw+kDHpQ8a/WolSWUI6UF
jNVsU3SCFG1GYwd+O53lWs7VsiJLBiB1F9Z9ajO7NqqDHyWG/7sEcFRNbz9R8xwK
6gacxKmlNzEOCesVfJdgAvCGloCpPHvPt7SeCo7WUZ40Br/FeHsWTpWWuyhDrAGi
Z1OBOq1+8rG/tJpWeN08l5dpi3kkTwuBhVeIm+1IMrF1w4OpxfZrrTDV7kOLJfMS
ymn768ow02v/4C5tH0APbzyZShUzPc3YCkvNtBK87R0Xw+0TiwICnx6qFFbS7mlK
AsDAWXAKD1M7Y88DDzYOUx1asc8zbY39sKYy4F6Et7eVIjiuynYnmiqvBfQB0s7L
m5degbIUpbJXc1014bfuMEbp1MUKs1CpsHchltzVgFTTTXyTX29sNsBsbV5PgRlF
rOaRGov/9RRFr6zt7T8217xVwkisQn8qZGsnnPP7UXdJz/HZqg9PaIfG/2OqpTEx
/UimTiC+s7BexiNMqV4iubLK36TRFAP8aV55OUFhf70BWCARyiRUsk4+0R83Fui9
S91l0EoDg7Jnejzqma7xcDaLXuiQ2aMiTwoRCbpL3A7MQnbCr9H0jkCZBP/xu9lr
juN46fIwXfaTTj01sSxr8Nkb1CbQYHg8k8X9zt+KBL0mk4HvhMgYC7qrytdockBo
C/dkAcFjtFtQ0U4l1SPJkDrIcf01APNDQnaP91ny4rXR+JHu41nY7JGs+zelgcz9
UCuUI3gALsAlt0H2yzVgxVn9JhBkCB2xRbi+gqd06H9+lFfnOONSztYwzZDk3ngc
izfayW/5WontHnqXWERM5QHX+NAVbDHQfg+9yX+9Nipxhn4W4GibpdiUIaNoba16
gJgBpXXnFD6CYKVsOIyJBGX92nZHvS5+I0S1pspx9R0LuGx9GbmbbBJ8ZP2CRDa+
Uz5RIeWIwre9VM9UosF5ih5DPQ9qIpS5/pXKG3bJMKh3WeT+LK03k38nVwH9vK8n
nShswD5xaadXlPJPBKUd28Byb51r/1V68LLv+e+ePCCbbaTwfMsS2+emui8vZqBB
PfIf2T4P2oGlhQ/AlDZJEVANp5p2V9TyVG41YkrANGOmYHRqtsDUy9Y4EAYDgOAc
zeHza74pZ5Gr5vpSWbGVsQvXClaUeZEV4CLQ3nmQE7cKYI55qcjiyPERmzLqd8Qa
BREmhKILHUGOatVE3PxAxBohyRdObj+T2AC0xvb5dZl1R6/PaXXw9oK9YE4wM/NP
cu0iqt7kxq7Q7iILe1iG7UXc3qTT9DnICUUFb73JQGC7RptGDUagEmoFcN1bQSDe
OZ5uhCNPtq9p1OpgRtcFPVmlTJtbPaBdmtB32db2OSDAlo8wBV+x7vuNzozEXFNv
0Y5LU4BsNkuKySCBElSmVNxN8QSxbtmDQKVkPcGZ8C7EzBNFwd2nBpCBCanngG9b
PEbj7lSpb55NLqhL4Pu0Lta7OEzP5NF960/j4D7uN2Ad0K8q57XtxctagiwxcHHv
z9ALicMcUdNdMkA3YpgJPAbc0hCJjGpiKVAWmuaYNYUti8ZXyAgjP+myZqVzk/g+
PU4OZjgYyO+AFBSU5LGC5XHbp/By8kpBjv05SQKDFvCKfXrC4tew2TT+sJKkIVHC
uD8aCyKfBNJ7XYB9Rux1cqThcLI34qEnnrAK1ycUdHNWiU1DzCGO0WdiRxtLkIpQ
aiN9JRs39yev+p5Zgjcgg7zlD9Kv4MTnWsV15UPbNnN5BwwIkbPejE9Y82C8hQ4w
u/1EiFcPDV2bVOxW2znXNn85IFvHvfm7SIhNbgJ8rUw35v8P8Z+u8Yy8mUQzrLtF
EJ5Xh0VRGlDT3TM97UQXUug++6/clB1pfgM35mvNNkJ6Jjk7FfalX5Dq8VwAVugI
TCTJsdqpk8XmFnad4XjLS4vPkSgGV/unXglSoujPan8rj3gFTangmi5Bur393iEq
Es2nAANuFFfZNICXXAAq05nVixdZ0zlXPqfYsish34/KgupkSgUYw9FAEf44VaVu
PPAnTVJeSCoyWeHA98XS99GChun4pZL3bj1CU3vnKgz2il3Di9xp2DIrB9xCuAeJ
blq0oD33jwOf4jvMOXKVhfhEFNAX36bRHT837udRo2KgSEX9HOmpK0NzGj9qj+Zi
kUj7i/JIZOOf2NTs8NSRW5SG4pE2NmDfQ+4gLIQqKeh2FVN38ungNGpWMlxa1bVC
Dpzo77pkL3VLie1XPbStx96ZCRVWSZNTXkNOHKaw/fgEh0Xm4sjpYVDAfLIXO0Cr
XEPDyoq9UQDuUXT1deQE5prJ6MVlFhlPA/60fUQFtU9Vv8USb6vN1wC1fpDvy76w
XAbzYUzq+Nk32uHP7lz+nJCnEOEfCn5iSluyVTAa7z/ESCCwS2fnhB+l4iSn9ISe
7Qhs0FtbAQ6Q9TB/LiBQB6CBCVVPjvtaiJ8YDXfKEf5reAoAUHFl2Ygegqa3vpVV
6w7+IzJdouSANJ5QSZ91/r/6sr3faynzCBOvXljLZK5U7KfEzuFm7HnmfpyNjcm7
FNCrgcOaPm7UuB6a0rb3lnO3a2fLiGaDeNL3RcWJsT/YTCyBcgafqPRHlQk6hBm2
IzZ262+4+WMWs0Rq9ZSBNQ0g5HI3oH9Cj+Rnn5AOb5+rwhhZUZ6MpvWnopLrhB8I
KbU8a2UFZo8NWiLC9ihZKfKUinfzIMQ1HfkwcD9uZGbc4pIEMj7zmVHybz7JmANr
f3aEmm7I3okdFCwHXpvUymj3S18G3+zefB6pEBXl9fL8BEYD+myvaAZRgv+O0n73
mDcETwXBK2m+CfxsMxHJOFjMy9GGiHMMtLlCTClHHhqi/bizKptpY2Wktx8kgMtW
lRlzXjg+aTdHK52zYmj7nHbJQTg1w2uaT2+FpBJnVmv8oE8Vo5ogxfvcjIvOj3AT
FGoQ+Pnqe2Zus8vZImRqQwRQ4oJz75M5i6t6n14tKiUi21n5tWGX1qYPHpEWAmlr
7H1m4M3HnGE+1ow1gmdjlPxLZRJU5Bfkdo7Pt6Q11hzc0WfbGyrdrXi03cMuMydg
1XwtioDKtyAJf6k/fZlyVgI4v9qd9otnQWK4b0k0R2Gmk8x7ZK9OTk5vvkjHLmf6
ixvcnmPxD7uJEZaix4cg0MmRNOoFeZwYcIP63vCXyTt6hWEoWP0qRf4r5ibtXDqc
+zhocDfs9iwYm5OvNpm7VVhccKbgMN9WXAP3choEsC3H2nYPfX6fvmkTAfyvWFyi
lUxqyVN2AYV3dMp4PuOvgMfGJRuIJRkSma2YBgGtNxNExegQHmg9HywI7pzcKdGp
7Rdy1StRcczCt95kcqTDaa8pjtm71Nwgir9Qo3EwbPsR6NCCF4PNWec62Vnh37oL
VlIa/PBFiWHdu2uazHtPwz/WJwrA9o6ZMwsMfuuxNnDOipkVDN63edQ0hcg9p1TC
APznYcBp0JzhGc5xCjLVnI3AVjp+NsZAsdyXN9q77EE1uKnmM/V+oHW1m967X8pT
CviEAXqVCBLhrdkGX5OVWVDr1dR7NPgbrJIYOLkEHFCLTU72X8VRnV4EFGGZFe7v
/q+cTd4L0viMhFfwDdDd5dFJkjEEKsHc1g7lYQBQY8FxtBqEMJQYWASfhwi05rPM
9DYSpycyTQPjgdBS0SLn6Muw80Z3fZApQD9H5GB8oC7RfjYU8bwOpc8kyDm1TMsZ
gx7Vq91Bks+fcEl9sryUg872WU1n6667RLezwTVqqZvGG0dbOcgsAJ1wiq2/N11a
ti2zTrC31q9ORgb6mRcbq/wLYyVyKFv4twaqdnBLtnuFObnhB6+ofNpMKvvyqSyA
sgmdqJjtwmOer/43CD9fjdwzsMcsW+Z3T/5SQyji8Ei1gQZprGQXgENW66wV1EEX
/UY8FTu8XA1GzNVeGLwJaUNOJNSl3csGra9J83J+1ltBAGBOGsplhZYIukatHbGs
/QvSqYIAAdKuU/wMk3qGs9rMDkPP/1H6qIGWkevkY00WPPezt2fSOzp2nOMFHtoK
3kkdXmEHvuikYXbi+e0Xypt9ENHEj7zX8/kkqZvNaJFpzzudBAKRxNJ4Z7IrPJnX
KB0mme0bvy/8b8GCK/HF//ig2cdXL4npuqzLogkH0tfe1yNIoXRHFiZ+XYAEeI05
6Ka/RRYIkKOozi9xgd+5GretNa3OPXTQNUQKmzebW0u3T+Foa7+wP79wKlovvW4a
vedtUS/V+Z47h2K1ByY3kHW9SlmRaxa7NihHcC8HWYj29X0Qx0dqkzFg3DKJgBsy
J9XpcT+/7uxCjCNo4Hp6OZ5pI8CBpD3e1XN224zRp3LIlqhmk7asx5lZnxUbjAjz
AT3EZJ2KwN8iH6A8DUzOMyRhPc5nIQm4I0SLiRAZNGT+i9uxVxWwbKDrdDzfzXiY
DWeZonqmjgN0MxdK/dxmCjJGeuQr1548I5Qtc4igirUH9Dv7fJL+ftSH/n2aMVm/
ndM8F1K56hUpllNBojHy9PqlKrVaNEjpF+xn3PoffsbOHxuALqAjhOJDxh0tZEts
60/Xw8JRlmdeK3iSu2koKpdNKejH7HLDIcE8hP57+JQo7DyScWMhM5DE6sYviCS5
0+Z4c8RLq1VnlaRQjWA42W9KN8z/tDJ7odrBzpHBTFl5vkw1zHxM0oH2saWUtCmJ
zxnAoxYrImNKVTbpvTU5le6t4/Rl5wbB5sNQE2m2PWSttsmjnluiklYaxpd7JXQM
brMBuoSKYGrtpKX6rebZw2rKKpCDXJgQ1HK505Piybm68DHSuOMqm6nSjTLcPQV1
WK8CF90o6uX1p464DlUyQzCTaMP7htGjDhqzLZCvKMVqBmEgvsqvweKc+xHMfNwm
4YwOtKJMnQDf0Zd+1ejwyv3D0igqjf4z5ldWoeuXzKRb71UxvVGSwduHZhHOdrUW
xJlb3DeBzsHoqbIw778agYPRr1XLU9krCvJrzYsdbYjLOcQYNtgYEo0SNUvUIfwq
S8V3eLKK4BfbPrhEYET19GDgBkFc37LXjaY2Q0tA29/mpLgwSfgZaQS6g4RnTojc
PxEHptyDNtJTz5sjIPUUcs8qWWiBX1cjjh38dSAZlkClDMeJnpP2nbhMhEkuP6tT
+t4AvsKOPFYd/p+WQHICPczMW17w7Pm2FNsyv1N0F0BN0uO8BHZEM62CpqOrWXMQ
/bUNCtt7wJCIMOF0clasg5lmrtsFOrpefb1IIXLuVY8jllJxo+7udE9Ub6Cyo0h9
CUR1C8woasb9zo1WbRluyeIugdjJZuukDHWX41+SCeoVCoxCd93QmGzcWm4eoN87
VAonSyCpUyKhRkZ7pug2K0edF00EpeQ9TaOeUMdGIKiqvO+MT+g8SfdRurX3sGM9
pYq3Lc9FMLlFgxeMiriS8kgdSZJ+3U7/7gcrBG4kURp8W5YSoskei1ofs/8EFRsl
DlTqUvG6U5fm7y9XhRs46Qj802gKck4NDDPWennICf0j4Iax1YFrxA6A4cRspwkU
sEPwc5HaJHA6WWUUciyIwSfeAXzXSNkYpg1fo2Xo+0tWHfaUNlNkmMY203iifBpx
Ufqk32/fyQfWYBAnYJVWqryvynOvO1vbqhfSLw1q+uTsGmKLQbWsjafG3NdiBjyO
KavbfLzPz/iwWfT4N2dvPXkpR/SO/uJyKcQ7E9B4nBzq44Xu6EdjoSL7picbKkkV
Sw0fadISWEq5MAJPmbblD7La1DcBoBEPUKbZpumY5eOPNag+/57v3XCZjM+D7M8e
pM29xrgaT265O/VtEzHEzWcDr4LbCaKcLvYiJ1mad8n/f3vXyjdN99P3xnMQaDEw
uWKON2xmF7S0V3RDL7ImxAptfvOe2WrrIgtH+WQLfC75fh5yh6A1b9Y12mwdnhJo
lorQqUbFkxKRZCY11y+oNeaVESTcjtE3Fuk0riep5hFQmbh3me4JOp9nHLTmHJQE
dDv/9nlGN+e583Z4jw2O2i4SfGGXVKEJpwC7d6iOBPmTXnSo/ZMNVIdqoNX6vlYq
r9fQSbH5y7GW3eo1oFhNRDO5dpjFKo0cgrPuM7PaNQIS5zkiqyX5tNi1VxO0l92N
BubZIMOF1R3ZE3tg6kDJCp3/tT95ZXVdx8EykEpdbofTbYjgt8/LfFo+2uoxw4ve
4243WmT8U/EUB9f88gKJe7Ugr6ofRG36VMUGsBCXMrvBGPzeTDL2iuAguMFOg3qt
+tf0VqwPm5WtRaPy10/w2BNf9lNZzEVKH+Q7oNJt55DVmsst/ucffkCxYoNbuiu0
JFYKQT4dS+l7/Nlb4Ujrw2zmeuCYHAfAg68bOawHZ1JuS1wwAACrim2O+9dzkGMb
21E+YNNLoujC+XPu0gGxDR0b9v0Foj57VgtkuFcZ31PJMazwQKmPFryRAdV3SFon
KqvXnAXKNTirs8Y9tll8o//ZLdyHh++O4LJUgpesFTtxjILzZYxRSp2zJrH7qpip
+5znTgOXVC29wkeX854JHmyJnv40SHWsgzeCsQyTiXtLIVOBIaHgXoRPKKiM/OlE
pWzyeeQHGxXPLeSARSH6koZJHZQNLsTsEubQRut3cbJuVyj5xHEZvCVJHN9Fo5Bj
6zF9VV6vW9kBIGas2ZQqx9SY+A6mpuWAtnOqliHfEhaOFr86haD7vdJhTnS4LsX6
sWdpBnInD7LnyDXAEJbq+XRCt3i2KINce6tHCe02KqyQ7qE3mA2maATwTv5Ajbh3
WCcAWl5HhJwmSf7wt+5a3+GwJi85uzpb6uS/uZW2ScL3qjK4lRBi911qvACB12Yu
6uQuBIxG+5Hnj2Bu7rKyJlUcx+FKXWB8rC7GKIQmadqNvq04EqnrbToAVZ1o9CcD
VyVSDPnHgtmb1+lJ/z4H5EFXDyU+BoIwVPUJt7uaVSm4EtpZSDuIsQTg9K1pKkV2
vMaPN5dT5lPEXcHA40537lHs1WyuzdmkROZqbuVwZdCbyXXj3cf6WS89xIMut1zq
mBCn4IeOwJWzFARt1/WYTCkR1SNp40BDMKGUUFNB0uCB2eghl3sp8FEIi9sWuSMO
KElPAM2RCTDKaLtD0YV8Vj0B3QwCT65uSBvg3xFRmyIofeKBgrUHFLv2yJL8u1uh
/SR9BOUEY2026r+hRu+t44l+eaUgoxhNypHhqMbL0/lLW3VRlU6ORKR69COSS4Cm
GFPJKJBsx5eWoSmAfV6HvgLIQ6pI5TSkK1aYRnjY9IVp8Y6lnj0SWuCID+WiPw37
rtcfoUrxbOSKIRjCwgFaFv3hKAgkB5Wy9mDeSDlTVJnsRUFrhD76qZFW74tu1Lsu
HfIsBZMPCybO7atP8EcdkuUvTe4ESh+kPyEClke2aNQz28aZWKg3zKD8mC3duSfO
5JHX4py8sD68W5heKPo19yWpBiCNHr21Ja3jzAjdT+JN9sQDF28aNilwLX4k0pHS
6pvo64uwXnc1MAMY0bQWhtl2tKmTqirv5FtdscVPXI/IsAf361IVHOFchPFqtB7r
zzqri7UOACROHxRD7Ujhb90EsIQrNtXWipbSXuLe5E0u2637ITu4A8zjNzBl18kX
GDwOjwjh18Ipst8VAe+FjBetXABN7sDr0M8cxp9f9Zf/Ivfigqf80lzo+5BL0uf5
p/+dlHp7FfaeG8Xt/wJeSgZTCkIpLC7SIwH28uW1Opja93MzHJdZZGVGWgieYn4x
1EClyMVH7eO0z7mmJu+UJqMmE0nI0JLCMDlRTKp9elFxftZlA/X8yupx9ijul8/8
seagLGeEKzNBJU8RTCY5KyLTr5KvL1uirrVqIMGdePQJIImr/jZjbNVdpx1eD3pk
hvajsLILbKIctEHJvWtyn7kD4wh0pNWsgDzqaoxqMlgxadJA/4eA+1GjW12GY5lZ
ESrlMdaFRq4pbS4P3vbhfaR9tx8HgiyFYrmWMYLrEW26bFx/7Hj4fLTNdzTAYx3e
dktlA2DUjyNn+/h1FR9cT3kgmYgHQXx+MzHPWvrqee/KUhkkf4C/FlFlzhL5k5PN
J9xThISJYj5ixjh7XMW8g+6HIvbGpHU6fatLKl2+aCAhXev2/K/vbmO/qGBQ3y2e
jfZNNoT0mIH6z0wUUFLFsaWRYnhY4h6cCyeOUIgNQ+bLb0tbkQMR04PALWJceXdV
qfD5FjX7fz2V3ZdiIJO0OJqtcS7xkHUhOP62PDBvDieZKG6kUaJP5CATE7VFdDVF
KtFut5wBOBZIGGQji4gK4VerulHBrNMPZqlhfF0Rsmq3YpcQ3Xiuo7YNvjyQsoet
Ps5/HUmyc0T1FGcFuMmGOllB/h73LoKzDAgNaYejMnpJwJJmy3CJwf1wlc0RlNBF
wV0OucZnYMcmCLE0krslKFZrBMIeTdL5C+QJm3YGGEJgJC3GaEH8vJF2tJqu2bkW
StkduZqsspEabrasWvRSePRiCrCjsahlYh9zlNRxgbDibIMZ0jsrCcwR9a24KzpF
Vb+ilyP6TbFFsOkrVgRHPHWNG1yy5lsxcjJqanP6JdXy2XkdS19ap7CDK8akDNLi
8lEVYyEgzAjJg9nLKR+nFjPFaiJq0t3RIXwT/OqY2vhj8pDuXiLXNLeq6vd//vg/
uE/Nuy95ql0Bluh9b+/isg9aM2auFesZ/fOPygZZhRgfJ6vFb0wiE/0qRxGNg772
rBiSKAxqkFAw1S5ugSlHlzAFwbwBAOgvzyZ11VLE8DuN3pRXzsNLN/5FwAS0+zyi
R+2G82BfJJEFe9CSAusAcIO3pQw1WNSsBix8B0n+OiOS2Zdsuq6R9onvWCIomvzT
nfoCD0k6JaRyyA/VUZIt+O4qC+51EIr13fO31ajp9AZ5y5Ma4WcuQJ7h/sp0mD05
bFPIdLomFiyubK0yRP61g2a+3vPrCNAxYtXYaKNm69VVT+sWbnBLY0cCPhfaUsI/
quJfQ9poEDC3TzWWR0fT+8S2upHRF1Cz62DBKS4qlMjFcC1xqa+7RfJW43yXE1ab
9m+umOy31tRjJDM3DBArycWWoJd/MxT4oHI+yoj+/8jU9apO/vVGPE4t87SHrnlw
rNfEiHh6i1Bjkr3OEXts7H9TSk86V/7E5PtANOWpbQjVFXrjI9b+ebBShu3Bx92k
NlAnWM6sZswnxqAxLBuBEsKtaACeGT3IAhH0QX9wVsT+5XlATL5M6PeDMz6MhsYk
r4RZ8ZeMvRNIkU3lwrI9TmzncDrT1BWVDI8YBiBBB9RfRO7U/v+eTBtMm2KrjPsq
NzMKozna8qKAvnLYlG5n/Miys4duXpUFOhg0qXPg6oRr/sjvKJVFnr3rBWMWtxcB
q/vRvAwmuk2BenP7ytETP0Co5/ii3e9Ut2Skks+AWZ8gsW3fpGpB61nbOjJ4oHiV
NUAM0sFmFYAxUmEHclxHBroiUpIIu/S0FFcMl8D3IcvnCTyH0EYbsP7ZNyCBHvn9
6ycSAioBFVt8JjLVVDATkQb70JE6iclAO4/8AIFXJ0ygIOSTw1w0z3wLtV8MSmtS
Z3qho9H5MGIra/G8Hb0aT73hmI3NgV+4gj0AzcAw6KT8ggqy4JzP6+EWKcOSrnUQ
2UiCMjcvuZ+fYPtIvQQBJNMUEooC9Ozl6E4Bc//AO/UlC2xkvN6ZLiNTp1e1+mJE
Q9SuyRcJuVyhR8Y2f6w+i19WHznwK0q+hAhIWlW9BNy6asCShrNneainAKbUxfS2
UoJiQR1PBDBlzvNPmJImjkVpH1Dn3xYP6GuUrJ1nTp9FSlwJzSsIGjbZwcj8Aiyt
Qin0DGvC07rAEcCNwVMqLXxi0KTTiy3iZkCDZWw3uXaxZGUOKTYrX8C/jFXM9RYq
IvPik+7k3nE4VZjcOZOvYC5amV3uiHAjrW6dzJcWdjKIfcDw94s8DhqMyC0J1sIB
BoAH4k5pvITaKMjdM2UCntmaenhG2PWa8sCf/idzmFiTSaIVxZUEYJucqfNuRJj3
1v60qV5rzDqG0Y423au2++kzh8hHAAZtstC9tAHWfGc7yTYnvV0AjeYi21Dl7RhB
f2OW1gA9yElPkO88hICosQu6MVbKh6Bqntd8LWJQNekkoWzluDC4NICTNvJmo3OM
PzasKCfY/4JhjOpES0sVfGhXH3UADXGPhOg6u+SzBB6aGP3hzOucAQ8FE+Usk0aT
j2zD7pFp9fleNSOg68PlmO2VpsLarTEzbJ4RW+FvVkii/gz4xwB3QqivsemZKZuo
YPJxIwjzjbPGcJ2oKsYtSfDwynUFALhS5H1UKrXoKI22oIELSGsO2eGTX+VlkTK8
oNNydnAz+MRUMp9JuhM+hwUH9yG/q/pF3RCRLG5l3MwLtNCKTXZmX8CJAn13sWcN
eQL+ol4CI7v85xsRU0qenLC6OnV62XSDT0iDeLWuuCiJNaRCNKAr/bGgoYmgxSdC
wQQlPvTzOFslSvupBcMWcNhaDHjPpFTGtwLrq/+BvIUjb5OwuYPKYDcvRRm4P1me
5xpheu+Z4CwDVaV6v98CsAjljs5O9makHbShUxW1JxZiqzcOxe0q7D6rTcLZPHtV
Ccqnt3rQe+bpgC2OQs504Bm6iiadWKlGv4dw6+zRDGFGqQPL/xnBm20MH3OsfPHA
t0oZEC7X7C+mw+oXUrjBoqtsyY2fvJ3rIEK2/6dFbJhBTh5O05kU1HR4CtONvpxJ
YhITWbknQURDwZpysBIKxkcgKh21p2mjXCya0ad37hq6VczRGL2cxYrK/h1op4Hr
y0fbXUXh/iZsq4ZRU3IGZiUJf8gdrwq7Qz3cneypBdNmerZEBGEB4d/pvDz/HLHJ
bZ2uUOXHcatcRc2p0SX7RF7AuZXB2sMapBxPcvuT83Q9BzjGHrRYJo5lQWmCW4DX
LGAP/aq7GCcdisVfXrWC2oa1j4ubQN0LYzJA7ssdlGgY7hc3ynn5QNlteZDPQoZk
DZbX8nhql9cehI/258JQjfsTyIQ/m/M5pzfh8Ohk8hqz8u738JC+CFU28scF55OF
1/M+7H9pEVi/Zb9fLw9Jc/cQ0xHH2QUFmoIOVetxXCODcUm+6zE/x/JtK00ZQwoO
nyNeb9HI7Ocx+baP2/x8outuEgz/82WAXlXtlbF6W3R5T7seWHXTTPhQ24KjUwf8
G9dosyLBoo2qEB+u5AxJ3pdFOq8+m0iS8jAYXh2kxDDHRZocOlFTIjBY1XTSGs3W
SPxSS8LlRxglyN83tN7Er+a5aO9hmdHYmpW6QmusQgbDLxRvjUpyUPnPM0bJ1YIF
EAz+0EgFIUfjWQu4bzuOf9I0rM0f1HJh4OfneouOGs2WoUp+7mIrnS+kBh+SeEAk
8cozdOHQrEhVNk6gOHSh6sO+hym0okSDT1iEIB+FeA9p8Ga/lwvKNMkoY3aLCJyh
Lq6iMgDwki2RIZJZQ6xiXDd5icslFjdkYdZf1wtD++GpKc8IZ8RfC2B+l9ScFbg4
+lQTDZMcCxImpxS0oEbmmlqoB0MvcAtdaiAYuLWnDKEAZ8CW+07W4iS0yvYkcmUo
/ys/YyO02OwlMCaxVW94cZuolN13Uxr2qzxFUmb4yrifdIo6i/i9HHSvolE7F5q9
q/mPPFhWXLJPvxUcDQr59UbY4NYXH56SU/s+iREEUpD7ZWpqQ35vv1xEAjKKhG9n
vMHRSR5phcrQ7OFp+o92aNp+vuLE1mG7Wm9Uroa04oMHIQg16Qh2W8vVAbb+9sQr
DfBS4wkw3SwmDU5etLY4nsF/9YZYNlx6G8IBGZnTVOVsJ5hDXCTAMEO6r+kjQCTI
izgnZHlKlra1NYEdaEND1XznEl/1bgy8mlU+vxH8ZUSTEF1gkuuUGYJHoBnUlPKo
VLAeb+Ep7JYclGVUaddjp2mHx9q1nOivS3US9ABsttRPa3//SBwgL/1ytwJJOhY7
A2Go99ApVnxKhwqveEw7ZdCtjq3QVC0rtxfZUsptRk2sDnVc7u4/g/AUchfmBeA7
Poal/v67J8qDoEmyqtJ4TiwBpE3dCR9qAuK6iZ84x0rlz6tV9YxiUQTQ2oa91a8n
LwoX1X5tA+5TL3v3iDK7XzwhYl2q3oEmZdDUg5J9tzvQ7qO6Wu+9O9mIj7l3oOrT
FvLsnvEV054w5ga07EBRsx7CGDKLD/EFLJp8QCsTIHYMsTz0Zt3D0ZGW4lU+sQgs
aFsEC+vT9GS/s95Mtexd2sfn2MZqAaaR1ampVEuglidOc231WC3ZpqPwYcHlGFcM
gKTCTd0T56/74V21tckinuwsXOP5rThR73QTmyDvv+6ajnlvW8MzCqOnp744AmEM
2fUUUNNkVHzGiBjlhAvfd8M2cxQzgDEUdN+OBZsJxaYCjHiNmBFFG4l+Hg+QVbWR
yqY+C/D8X/X+HfqrKqTwxwK+XYnlFXjFl3iPyagVfw9+CAlRFSmtzD1ny3C9C9bv
aX5KPqQmFGltyJZasm2S6+gK+xG44XnwqNOTAT30Uk/K6kOYzigMe1wgFjbn62tK
m9+aZJOsgl0Psxf1HQEqwy7+SV6pKsJvjlDL7+PxkOq/TJJQLm6V1UTt7IW5O+Hb
E+jcHMRzDh0uQZquS74/D7QhpHZyffuXxWEHccNnwuToeQqrkDetxhBpAxEsonYz
qwdX/Cz1809G2A7rtrfZ9cbXro55Q1y0VZZlR3hcgJ7oyZGG17OmRuJdu1vMep3O
drcY563sFJijV8GWQgrSKJibRYRGlRqlXhtt2VTWL0nbca2UmDL3IJz4ZS4fd4Ih
1Y35MTBhKeJoxndKVkIXXJ9jkyjbxoLpXIevusah7fajrJLCR/Xpp9tW0tBTxmmL
hKpFlNsl+a85EyRhFAA+AhvxvSUawAC27cue6V/HnDtnMnTKfE91cMuQ3sEi2OCy
nvRW86XZO1m1AGMNVxmAHqdllzFuLbkrVn/hlZ705AKGFH+HB4oWSQQbl9IpvVt6
hhAc2fsAnPEKGEd+/OyPihhu5ozWNZmfamMdPx6QbMVYak1fsRuRE2gUmSRhKJPs
AKyDj02Qvrebi1qn8dZ8fQeU16AiNxiBCCJR8p05nfpKL66OLZd+W42YwoyrUsVg
Ph/59GgqjXCpWEPEk1SH4MvSqGcmdoT3DvTTbs/JwMhgA32RM2YETwv1WOfiJcHP
5rUCD2OJtr9aIz0Y7n+MyIIVrNWCwPmUzjB2+ctXQ+zYTpMSvQIauif6DCllp+3U
YbedAzyRmy0wB7byVngh26c7xOl5qFqV4aEOQpN1hG9FPamU5T44ErHX7IDHofNS
buh/9pqJAFdbY4hDnFtotRZJJJ3FURdOypi/GOVt9Ih8Cqn5Rv6U0zT9w9nVhZlU
SYJ8q4WrDvbGX0o1OTBudNu4L+nd272YpI2s4F4RzinkFUMoVNDi6iuQR+YQStvT
JWBINp+zN6g7NoJc/x7bSg80REnNEe6SfyTKo3XiMNojZiML9D3jcsE5H5RHBUyx
OOwIWRL05KpJtX9eZUd05AL4LdwlIvXjRzsivCfUploJOBjacfAhruPdscMdNjTz
5VKN9HRnjCXxnrBCh1Im68EkNrD0UHP6OroLWMKIwzPwn+pUnycijqP6CxVfb/+r
ifv1SmSrr+OV0or1KAkY1kH13d9coWapse/xZ10fTdas8sWXf9U7SBzRb90o7LaN
BHR3QFDhb83bFcLKUwDVjDg2T9xRAH3dV+zcwndVeXPkO/497BMkZ4f+l3smvGxC
Z/FDmCU44LHyvHBxeRvKP3guQjom9WqqPEwA4iPFN8HrVrn87pN4SfwmZlf6gPhX
1K2LyNPbhuk43+1k6fPpd+1IjBPe3liLab3A5vPOLkWnaegOjzMujNO8AHY3l69y
LXeQjYarzzMJ/yII85/g9ibZKnO3ECdEvFKWg2r7n4L/5zoFXeANsFo90Y11hJeo
7xhrGFMFi3zG6X3VrrjLlPsE8vDZgvs1errc6wloWQZ1BmUX8pSyzyj9VS6T/+ds
aehskDaJDKEYThS29VuvdB3uKKZAvrguvBPxtvLapfquJvBcF7ktBPgCe+FHV82U
TJ7YmbuiD2mScgcc72QiOWNV1WXrD1ZT47jzdkokcWABuo0g+GD1I5nBAOXn9z8M
4Nwcy0Z5z05caEQsxG3laVyiFCe22AlHiWq5mALD6FZQp4S3m4/rZIQ1/+I/h8FX
79fPPz9HDl5R/+rt6W4PnLrt1bVsmJGvXOCyPDa9Q4EkVSzrrPa7Gtg+4RXze2zl
KHFCMLWDXSKhGtjg1jBtoc8nruNckLjmSc5DycJi6aG0yp38qmKg0JSvPREkrvBG
Pchr85Y6I6Sag98RfPp/GR8ag+Nv5Db0So+yI449MW+9XK3pWxYvvNoVUesZW4mA
PhEhhI54DM/yc/qAMIC4aWVK1zqdMf56P7nVYX9bycgz3YXgonNCAJ5558t+HPBA
KHjjRd5nlxc8fxdgbP2m26KvjAepgHhgIDb4wWgD/iAw+6ElHzI8zittnVzxu4I+
aInW5C2qvql//4cGMIAH3EW9ixVk5LiK6M8QWfEm8Zkw3l9BV2G+6MyRPyodmpnK
Dyrp4yQzCaKi6/ZGCAmbZe+6LPT9Cbc/OPvVDJowg3xBZY1B+Q7+u/2ttB+c5iHJ
3K7ifGLlcxUgT2uo61E9JUn14/4Z23idLB94CGfjpLa7WdMM5SNtcISTq5OTzPbd
La5rJEYex7tchv6tZUkgBmePtQVx87l94an4v7hJHITojjMf/eZKZi6wOaGeR9px
AfI7hPDSxA4pNftIyOroWwbqOSRp5kLOgPVz2TdF/Xn8y5jPpHA9wf+Ypxly5Fn3
BHyvtkay+ckUTZmAj8CM2KwmPKFAXkARKMn0czJyI9NWDiXUyB7TROVVdAItraR3
kWilEGFY1op/tnVUAJYIL77xZggLGkLWXzhht7efWrJx7fB/wIaqPEz3ZDjUuN5M
UFGU3b4q+J5I/jv9bay3zmtNh4r1Vlkkai6DLoFU3PgxJIc5HFYX1qeGUSu82eZp
6KHg6o6Il6IlW4VV7KdLwLUo+kKXXEax//YzvM7xc6Dzr05bCCDW4HUFeBWF5jvl
xiTs82W8P+vmwcFRHm4/lMRSWA8y3kCpXNj5S6LLF92z5quYE5nDlrJ7pJvau4E8
9Uw7cKv7CjGi/3aVczAa79354GgiHyIMfNKJTYYl6BOQAueATXk/ggx08Iige/kr
P52uLqODmot66e81lK6o+xBZnGYVaiGU0YJaNDjzZyPDupy9oIb3+U+Ct5sRhsOB
DBDOmh8xgFy7rnb465CSe4RkLSU0PFu1QidKZ9chbbz75X8LnkdwwT0fRTv9IFom
20xz2SN2OvYcXlTaGRj5v7KWc8ajhQsoh0T4NMt6Omjp9OWNQ0GGlZLw+JarlkAq
oMljsTHVJA095y+9oNfgEFznSs7e7c1dK1/VhYKZC29q0HLklggWtJFEoce25iFP
jWzStyuZK5RjjFUihywBoArAzi4pQK7NtFtjQCjq4VPCyCgiGceIk/VtnEDEroFS
FGKy9FJjlWOVoIHrzqOgaoKKERHfPXSzcOm6mXVPeUimyWyicVqEAlnaqL1Kjr8w
RTEa7XRYosvtBtCb4789W4XfFmommtGSeY9of809g/guFfEfsMm5DAvTEIhcBZXt
lAGzsKeo0o86opXM5x4JegUc7yXAixZQuh2NaTtWMIjie3AoOrcIOlxAYvod0x8B
AaEW6V5jV4RIre04iWncTOFlLxEExjL+G7ageBaNdTxnUwfQeXRr4a+58EkE6N1F
zRYJ+WVlT6EwCBxi+XDlB1oEVPsMeDgoXNammztG9Rb5mlvaMUsf2dgRNGN6pu48
haH1Jisq9CYjMjo0v4Okh16T3cPRN1nWe5umqnMf9aCpmPO1Vv2pyYG8aQHoB4MT
QO8/Ac85Fv19PxFkR89Ofmt4fkURQveLnmH3V5bwH/nbrhFz17ZWFj4rGFP9u1Vs
D59KWCo+2eoQzlxMkYaI6HhTJRblZ7zDb939967KR1mv0/EqfEwlcEDK7hCLCEzi
wPCuBIuLszvqxuUONuQPk1akYrBHTKRJrE5iyOoVsc931Us1LavTDAJ3xx8u7lpA
0Co72pKpD/D5uIneQ+8LenaiZKmPM8GkGa7nbJZS2nygpnKkfH4kXfDUELCFHWZm
IiPdnXxfwKEpbsjOOGlAknbflSqutYTkfJTbj4cXc86Io7k72TkxTolEPeoE/0FY
ep+jcD6dOH4D2QmHlukZv9ExG6AfkaOqW1SDl70Fw+uRT/yH4ezOT33mxhI/kYUj
Km5wUl8b0cR9prM26RVZnX9f131Omu+3VOkPm03Tpr5tVy7jaaUZNiuLYDur4U3M
WW8TMW88bN4Vx+OkrY20Q9a1AEDigMd+mfocfCu3vF0ocZq4mWuriujDsJL+xzyh
s3r0mfKDo004v7g6PFRhVoaypQNBhWnABXodQQlytPIX1v7VXk4ZrTwWNWvy4sMj
rAT/2bdvVOp4qJR3wbuBx/0m9vITfVYcHFxzbwd3x9KmrK9c/CvJl+a0o6N/hqMe
O6bYCtBtjcJ+NOcOpiQLirLi5LLbSJydIsGiUUibCW32oM30lZe2Mfl84nPBuWVO
YrYbHEjEAPDFqZ1iZuvCWjnjyIFaep81ya/XHL6r1tX9kqd2iUqwS5WiPTQxynJY
yUnusbaAILpJU7dxTvgU/N8CdX+hrxoXy6o4uyuBssfANDfFIyDD7qLmoja9NSX6
Xm5CdIoFvKalU8tfXWAhh5GUGG5I99zbT/YKP6SNKKnNMr/OgTZp1sfMkma0z6K1
t0dSBJWkGbAnlZH/v25R95Vtf/sqmTPYl3+Ue2qLbSnXbhqvPIVhbdsw/csfZsKY
i1vf9pselcP8NYzjjYzkgNi0djLU3LMWSZ8jzfjM/yUqRrs2HHeW2fG23nASHeX3
UvrmcbtbciSMFjO3lRLgfLXT68IsaUvPTE7uYdBFgBAgnSA9U0wnImqH8qh4a+yI
9V/dYODK3Ym4B6X0J/cugGUMUKPH8s1rqjVVgFGurt/a1TZ7Q5UdecBCmbwGfbrC
x6YGeUJVpd2Z+PAgZkQyRL2y57v2//CUatXiIUdJDh0IAad+Ahuak78OwSOBnBoK
pK/X2ciHaTNaVlAFLrpE3CnLJyH3TVueuUCLNRQPMNLScRBf9DYNZuVConzga+pP
povffEe3vjDZA9RK4AiznQ/t6/chFNQ7CWfT50uAW6pAGj/+JTDMw7L5B3wXPX7P
RSxdJrRQ1Dxp2vAd7NS7mdB42Z6QU/simHwWipYirMSDlISO59XCT3AdjKVlB8WS
ASdBWYMPwtkRZXXp0QNfpCdh/Ar6fMTec5TYyk3PE1yJPfon07eDeG7kgh/gPfXG
iA9BH2UekkOftQ9l70rhS2g4xHNY+CMil0VsF5SX+pLC2S0oVRisSW18nwkMjJ0U
VGuAElq+c0bu433VpdKeVnAXqVlKQqv0NxPK7GXUnBQK79RqznrxSpYT6xlV1CDm
2P2Wktt8yx/CYK+o9QhZvRBNUvIMi+50O3gBMLTP86HHF61riVak7fLlzd7HfNUM
lwtYzbtG6ssmJ7U8odXReGnfbo5PHZl2zLnF+njrJw0GIKJk3WL58W/NmiVLJ6Bs
2vd/TrqOBV/kVGWbPrpEjsCwB57TMVRcUMd/K+EV2/KObrpSYCH7jj+c+XQXO2bc
SzU3MtZ7yLf26ZtWlP5pDW4riD6XoIYStkT1n2HPFlzZIGsK0ZN5SkR//0m0k4zQ
uRIa128ZcrBaURqc695yK4PmqYor5cHG/KhHiVAedf6T6ZCOvNHU+DrITCjrTad/
jpg6r+ACJxclXrggQGOcoE2Hrx+RSJoa8dnjuBot9dlbypRyt5HdOhEXPUpq3Imd
ty/L8EVESGvvAlB02Ev0TIEkIbOvUFi5SaOBFXo3G2NEHUVuzcIDEnEPohN110pg
sRaZnneG/mQi0rpjZ7/NcPBC/uerWcHZHi5W8L2lJjXklDgCta7Xr0d0k8kqW5ht
HB5uS3RC0C25fc0U2VOlk/HbxdUtJlAI2drF0N+9jM60G7IqWw9Prl3xla4SLHl5
aaoBmXdHOwT5tnr17ReEQRdK6Btq0uAqhNA2q5Wh2Z3OMF/W8T+YazUr4dSs0NiA
RtaO+O+6GMfcn56yiAs0GxFoDB52sOEt/RvTpuqbribWBAzzW1ug1iz01g4rs1a2
GhGzEiQZEYR+0ZD8y52/mTYeqmlCa/oaJ1bPbtj3EElN+fAnYQONuvWkZJyy5jm1
bAN0Axvr/4X/IJlSK5imT1fOZND3f+uX2cdAUnVotikwYJRWLR7GkKuCS2wWtdf7
bK6PjBIbPQwJxL16CBYar7xESRDnmA/nKz1G673LAsDlBkASUqiB4FCM1LMipPsf
X6pb4Ni8Nka4Pp794CvyCUiN7RCTV0uSJyR9BUBtbRQJ2IwnTSWV8+bSqJYQJ8sg
IJaZm3zxEDZbN8+qKMaSqEuOZ54oL9unjPglS7cf+q2GWpMuRo5JOCe/3ok5AAhr
otUfF7+KhQTXYELgTTviaC6X0mW46DzwBejNnLh6mGhCnokqw6xZew4PUuNKGrh6
xYZ1c5XTCuOZKbP+ISNbTlrjlRG5lYFwEKEY+Q/v0aPUPLVr27naOksR64KtPBft
BWTnZF3Cy63xdz6R7z1IO64Ma9Kav3ANyF9SCevkPDLBwVT9k59qB/R0q7LAGoo0
F3x/9VeZ9MSXOrukNYqJIB+CojStkXUligc5lLEbbE1rL+CPBSXu9Ej4KX3UCt/k
4NOOzYFazI8fj7lrJhkhTEVz2zZABMkt63pvwxLwDrrrxh9vlFuh975+h3w/KhWz
HUdGLTAYz4YF6ZljtRZJfjLQe2B0YUqF7KIcl9kc58oR1kYPk6GPVteSI6dZOOeS
Pesjv6R8kPhq7Dr3pQjzRgblmgPrH5/8HPKGIiYaqJkSOXRLhUhWUkHW/rfvZNr6
a+C9nwPJOFKXxh7Z/T5fQMGncdY/x6WnivKj7fa10ZFGdZMdTCjuXOUewAALl3km
OLPgUzsohWsEnfhkkyTmk117bWJZYnxZlTTF8x4L8zGbABdyPyxrfAWq9oEWaZAt
P1YIqnNMsWrWFgG/lRLrB9PRYr4JNAx04k8gC5J08OiQTmwgG5ic6HHceLIetVOx
SSyLuXgkcARaFOf8RYfbxBBZojibVTku6xJ0ODuRV1a5Zn5hfb3EDQyYnbiJL53q
1lDHbRkAlqjSFJNDE+tmR/SYEqM5CEMJns7lHFPR2VvxSkj/kG0I6pSU6BkGF0Yl
CwAW3VNlCozZosBGDiTxiOa1CbAlo1CvJIFnDCiHJt8P3WBq4bKGr2TlMMQF5irW
XWUkC8qhmbgCm7kGvN0fw2GSedhyAIKozuahrqL7YJXDJ5e/JIsNptvy0m79we0f
IvFYKdpStXjRf74FPMF12QqZ1ZyB9/RpsCp6Yj3la8UMsOFfvJm3lW71TDkMHRNT
62L6fy+Z7cQmcMwz2rNPMRGhjy3A6qqFaCmlXZcMIy0ikiGZmxlFwVjUqlCOBqu+
4TSsabMtXZBWrgAJwRkkey5lIK3LSQcOM7p7gCkfK2i0vyn3ERJAeQauJY/ANEpx
dU4j/ikiuampNVZYO64Gi4cjWq8h8J3TEPBujQF2rT5yPfA9Tw08br1COP2Pbir3
EUaCLtOeg+E34uo5AmE8qUNOJeKWeGBQs9RIDOEAL93wicR68ciRESeRYmRkcKbe
nnIz6CbFbtGSPcuOY3ybGbceUGHZeSwsPv8TPAIdQx/C1DPYtK/UPbs2iG45YN6O
grS5jUrpZxFhE+0H22w3f+XcaLaR2Rs6FTcgRCLFevPlDYIGDnWt36k4bPLbAIFW
GOhzre2II5XA3kWFzQr4tUoDtzurctYXlJnmN6aON+PTYrE+XAXXu6FtP8qweU77
e7q/hdJBnbo/vAOIbfcWVHuDwaCJ738Lf2VWJM+ep6B4Tn4jAXoYfwqkSEvTuyV0
3znoCgC2TbsDCfhAsJi3AhVqujrDtUTqFw8PnjfB3OHE1HKlHx4hlRR8B1i5yDlw
mo5ZJxWXkOwHLYEz+hFgaVYP4z9U6Rl1Awe3eN08WBJ4xQyFvqI6Kyr2aJV5FbOu
LSlwzez+EXFu2bL/lqiai+oXt/XecfH1/OH1aAOeAGMeCCwhxtTfAoFaVbx0w+Ts
YtgrHnO2O0Zet3LGxb+KE5b8lea1nztsJUIq1Fb+VWayHsi95/KOaPPHoEpDQibP
4nQqaQSOYCFUnssC+tG1DMcLZREkwDuxmbv3z0Zdp6CQ74udmVMzheekFLd310T/
Kv3zEBxUcLTPWPmFYCBn9Xj2v54GNIWTGJakS4FPqZSbShaGdp6x6Hu6K1yAfSAR
w+x7sJD/CZYrM7vDNnRppnhULBjUswE9oV7sAda+XJTJ5iC/bIGMwjD4SvLu+MtN
TZcvH70o0xyvZkHQ64RQaxyDf9WvB0Yvb8MwfKTLQdbaSpzT3omWb4KaSnSLddPu
T1qwoNWsk+WkUcXuxZvwqIpAIrOVI587ilazXTFtnSQwlZsud1uoK2C5wOTkq/bd
nw82nyJ0e61VXcnWAIQQZ5/U4ELHP+ixrqD4YWF0dUoguAv51tKn3QuF2OQZQfrj
67QafwTyWeQnnbI9aLNlmvhFaW1cx06AYO+6ERa/hiXMDyE0Id34oRrJ6tXQ2Zxo
5sirwJbKcp5V+BUfYId2UN3bfLMs4q5CCUT5RdoNiDaZd5WbmJNmRggvB8cMJqvB
X/5crbcWXJkOOnQcE5KIF349oF/Ezuu1ATloGYvozSHltRsfAsFQDeGRyxCHcrcZ
uNKhfFUK8SZqxuE+yjkxrZ14NeOM38dAjfnhknqf3uyI740Xe1sPiItF6Sh/6C5J
MJyO29XnWUSWD279ADA/OH0a3x6o4Do/qaAWAkSWvJjyGGIWwzErN3SqRBuVaWCV
1A/MzHaLTtxx4vYWIA8YNF+6EVs585xHVUGDflaEslWZXso2g4IagonGDeeqmlsC
vbkjo2/oWWj9CgLK9fV3tAMqNb73GSIjXEXCTm12O/8E8+QgRmzlJ+cSZm9JldaJ
Eu1iWg49RmtTo1YOHAxyEoNATYvcDLT4rCNBrPnYvZ6+DZ8RbCnFCu1vSH4TR1tX
uWHGfcbWDG4jGlBhSq2YerdrbfdFRIwY/F1fqZpp+x7YCDXJWvVC/U6o3JBjF8Do
QosIYd8FWVOdxbU3nhec2H5dgq2W+C1eIUZ+nuXtSvuIwshxqsnpzbnZJjmlMzya
W7F3vv08Tf33kRkdVejFIXJrkrqGcCAts1XWYszNlyl4j5XvVIfc+ONX4HTwajUy
Kt5WD+ChCd+0uckvNqqh/HH6ZKnWKwbWCuGFsmiFv/1hawq316yHJmIJDUQCPOkP
62sSgpMGFDiObPOz53rUXctKI26LnsQtmfHAEvu503MvXxZyJgAIfsAFRaQHNKoM
zFL2lnnXN9TYfaFtA93iGWycsyc426uQaK2HFi/2F3NYFkXzynd+xCzTnHVnOVY4
lHuZKVjm3vYR7gAXyMT74jRdG/ybP4d1SnpjIrNSSQbpqZl+6/0MnpASwEifhbUp
+FZShfE806QOgmFaaOS88jJ1FhQoSfjs88BRH4jx/NW1FXIxMQNYQKVDrjbbb06P
meCJyTsslRSESlXgoIsk9YnaHDnK3NrC343I/FMu4Fv8xun90CBmHHEmfgMlz9rG
VpTwyJrVV5GZcZ9xmAa/ujz/+oEYw2Dq2OiozzfBCt4c/scYkE+IaDBDs4HTNTZ1
FQxPnZAfv5HX1fzq+y+QxnyQUDcAfVxtjHNE0GgIIG3fUjsu1y7yVT26LhuwhK5J
xBFAc5jlUYAI0zjcgspEk98syH4YuvoSDDrtaUFPB4FC4FOuVVFwotzodN+azTeX
p91HOFT+ri9gMjoq9ps7KnYBAKHqlx7lp6pny2mp2Adw6Grv8BpL9zwnRPWYZokI
o3rqgi3pCHLMwkDgodj0Bua5+ZqiRtWknD9VX68z+zUPJR4QqTd1W9uX/EpfqRuq
hPeTZ5SwlOuRmS6diLNj47b26/jcmvrMiOB4ayLJSwgI/z0ojev65BdHw083DD0e
eZ293TJHxeGSXe1d8t3PaCTHQbU4+eXBgj6axdcmxU4kH72cJ9FETHRKA54qgINA
fV7v4DSq4l3bYvJU22lnxl+Tg+hZv2k8eWmZ5IPE0Xpm0I7lls4+895e7zLCXXPh
dsg7X583lQ0ELHiFqFAKnRxkEzO5ZBfoj3dibdu1dV8XvfbVrqh1T3c3f78OQeIy
2+TdbsFYsoQKixC4FEZX90UeFDo5pC+WzifgQI5+rN54CJOG5ZLMwd2lm20ejbAE
5thjaokr5MMFK3tcUFXq6ozMdISNTXkldFYShVDrxpnvJXNQCtwjt/ZGMRjoHr2f
yHlqz2m1b5Sz6GLaYE7hwOs7t1xOsDYuNyU5H8UizaBprUdgPF614VWSxH+3OyEM
YutZw1kx0dtC3/MN+yjqbUya3+Vb+pNA7Jr+uhVanIOlUF6rEQkGlDnlrKe+Aitr
sgMb4fd1lPLLUKbD/HnX4uY3ISk7qhRg7aB513vOzfvuof7h6SAmmEvxrhKkTC6i
d6VcElzroKpuWfBSkXdPSasmvtB/tRRPHxBD72/SFwRcaXmf3DrreOpQ7hHI0/xQ
XoPkHxcRhijU9ChF0EaMC7ib4Sfza/gS+chBN9kuay2kPl6bN51Mzoox7eBMie+S
y+SarJ3YKKVdpcW6kVdA0SyzqQMbWM2ZvurE5oUn2kY3BOTwHe+mFjzCl99UAB1O
2X1JxEofMsssJgOeAaFAdnd3fz+mma6oPF8RkgMUlY/qVeTNwcyKR1W7h4IA8/TL
zYooGbU6OmhN9YDV/YHS1vTkKuXLrQ0iQrpPAI+7GNY9UnIWpPsOWKNvIIKSdH+h
MdeiGwJ576ym/a7lgf6fdW4m0whFHWeZePwQyOlsch6jG1igRU2dzMcRa5dPEFmh
ogXlPFWB82P46fOGvIfns1RkWs1caoSq6rXzzxTk1Ykfu7kDjqyzc5jJffk8UeyE
PLtCQ/5yWEIwcJSI63S25u65x8ig6VIjcONlxRWKBeI843BP+bUHLfBVg+3Hyuzm
BhIw/MFlzcEW7MlZQSImNbKaKsxENJ5oQ8mead2VgZz4YWzNX/wvQ6UOrhj6zWrW
VtsY6iVC7IoqP8+1faT45yuCaMzaX+eCBhOXW+apgGUhTYVv6MyGw+AZZWFYVhZ8
QzlNgcFZUblU+7MK7rFc1RLbp8SCZLZ5piILgbJa5MEU5ZJH0fNvnJ17zRL6kWjN
Ta7aSE37DciOg2op2QMUd9eaBx2gtadRuEd1xIMAI99r7U+rdSFMnVUdS9eptm5u
QgNJYuPQ5HsBtlI/D4O6vsDOurqvCXjVaqB/aU76vMtewCWdIdszFDJpUuXDVKVe
XLxo4e3zrXljnoXoeTeovsNGmkxm8t17B/Sk3+6uoVbd6QQtHlzjsJnYTiteALWx
pNJebDmTkXJtpw/R+Gl8xR+mAdV7uJBoK2++N4hcacoKbpp+TiSudtNrnMUvW/yZ
R0wyjjMMoTVNOJSa9noNM60wg+cmdO7WPi1B2bC8L6yyOuSufZXxQfC7C5w96Shu
Uxre7DZGi1PMWLGODwb8BP6gqhY0qFfzVnyj+oCfmtuhEH29Bevo+0pXOSkmFKls
Jt3blQqZJdBTXHOo4jm3GU+niMhkqA/pih6BeamOZC4n99GILHRlLujfD4acgqFf
pibfnvX1qyfPtbtpczEsuZ/IgSpZWTdQTmyhHw91gDCimiLfyK+3SUK37oZMLAds
kgeVEV6CgT4SX8gzZGYSeberK7Q7yPFnkF79F17+Vg07VBaV+zX9Z/5GMa/ujKho
j9jhoel75NkL3Lu8+rn7LsqTQjSeXuFGBnXQ8ka5t3kUiMwT8tSLIlCsLvpVL6us
0Thy6e1z5jWsuZs71iyGMbJH7fAHwFmbKZqwcmFFqK5qFgRSnYTXz9IGlxeJqjjB
soOgUh22NccWauVPl+z1t5aatJUL5lcWB8Y8Cn+ceeyuxgzlDgvuKblMqkKKrv+D
zCX22kM6i+i1HI8fF1ZOwMiL7OXZuwMVqB+z7vlOVHM4wOZv05gorKuHVxkqil93
biUXTrf52ICbOJk0B8drEHd74WDdUFAOf3lqLLlAVCp5bIrXRmlAQcRbX/JL2e3N
X+G7L/3NmJ+4EMSW7CY8vYEgFAKdOkfOjhJ2hyKyJwzyPK16ZDI1HS3kPuZaP3ac
8PGUTmN+tD6yh0w5lQMw/cdL/94tLfJHA8zn6Vieu0Aqe46Y/LcYXW6S3pnASMSu
b45zbtC/vrjxwX8R2/xUdjFzEkV0mDvCMmv9mvflokm3u3xyaHu5QA49imqN9+ns
Xg5sxRaMnIVSjNCsFQoz4RmMWIdzC0bF4s0psRBTo5Yi3E2/iEIcDmiA+TlWegQG
VCCf1I5PwNbejm3Mms1BS4315W5F9FoVhnH+7YIMJhjtnVK8ALccFciCuIkr6GUt
lTJVwBPW+UpTjbTcXx4ApsVlcYR0uTJckjUXfWYXu1d5cryX20J/9tlUQ72ZRbaH
4WfplQy+GemW/VNxdnzHm53/+YKgu3UPhqF1NBqTuQb2I6qS2Uoud+YVwT5kz09w
xIwrVM2SAQEw7oLAujQhU0i7YHe9ok69KgtF+xQ6GE573uJh6vrHAh/madWmudME
QweNtDeaA0VV8+Qu3VKrt4HSFW1U88yVvxTlcMC+ySpeNa96GoToywkRebnhInlU
q3A6zK2Qy40/ZDSE8NhPbAI5+OTSXhyRiYy0/hMD2o5ieh6nku16rz6D80vP5kT0
uoKL7Hqdzo2QBnV1U9iWPjJYzeCCX9gdBG9H/1Y36qD1DQP6XGqJ956eFl6pp864
WJmEByl0D8Ql6SCI9md0115XH4MdH5W3afqWQY4M5K6KK0y4yVSeogOGk0ME+x7K
xJ94lS7+dACzzs3HI1EIUA7bdfXygY5NcHoxUBUNiEwIt50AuhfxBGfwso0C3bKf
NqcN/VqPooANSCveU3Io8kbqF4rZIm2unbsBIgGVgVly5CBUd9Cc/cdabGxNg4cY
BvyuN9CXmPZWkOcBrp1naJBLEaTKd/DVR8kooWkZB6KTjsUN+R4R4G+PJenHObeC
onz9snqhoAuB1zEbT0SCan/EGq2iuAu8NBxHqePlcOjcgT54FOeZck6AYbkgEboB
GcO/B7RixKNl0K1rMHQldR++2LIOD6/XTP4S/nAkJ8syZd6h/UlFYpRZN3fPJ+Ol
0SFPszOGfdzozFMmPlDluh9ttIfGjJSt4SzJW2nd8ipdIvjqolszJ0/TvL7embo8
ixuyXUpTNH/fHvl7ZQlESLImxOCd5xQVmacHICxP5kkdyY/+9yP1QrxSQ0h5fHXU
ILsvdQu/tUD9Fb+mdPzefW/eLk+rNfTsaIa+Kdp8BXyD9iGeaADfUwS9R8Nl+FmY
rOWQC0SLG4A+17H/g+IwJjeaNtcpuL7iszZ3nOscaM7Yc8gLsBioA5LO5a/szQl0
5fnqeJbV61s546aPbP7Zpe3qHN5RdDr1AQlxAiqsbzqlvjcbe15W9g9/YA9JsjK6
VZVHACkc0k11rnQBF5W3elcXyKivWRiwITl3i8CE94doiktRrR5AUMcixzhqWrFp
aTdZtQ4+RbM/IYDZgUaux/NymfLoKyjzfvRO1fkWQlIHkdk3RHrxfS6VNFt+S4/3
6JPR5se8ZdKU/GJhUdv4nKFuq35PPppz7mz0CgkE0CdjgZ/Ncu0nmn45I+2d21lK
LRY0mTRqs+2QxAEQyMvN+4ajlTQAyF2O5xRgKu5frS1mUca4ua/1TDUySn8+9ZXy
0R9ccDLMVuNpkz75hfSvD4JM3IjZWyPVogDA5/38VopHprmtTzfC7/jlW25GJX9+
EMOi/YmEI3gxUgt3naB5PBMDdmPD95R42IhveSsYQl4aHlbw2RxSh0iAalzhKClc
3N3ueT7x1RR6VB45MZV1VZXk59fl1L0DZ438UhQFKEPMOBAy6DuiI6zdw7T4X+Ei
tFuQVk4EVuq3/utjSIEZnF9cvot44UkjEp6fojwFZ7zRZGuVvfExvJWkoJDfn+8Z
xX1dB/finqgBeWEMiUZ/ivcjPT4e/I76xO6HuScWLpodW5VrQXQnY9lmhDzQqjPS
C6WcYENHk8OnLZqsVdyLSo0LWqLcXpQ9DNsYMI0eMss99r8OtBULGLtwyaW7HVsu
recCGKU3aXUZW94ezZ2ztDQUsDqBYeqcLgGKes5eBiZROQUj/sdPdluhrlM4S1Ch
t7vzt2VX92+0iZ3D3yZJB9kkaTtd2Jp0V0rOokEg8x5zUMksDnm7ipYYYh1hyfIS
+gR7Dhe5uqNS+CeNifjDmnCnIsQahwV5Ev6UyJYayCO/eBtnRWzahNPpk6qTggvy
/bvEYWX9fH3HFk8TXdUXPTX4vo6HZ2ULEsgpZ8eRx3v88ud8zX1kWc5TiDold4LP
0vads8Q3QI85jnGT3tVm6eeY3RCfGwddLOzI+9h6ZWTRqEYpS9o/wysH9aE5n2uZ
FA1Ul+D0wrhZhr/wse48mNVo1f5FLpR1h0GfyB+fA2Ny+E8IaIWS4utIfTS9JUnt
1QAwPUgiCa6LpXjgMKtcne3RgixlZyvqpw8HRuhNWsucPVBFdqmbW2ATd1KO6FgB
cFAy4cr4b6P559gkhYeaLXec8Rug2qjZRfJpmkDH2vYkAwWCP46v+yQFn7F0Lf1r
wvA85xY4GLYudicVy9wvdslBY/f0R7nb01PI737DiQFR0XnwD3fzjXtKUFYdLxYS
sN3mxgezryQ62CM6e6ya07pYRsGZ+O6NllRjfUbYMOYaOCeQODJuvpxFecXqT77n
IkFHpPmj0CUnsKLLpRrpGh5xzC0HSc1GezWfmwsRpdr+I/UZa96K8naHfE0fR3Mw
+U1HMm9jmDxOCKoTpkNnOfIknsvY+ICbANmoPHXw5M5hA8p4ohlITLwztAsggAVs
Cyd87vRxFO6eqE3c7VtEINsqLqvYVlj1e9g7dYbrgD3bBRYoMfGKGQF5dWiv2KUq
lKz+tXM5MYlMB+mWE3tWDqXDGk5vCjT0X0jZRn7lu99deVWdMRqFvp9R1HmordrA
F3e8cP1T3h2F3SsP/NfgORohrbO33/pWfWDvxTigjabIpyoGqM5/lCmLBdd7HPUX
pz+3eJsO9VzQaN9qZ6Qa6qCzDcUj69KCxhbpIZE90XkoCaUZH5TZXY/zvXQhXOnn
GqMXyo4vv3qw0L9B7ZIZPB+SbeJW2UOJarOshpJTyWDUIGqVodJJ4J42/5ZRQmGo
/f9GTe10JhSFNHyX99ALVvY6wULjiWcnuL3/RGZkey8WaqGD13SfP5Pnq2/N6iBh
BiXKaXhmlliTmtCB3tfMCx6hWLjhehP7/bVKrgQVBeUImfVotEA9HPLwHbBaTGY+
8/PHGOtnvf+k0bHMr5tYXXc1pcpYo2DU4fOcTUJxeLYMOxmB66w05eFWDAwvJb77
dlMNp82qsJqbUTZa9uyrrtSkUuRcsoYL+ux3bNrQpvM34tI6xPAGFGQsctaZbkE8
DNhAFL4ljnLK3ZTc1qML1um7cHbSKD8fEc4Pezk1ahrpgeORXCxPkJthMBQgCGwt
1oUO7rtTYlPr+fKRQtvwfNg7r4cKpLSV7e6dW1eiq8B8l26CcWBTTzhBzyR2BQwh
+u+QpqkO5C4B1ru58n2Y6N34nQ9wJyK4A3Laflyg6IDg+e3ZF0ZvBwNSWdy/84a2
i/LvrgdrJhgf0ZExv8/kEFecOX640sT18ULg9SyqdHjYBIzWgREtajkqyHzmsjUg
Veqe1vGarSWaERHfjlaOnO6a40qwzW9kqHt5ItFhgX/rVb74uVkRIV9qJhUpGG24
H2xOOxX/4zeKBSNWiZfo4AiFJuXXDSqSlDpLH1V9FbO5ZDo7z0L1ygB+m+wKOaIh
UYi6AFOme4YoWcLQb53ImgArAJXoHhuv/DYn8O4D6t0o3WdoehQfy+uuSwMnZTNq
JPHLUbIj0TI56FTlv5WbOGWlMVDlxuAe1RHjE8zzFHByXuImgmMU/SCQSXE/QJaZ
AWyCSV5/4nyC+hzSgnrxQ/JrQmKO3q23wKrL6Z2vf2YiNTAXQSgm4t2mgeONFPqa
jmMhTMP996XTyvYQQABqYTD49AgPSHzZY5wO4cb+ahYEAeJr4PoFEhZcBlbfxSvC
LN7kVwK1KuFkLUmUI47TmyjZGOe1E8h8riN3CY8zP5TMplIuaqYlc5Zpicm5s4Ls
uU6JjJEE+l49mpiEka9moIHCxnaD9obTuvee4F6M9zB7fcnPq1SUWN/mALfEIeKU
dG9uVUrzBo733F4jR85DX++Wcl+rJMgXwXJm+AOiXvaNeqKaZyCJSE3hrcNL4NkM
PRe30l+TwL2vXuqdZCdJA4HJvVRjrGXjW/W6ZHt6cUtQSD4Pa3quemWgd0htnhp4
jUllUEqLirIX9eBFwbLYDLfP33Pt6yoaxLl8a6TcFmrNBteh01WVPbd1bUspnVm3
WaRsCRs/o7HNYYPlqI97Bvibqs+79mSUBCKLKKdzGwKDZr/+7LU7GOCK3bd4mr/9
1G39DoA82aP9nPQKrqIiTB2Qs+26/miJfs3H8SqPYW2LCwP8iMF1PK7iw3vLvGmK
7Cl67/KXrK11gdVhE6RudlZUr1e5sCGWBFP+xteHv72Cxn46t5ywYvGudKgPmslW
i0/wvHcFgP62Y2sUkoiZHsKOdFbF9ylgd1ZIl7yVby1k8/JfBoYLwr7M1O5iTsYs
ou1jbJgWX8a9SbDBtsAD0yWTpXbKR+PZa0U6rz3WFInA56sFWmNActX8VZdzEbqu
Zye5TcolpLOwT3gkk0+I90rtpXcbDvtOYFDGhot/j6HAAQrd8DRU9+yk264/0Drj
HIVnEMrZHo+ks6ROx9iLUtUzjC9f2IW8t0kfKZTInYelM2NqhZklPz4vQ2FGF1S6
XjKArOaDGS38aOPyEOqNnsibdK1t2IeeHnldn2u3jj5h17HfBaHSlkmTEKrsMyCW
Db4N0CKg/1lWzZBhRZaj+Dlj7OcG9vuemYwvns473lmkKrUqUlmo9Mf1KSLP2njz
q+uxP5mmTpjqWUq73bsb9B6Lbs6CF33jZqq+bXZ98yYAFaaW/IX/cSBK1eZPKdBm
g1IOszlVKN0Y3SJOyn2U7KMa8g0Z+idvz163+vhsoI2xA2GLVtLwPYC7QoBWnDki
qMbIUcrj8QGsZ7RllO18kn2lzlR3EJs2teKkiYCwP3FspHLhwYr32rC6ka/AC3Tq
pzMqaTbRYlm549ZoQCl6F/EQoeinsN0lAIcV9gH6SDGmc5TtNc8ZUuCjy80SGh+Y
XnhQ5Hff7hf6WH33teS3X9i+91XU+kzpq8egT+QuC1SWNzlnSAZBEqAF/s3hB6eK
IANHCi81zxdcMJtA+LliyLXARxp6t9fL/moEr91O6CYxJpXcqi95WXKRjeRqvuNo
Okv6yeFhdW1u5tptyrS+fDHlX0aw5FxF/QOMDqlIyzEK6z/j86UHhUhlgy7SHwln
Oia5+kicFHET5w8STbMSTJfbJfyEddkRCmOXjUNUDIHvfGX9ZTK9A4Sc6eqP6Qh6
TzwJc4WDkdfrsh4cryZSgVv9ztP5eeg122edrVsJHQBCAjODDHQTz2iV2t3WCOzp
iK/JqFR4OVYomiPv7T0wz/0xKSTHyn4pk+idQenH/XzdfPsy5+3fUwES80GlkC1Q
balRlNUNEBLtqMJQ1N8eJaVVwoSriAvFX71e1zuNGNZiZ3bNRwMLWqpB9U8hl/eY
AX0sj5Ep8dOrHbY+yVrHWjVT0CQHzm/BQtsSyYJCQm/O6UkszPiguv/X04Odw8be
r3bkKMyZL2Ey09OjoYcwKhkyeE3sot3/WkUSScyJbj+w8gjHTe84VCZTTngVuKz4
GKgkKxLA1smsbMSlDxn03qziWkZfrlrmSS/t5TIEw6Es5dZnboWuXxNuwRril8bk
4/VUt/Qcwz1G7Z2SPY4O7EFc8nJFiLlAf78TiX5c27aPXW6nEZ12p0jNP3/WyZHo
dsY8niodAJio5ufBuGtfXsCseuaFFX8heHUa0+GQ76tSBr7T07fC48ShbMgUCgm9
owlm4McyYUh4VC5QQ5aW2ZSG3o/qp2zJ8E+BfUs+X0J+E9FxQAPdERH4TzrAXn/A
bOV+MAw5BXFXPrIJBI5ojFe+Sx+OO3fX9pTnNZcs60nD2uUhjfYy+9LwUpWbz2lJ
0L9Oj+/ejEmFbPx7/MbpA6FZyyEpEOlefAv2oXdC8BHOpEWhdRnx3FXI6MwVGH57
bSr+s2KdkO60DweSaj/bkY+h3j/cDpWIwN35DCCPnJ1J3T+uT4XYy8OQSFpJ4N24
XW4Touf/PtamYiqFJgE7azI+NJw++Q5cAYM78QrMfpsYhZfzR+8Mdd+xTy4M5wtU
hWXzJH0UbobZ3/FDscfweTXlg+Dcdr2ZA+PhymLf1A41EsJZC4KGck2dNtzY1yQj
LD/28hsr0E/2f3BWtX3SuqqbvVmEBPMUZ0ZWHil2DdFxsRQ4o0TKN/hgSea+N5+6
m8+/MVnvGLuZL0u++lu/Myf2Qr5KNfdvQepqnUiPkPK00zanf4o+5OewWBhWMRFT
iwP/BGCawiZ6CrCx12ijsL+NKPB2iiIIsTQbgovEHP1eArkYGuVyNh3omSGq/DzT
dhqeWhYmY4JX92rBsMOsV1hAioohhv0c2AOF5088/jEcTaYRCJS+Qaibyd6l0uef
z+W3eRWdGOCOU2+NAG6+9kQOeIhjjOZYDheT2sol1OCtGpkv4uIfiEk41rEAqN7H
MjdSxNIPw49+FxYR47vqjIZcJ2ErknnnQY0f7u846I0Dki0GNIKAnAPcmHAIFde7
KJpQ1oIoR7wG6Ey1VAZXLlUMEnPmCC/3d27Fw2P/KRpDAubO4JwfO4CF4WyizBcO
pvqwM/uLVJZVtHgLAU/WFAzF8JuJgPuWP1r5OBGo3TybiY1PMs/AcniWn8T32gou
jJsAlnGFCFy3M2uma2DSsJCHg6RS2DmXQ/5HangDKQqnPSFinCIjD2zAlaAByNUv
iWv1M1yhf1sOchWRKA+FZYJ+lokB5TtoljfqerRqaA4swM3ppS5lvv83ktoDLFZF
rOH0e1fRjn3xVQcw6257oWOSBEO9ex51etgyA4pcGO8CEkNrR9c4f0Vy7JKuUoxJ
Iuh22rhCok15cBMQPxRIZ1SPNpcTZeMtTm8SPJMN4ndXjFBJll0N8hl4NHl78s4Q
PtrW3W/zD5JGsfdBt+HIMWdYA1SxAzGfyy2u2h+dGDR656Fw7N2x8WLcLVXMfydr
8qvzFCh22dz4YRIaeYoeVYtF4eZifB9as4cbdSsxaIzoTA6sOJJxcK37leoghVkN
0XDIxm4vqEYbFrQQc20U4g1AM+pbtrlmS0hhNpB5Y5kJZJwe9cFnKgjExUxwitHe
MxCU+UAvKS1CdGuxfAJGfJU2eiBVFHWkV0GqzjXOi2+zFt7T+MhrS1nUCOO72BCn
HMlnDZFlXxFiA4HpDCW78Gv+Ts9QQCkuuHSGs7w1Heym3mMPXvDj0TKtbgcrocGE
IrKg+FRE8QfSmyELVWrSzzrwPEjsjUm0CT6mvl8opqR3wUEOilnqbrTEuN0iktr8
QcojdLZXVJ6iudJbxgYHLIWemRdvmmwd5i2xP/fnfi4J1AmKbSI7sSlcTVSa7EmW
BXsvc16dQpJfNjkCOexq4YKTmfB2mqBS2yQ+d6t/AKS0dtrY8z+kJwbUFCYcOc/H
9NK/OrGkOeJC1pjpW0krAZfE0uNl1yjC60+zhoF0FXAVUUEJAhG4sEZ5j4ruETcU
8qaxkZAbMosAJL9E4wveEI1LGFecRHilRHXLSZLyTZxM7nnQdpGSAkTL0pFmiMIB
V9jAqb2zkb0nArGZJRNx7a+zX4kPCHaiQTpmWx5YyeaPXiKkCZiSu6iYw2oPmJbE
2igi2X1YFheYWupaFkHPPGMO+V/sdS9px8VlzMwwBlg0I0zOhmavCQSAg4UdUCZ4
KFyto4X8hXRESDnS3dfrqQiVsZc/HpSM+poJqW24tDRJfzel+uq3rJUryf/W8xPb
XFL0t/6pS2+7RpNpUpg7cyMDxBQATMVN4llkiy67baJwNc7bIPpcO76qrX5rYr2k
WX8AOlisrEY6ybClAiq1uVxWpCJtHTVxkjU/novrBJPPAL2Ke1iRQFUKUcHnMOXs
7AzsKM44yla14KhpV2v0TWX/p4tiRcpLOpyVpUjMmbn4B7PXtw1y30hH6iFh+GSI
O7GPXj4im5RhzFTRfIirki817h6i2cuc0557+d+ouEym7It1xFULCn1WeOlqF1hb
i1vID8tUV0w9Zp75FUTkNymwrlykudjqPJ4akXRsm+rR0yHL8HLOraO+9XPa76dN
wzRQJjV/KL0eHadJUNTkCdi3cMbcrJ9TMpevMivjsJJ0kkacGOsb2uwifxbUr+oB
VWjuBDuwWp0S2NRQGU0eNStn/Aj2TBW4OpoEltGZ07t81FLMEAZtrSq8yDsh+QPs
kZvbMCIE9fpOkCwz3ITycsz198j9t07nTb7TLH3D9bh80ZLZvunmJNuA59zjzKHS
2mg4OyBJy5T5r1W6h9+CIb4upjyk4oPkhNTjROu0zlOyZPfZFBoudUNNXNQvgKIW
1c5mX4WNOPb6r/0+Pa/og31W17VdglrXUVcfKUzISk/j1EwiJiPLZmQ7jLXnO8uN
7Ft72P56hmaT2mygPAYHmvqsioXfQWiZgCQJ/GNWzuHD2j8HzvKP+TKxHGxB5VUO
IpAMS4WdJFn2OTJqWsy9le3dc5wEvVdsUr7MLm4JwZmyJFj2827fzTe5xbYNQe3L
zHwjz/LCp27RAzUf2fJUWbmc4gTnPJfxMfVU6Nr1H962md/558QnRCE2QJb+mGDZ
4dON+j5ArXyepq9ivQBtYrqHvG9Mv5q+hhkiNwpjFEtO8XG52Mh5uOxsbwqsTbpw
AFe5Bu3zcKGBGkcvn3wjhCXw979cKrzoMzS40L2zFFJJHF1y1dUQXwBl8RiVVGk5
m+DFPk7YXWoAQ3KpSeqNa0znPDeT/eyQhMvMu5uO+YUGarX5Zo3jOIUUrffmkfAk
IMDp6CPWJeJHZ91rHghWamrreEHfI/PnDku5ZY2g5p+3lU5zcxvVrarxxXJeCH3x
PQZUu+VJgJlRvR5KYqAzd/zSFYGmI/G4vL4451f7PZiDgJTWeznsu+J/D8rLBaQJ
fzMk8buXj0apSLB0NM64TeorJ1PCpfcdoNoYQNFKLYcS6d5cJVvRIiLNAdk9VDOC
4jAomtnTSJ/hidtNv2x96gm7NW6mOZw+bjbPmWBazXS4dkw4s538ezuNle+BlY0T
f4i7c28l98v9uScyizmCi0peryM+KNQbr4TreFKyVhhhCxeYFZZ5R/BRnS545WTb
IB8lf3eUKMQZq+WWQhm36BJqGp5jiLzcPKjsJ/NhwoaiiULQSpRMxJob6TZ+54VQ
3FdANaQJfv5yHWbwc4OVmw117sbQ3escZNMnBG2ga010NdNFThPDYOyoesDQ2m8S
tTnwmRRWZ37dAEDTirNWsU9Jbh9y6hAG7FCmyXGhN373pjRbs2O0N8w20596xv/A
MVIuCMDWQ6jiywpLCkZcxtJ3wGP/8sbctcl8gnOILhkwW7pQgxTHkC3mp/d99Ia8
dVqCcMp7r5S0C8uh+fm77FIBZ/pMY1TgU4pdDcVLu0Jll72vC3PKBYAlkF1pZOj1
lCMAWmQKTE/a/FPVqsQZOHXj8zWP9A1VyD/wygTPAdzK5rZv/0UByrtxAjo7lqig
axxH04VKSRBa0TDyRm8pJRhzLTuCNvAGYhJ+xUHHOOUesDu/IJb7uRwdZ+Je9Nxm
PanmvdU0rYqmnCB6CrKdP7ASQpigdqbveBa2ePY7vfFLYgW5t6DtehADggKLQUKG
pdO/786B1wJdSXn1vAK+D4bWWMvv7NjgnG8R5rDS9nu08t0H2PSwmnjegWUJH9G3
BD9xfkv3+VXZzYkWNkBaCODsO3kA8asoMfYip099vc1aamXPi3U+EbhVBjMAZhcm
PF3v6yTxC9eI/0xJtU32uVv/PcT9DHMSJzqIF113bg7si2A0oJIpyOQdCzZtG5JC
FMIIrfmeMj32PlyDmgTPD/GoDgTiqGtLoqa06RJcS5DfU7kUa1i3nRbsfIddW05k
eQgv3kyT2sev9neAZKugG386tWz5e+DvVTLRS7NyFKeyiucz+lI4g9y2zh7fX6c+
Qb/gnBpzrOn3uxxh40BgRJCKpb0hyPytJBgiMZ8Ss2IgzazUMd5NPDPm1v3p16tb
+fTzl+1PLeNlVwLQ5PK1Ffl9NYYyOChNP9Oqx9bpWM4PrifFmM7eV1+gEpClXciZ
lbneNwpIJnA5C3hqMwHpFUz6KK/u8juxWapIblj27vceee0VuTP2pVOyhM/VBmpm
r+le089mfzN22IQUjts0soaqFRc2dup8TECz2DAziYqxAh2+5PxJKfzjYL79bpay
GtKKn5f0bXbva5mMjT9cCHRL+sgbkXRUQQh847McaoEoxdEtU7wUG8hPAumrAm1g
fkPNXwqdb1V745rQAcNCf5Sz5elTTqmVeTvlBgje9EipHGDUsEjjAzuCL1DSoaqM
qV0YPD883KL82MtHShYqPLaBM+Q7qzcMKka4jkrENWBqARGJgLpIfLlJdjxGCLpK
Z7RqSb7fdDo9FkpjIfM4BWzTNfJdhel5nbzAwA8IIlKNKS8zuHzENgVRLlrK8NCw
F7yzHxpXeLwEYNpum3EpoFivNGu0oY7t+dndb274sYZoQ9ghVkKqZX7DDit630Dw
n0Q7BzRV6mzioNY8iP8hYwFqXQD1Xuog1Od6i+frJqILE1QzG4B6AGimlxRr/5N2
nOUULA9pxo/XBX/eqIqQkyc+MsKgtTnmj3MgNT7o9eGWoBlotU+WJaRdBHNW+u3j
9qgczX4KRPztDOIc6pO1RfWSDGyrA24HpAWhj0YPKkiMAmZ9WPxsu30j0t4yewdG
UOLCD5sK6baTbB2jomc6/xYtGf5xM1cDD1JLEy/SfA6bMgGIPjpVJ4wGxz41ZiKW
ZFfItr4sPJg39YSO42DdWJ3q8ic6/ZiYXVqjN2C3XKPTcs+J4+IZhDtAThRLGYv5
+1QUO5FJxat81NnErdu7MFZSBQvjlOMJgARIceHpMvtJIsVBjMdHT71ollPJNF00
oKXJ0EMgex78nhvF0AfjKlAIVjy2u1pWIi1j6CsDfAXNaFwPMy7ai8dQFdDihZtZ
W8xSSaRFtthm7z48M6jDzo9uquNOGPWFdS0KbXvtfrzj+mLMv91gmqethjZdp2sb
2B36OTK+BQxsIm15rXsMvlnCXKwINLltydBhKcpIv71a0pA+Q6iefODXP0TGla6k
ooXmPC34SeNfvZTAdR+QC6X/4bbSm0VIiqDlcyWjlN8H6nbkzhWZQyPvk6P/Hiri
VMQsfKDirQV40t6rI8vHng6Gn36lM8K2iIcSXWJ/0TNUcmKrtVz4/NyTNKX/Zb8i
pV78IbZnMuEZDH/JThHXX+efcVY/qZUUCJ0Iv20zx9kZud8DJxEiFkCA0StjtEb9
++MAShdNly5xnZV9VcXLNVO01xEoczQkNM5025F42OClibszEEMIvtU+ohS5X2Am
vitJFIoMa895jB6+Ee2jC20Aws8sv5VqG3dwLdyQkrivP0ttr3a+dFcePsdxTrc4
UINGbH6nUT/L48AVwpRPGBVIbwiKTtgwl6D79k5S2Lbr1JB7ujVMMGjsKGV1g6hs
atOdCK0BOrwDJxhPN1vNjj5xac8hd6QPB/sgLvlOyBY/CWtkkf3HrEKj6qDgvP/X
Mzim6Vcx9/bFUwgUTyMuygcuB4QoSHWyeB3OZ0dru58t0vWYUMIn0UZZ4xPiU7a3
NfLfk/H3rBhwBva3/Vnx6mY2ngPRYsG1i+gED3I7cBRkDiPlDP23y/2ZYDfF4jnA
mlyw0fSGiW1Dr84cxqsjOwdS+CvdyXZf8WhJ/iEuYC3bDp4ofM0/PxMWe3g2sisM
Lb5gYzNN/q8WM3e68hc5BOKhkJlOF/jBBTpoyg17AI/W8r7s0W7AiDgLBg2pgc8w
/NbfifUbDId2xdrN8QOdWmBCrCnsXd39iS6zdmNnl2vOl6NPGIkCZDxlfvSdPHl1
N02AzSmVVM4JotsAa+qbZrT8m86tmWvyaVN0fNgd6mtylYhYEVy2CYiv9SXAFb+d
+wzK7xH2fcPqjApiUPEmbVV1D9awTpTDmUCDr5oMd66B+LnOYCYejd3I9MtTGkFG
lQHZ2jubURtX1w7BfbPHOoxQkMYVT2geeBRwHD+LFJ8UT3WC/a77UWNa97EnLEXu
xIpkzQ27WqsPGcPyljMkOuuP7kSWGt9bV7ro/I+ZWE3/eJPNUDNGf2OFl9ikoY8n
wC0KtEjNDAkRNklwXXHAZ+lmR99DdG499egl05mPrMtysHCnRbdww33sQpPMr6qb
hwbwgc5R9taX+a/1ypUXAi2X0XUPMCDmc9R3YtywQME/niJdjqYk8m8aib/IIcay
eh02Vo4CeGOax7USj+TpI6U465T9LrCl0NIyssMpkamsp/DvAR8iXXjlaVmb50GB
qt/u+FyrGNPod7DiV00jetEAKIJwFS0Fk68kQfoU4Jl//sD+7LuIlpoho8AQRDEN
pDJ1LN5kiLeDEm/PR6gbyfs9TcsOuuGf+Hg0pNmN4N8J3W0kEL5JPN1y0jTdEgpb
pCJ31K3nlrklUqBTZ0ka3W1tVMavssG3PdEEPnwP25Mz0dVkViYEGYjoiSOMYCZ0
xpigsMohQ16OSEN3GlmBfyCEelDAkBOJmtznjxyZy12NtZAgOzgYZd6mSn36e+ga
5vM3yobdJBZ3KIYIsN4RGCShmRByHmem1DiWJnXPrAL0/J4bEv5DVY5BpsRBu5v4
XVaeyIXU0B5052ZvNpQ7j2F8yWK7pRlNpQC8oZMaZ45bSjetyHCZx2YE4BLSw8k6
tZIha60kHPrQRLfS+k8UfWXzYxvy3qw9h3dp8ujWGQlNl49vfWl4WyIiSHSKhxBd
b1KO68SpD893sfOZHy2SgCNVgYjdZGIPSD+ZLJF6S8HGWGxNQ7vmopSiJFphdxMS
7wPvzIET5un0MHGwtFm1fDJBETBYV+px9gsZYGpeRTBzO0fHc6paeFomabzjlYbr
PQd+VXGQ9QRf0EdAoyr2BpQfT/Oj6fmFPH82xReC7NguO73y/clXBuRtf/1yaOKI
R0j3u13T0k8JmTJAEGzAz51URmdfwV1hjyEhHPE2/pyUeuOv1EanEFoTIubPN4ni
WU/2k/nz49ULmEJJap+iqj+eGSjyKakkgQlLyCEGYlDKPsKYfiVWoNIC0eyFBZ8M
EPQK/mDWqun7UsHvdv4fhWVdgChe/YVc/GlzeWHdo6OhYZczutDnET40klSZGTAc
Is5l1fmBq6ytGqdRn0AaNZvawLxxbwHSs8trPFUb8FdAviymtddC9TKWjWonjZOx
S0KGMHBuYjJW44rArdg9intYGw9g0Z++DpB95RUsklI1fYTkDy68vsl+1f0ISGuf
upQYWwgzUkPK6CNj3cW51bC+V8a+NX3WX484jvRD4mXYps8Pb/r9xMqDcdgYIlll
2wkJT+ZEbMUTE6qLoTbkaTRb41lyjyXaFIbJaR9VA0gjjujKNIeqZ0/BPK5FUvxx
1Gzi56PXfjVv74h6y8QN8H7Glya2NWe3otpjUdz+QvY61MD3mroagZGYsKOvLASY
FpbQtQobVh4Bc4mtJqDjGj0RfN1C4BJSOVh9F4qvfg2AUQOFgfxNqyp6XVGIVtU8
VPoAxTGJcuajzbmq6puIiMlMmOGXAkyL0FR+mhV8/OUxkvSMKY/wixv7FJ+yjkCx
zyJMFRMvfH3l5UCU4GBYxfy1IdsbcmBrWbuRy3pwjet+97mGQraMwSIFrWDOCLC0
nAgDL5IbTEdOwRPWWlYVIWkVp68wftnFjvb+yHlDhj8MW3yDGs/ljeMw9taWwkge
5D7xOoV0oefIYDor6i9MC0XiqGiDKJjiuvqxY8JCib0Bvu5sEWvSeL9QpmL1pB92
JmK8qKLHuqdN6ru+ORu7hxARpdx/rsLk0iibvxcvtzF69s/6+9MzPQOzeDKHwUu4
UJ1VsVg2rGpbNuke6afHjBuqnExyEM//VvvYcH3L2gfrRSglMS/LpdUtXJeX95zM
42Naz1tfRG52D3gAb15xvQlMtkOR2wadVAIIxWKYGk+85MSkrdFJW3khkLKFPxdI
iaRCJE0Ih2lEjOrss6Z+sbIWZ54rtZC2kUhltWRxVhWOyE/hP7mIdNZPV4AMhw18
mW1KgRjAuyXJvvzJnNWp3VK/j6q4X7c/r5cDyXuN2EYUR9qH2V3T3e96DId1a1ln
XG2tjTXW1dUC/6eUmhBu1BSzYR25AIAjmWOQsHniqCPd++6kNn0cnmutr8v2o+Ay
OjZGfyA+xYFJ8dxmkCzzzoCk1Qf2Byn1Hzz7ErzLlh2zEC08b5CTQCExmdhpksNn
A7aV5+zrCZUmQC3qp8LZD7ix4ojr+mWBAelr7xZxB3BS7YzzFNZ2qtnELpMPe0Iz
WyP8RICP/7QKan+zgysoURwvYuP6m1e5nHzNwRjb45t2TxgTh8769hDJ69IoS/v3
nDsBlpu3QgZCIohKOV7aZHnvjVmKab75Zbnz689h8okWRS5UBkl7QpM/zKee3R4r
m4a4wkyVfh4bXO6xqfo1xj+Xt3jjtHMFumcSS5pPnbDTXzm8gYJVAr/6qD/PpyUZ
UdxGXQZVlddZuR1ke1jWYrZMpGjNAHvD1qcqUnAejUrkOFDezEI1JObOuSaKoTHg
V0Q0lxloVAqNdEeFJFVhoff3XjqyDNN4pirXHE9YpwzXKmcVU/d7Ruj5HaQEwrbQ
MuXH1da6vVdrCIeTfj5R9g7jr1X2zDnXb/dsWdU7/viIzh2ejIbcCHiYyXMEQGaj
k9P8I4wWuJHXu1l+PGUwYxeDp3iCYdIGY+W3F32Wl8e1eUEPr+RgV/Day6t6DgAM
hj4bDvYOVD7GzejPog+65R7dWJ2hp/zpYbkaUJGkiheI5cbtP8uUlxaEVBvdbGB/
GOMFFghRsuttBKjnu6rE2VYa4VkfIstQxWskcdt4T3Mp9XV8KWdLREybvdCicSK6
zP+NNpCYQg59wNupMNikSDKsvQQqtfQybewxYr8XqRO6cEVVDzbG+EljjffZ6q6y
UDu58jBiN810zDTQD3tJvK1O/LxvxqmRzBVsXWvNM0kgJTKso8XBZAIaEMDQikRF
BCZYZAElv9kfzmE1uKCRqauUs8vXxADKS3CDS/18jSNaxRpniw3/Tow0SAoxa+95
sOAz3Tvjk721MrjkQtmSBZF43LtzjHxso8e5lmu+11hFdClk/2kOWE8rxOi3I1VW
VXrtNTCdHeK5uJE8hHVz+eCnYkeqcuhANXNFi2+pHmJnxTMD7ADFBRECkW0RUMyI
gWMsRV9Ecn7c9GV3q+yE+0tjNNeBnG0wRTFnStoqnAHqAZR/ioOlTUKl73U1x5bN
PnwkexLmj63Hz62b2A7c5Yv8lWYg2824QeozTTFBnnTrnrB/igtm7j0hUUtVu986
rgLf/NoCgQVRFTViG3RWFMuH/bIME/QXejWrzT3AK1ugrg1lqq5kHvHXGNC1OB0C
VjgDAJ8lDG8Iqlyuap8SoeoPYXzNwwA7Zfpu/sb46Y5gIbXJCqe1BqJACbm4/mJO
ucBCCOjbuqxg73YBjesH7ehIT9dR8kSEZ/kck/ZN3HWArFxGpSeTO6j2jO9TmqVd
a7/QoK8TVaPrIswU+qeg48mXjNm151nGuPz/wBnMDYwx4SdKIgk2bIwiFvVnQmRP
AJmx15AA2+0ded/00t0Xi/DtiUCvOfjsy7yS9jYgNCHIKlxLrapGMOfX3Ssqk05s
tsPJtyOTjY7tQkpRQYOMLi2W8YP/Bq0aaVLRdYt1HsATMrBAU4WvIg2ovE052xSJ
fdipNylIuv+NM38l7yXIOmg91YdHvffuw7aoB5Ofy2pUvFtQWB6+pWAzdfaSc9qR
zswVQaqubJCjwW1GgIdRz+J6OioNU50/Q0OZgwcqyUD0tipquhQN/V7JRnI5rB1B
JagHMmoQft0IC7gKV4/5md8LkyJ98lhyDs8YZnhUNBUGqnxayFVBv/9uwzlDMZgU
0OLJkgGMyoCsuKCpIOvO+Wisc1Qrw+kT8X96ZtWnancp4T3V2urZiOcAP63U1cso
metnQBzAcI0FleIF5O/yeAamPRKt0lGEkoIzTYTq72Ma9xJTaHBh3+lPd2cjkYot
LpEo2oGu6k4Px3wKEN1a50QVecq0MKMEqoenVdaKSi8UBQf61P9kJOPunkYfaaIk
dQXGIc5q83oe3ov8XVycGK+WzLOBCdj05JXP15vQcOix2cK3kpQZoEiO/jNt6Y3X
NYnkYtG8nDMsxWjJuy9RXDiSIPXJhcdWGUXuYTPvdCNDQXCo23qKSW5Epq7uh8Hs
AYnUpkPm1VXt+h94YjkAEW0G2RUpk53mWDq10rKmN5ZdAfLom/VootjyZhAn8qik
nO99K/COQYAn9ecNQm/W+xNgWNemXN0Xocfn+3jahYHOl2OuXGjq7YnL1xZ24EbK
wQ92EVC0XsJNMMTm68igpMDr/7MGnG7lef05OyzG8QayCb60lzxv4sZmC/0QIH3t
g15Snk4VPR4OBx+/ra6fbhfMZAVXYo4XJPTt/TdJWGG02+dFKi32J9iB1d7mvYXK
toM5g8Gpuy4rKQBRUecvNV61cQVkfUg63i/u5OOKpisBmZQxEhg3Bai6pMpykSC1
2BKNtiJmJZ3/VfwiLRytYLg+DEuXGSYssrIf9bd9P89yJeRBe7Hj4XPJfminAnTw
BDsdTH/l8xNgXI4XzJdZFv/QMHQ9mZ2ddKIo7J0xHYT3svIQHN51gIQlckGgyTQY
jI15x1OCV1lipoew7KtJhrOOOwBA6xGNz2mK0lR3XHlxG+v/bAYSItFRF126LHLW
adq9zBHI2hjb+IST5BqMTXZNNIkCA6EKEVNH/KZnVzEG7rwjNlzlxjjnksm+s4A/
Qn4sxszMNw7W2YbRN8hnU8gNgVGNYQQoG+0fH5DXVdR5vFTNkpF2JPUTTKzsFRWG
hYAXovc/Gm8ignmf5mgbJsxzttcmC4qP3bXCSMTGAeErnuusI2YR3QOui4PkCNKP
DSooDVlCDwAwdcBMweUXYAGxO2zCZDRkUowkUyD5XAQXQFHEted5vkR/s7TL05/O
0KDcvmz6MmagGuko+9WFjOLcJkLYJ+IKNEKsl80u/I+ICreuQ2I0w+dsUY/wBaQY
jfso6oAVVENve5UEzRKgyY1VHEXuAYxFZYzbHNSn9CXpd2zkIwRWELGXDsI0Oq1m
xff9dO2EINg/L5U2oQpaUhEEyWL7LQXcK7HGdn+Avr5/7XwTi/hn1HizdVd6t9n6
CXKMe/AENmQtQg6tnQC2Gb0LQ8o4NfpkjNgvAqIqJAjehCbcBMTyiep8fwhSaCTF
xivjg4k3gYimP1N/35gxg0/3EAGbDOMSr+rbWcE3g9vCyAfoPTCa3ZlE9tuYDQNE
DMX329243TQbZGmYH5GjE4RhlIlnK64OBP/RICSqSXDlTS+Nf6XU31redqXh4mpb
gFcebIIgh4ozgFwYUWUlFnZEZz2kVsXvrQc86CWheiMxcnmQI74WdMYJvhvPEpBk
LUNLnmrXQv6E7Ycsnsk1BSusjBkx3TNbVaULDwlL6Cgf3dKS8+lzpEJZYPalgyZZ
HoSogTnu1HqG4lKe93qYd5WiTaqtovEhUMMQilIrF121CTgu0dkfCA0EFjyPps2j
z4KIkGbBkfyTwj7C60+hzj78gd4syl8+sD2jzXduiXdJs7qrGOdKo22KS2/gQ5jV
bKP3bRC80ShEppporPWe3VJpR73jo2afVqZRiAAAo7KoXhz0A1fXzQ0P80qFxeMP
x+Nuf8sLtbgJL+5UHJI9XUrQqjNrQNSyzbpjmw4vls/5r5r7PO/htsVjEdPcM+tM
HZt+Ebfrao7zBsa3W1V5YkmjJ8LEwG9OtTNJJAKwRE+rJlhpY4MSjW/eCfbxIuYC
tKSf2GlcQczVzTk/CDnr3w3aC4DcOuUKk3HTkUg4hkrMDh+5qlrgFpdvsHXqG660
7M+Z4WupcdeK7wYPqYdlkAC2+01Iqyrtva4wBaTsT/PzG0Rot+UcdzYXqBmUaWr0
N7AhJhM2myi5QeNdZxNrsr6VoyYH20eLPV6xNqa2h4cnB+WF1KsGIscjhqOnXqTX
Rro0r1LGapyZmextO1hx8qBBlsZDevsacG5wzxQgcWQ6iTJ7cwzO95GZ6Tk64CsI
MtfnQxvDvOUs+aXO4XbfMLX5FxqfUCpJusVpL+ex8WFqz64THMk8LjinGCCrdjpv
L5E15dY/EuvduWEfaWA1OuJPk6uhxD2yAHI8Wcr6cKdOV1Af9uIPcUdanvT1WI8k
twnDZleAKJjJnRUbCPtetzvZVR2wNsWCdFrxbcvlrzLCcHIo+Cg7LrOdhXoWE5LR
hEr5bDpEfU99RSlVprQ65pFx0WSG4mS1HG/dFW6JqXmNhMqAP1KbKwLHgpeUmYtC
AqIe9JPiVLrm6A/0fApHXvzpg6pC2dU50B6JKjAoUzhAOhGBmtcfzGbr0UZ1DB7v
Q8XFJjw7DkPL7BPzCbGH6i+S7xizz6fyiH0GJVph1FmrTz3zrE69f7IZj8mnVUiR
4XPVH/19QK2oaeeHWddO+UNNBd+wCNCS7X9M2t5KSWVobjnEBX+oFRNN6S5WofaO
NnjiBx7Cg4FjSgQwlNhNCZmVR2FiKttzcNuweqgoTQawOp1DMjlzah8Q1H0DzT9T
aEzOwu3JI2ws3MRdUdpFecuZCF0us6NVsQq7vgtSrZbkrhzZm6j6N4lK8SR/+nU2
J1FPO1KtDYl1M3pyCPGHYen51DyFK9Hu4uHSibNNfj5Ek+Y5vWw2pbkohkGxVd2M
oGbx6/6ZIj5p2vDCBA5B3lpDgj4FdtiQn2mMn2zcz1CmFnn3Z6eNIPrDtq00/1y9
s+BvGzdojitVJOVgD5jCPoYeMQ3bDck1Ge28kmYlCXlqBrpkP4iQVTDwoKydThGH
pRJ2bkhXCbpUAkWZFZZMGiZiq8CqDTcHVQYS7Ptch/kd1kvxY8EVH2SxYetukmHI
ekK9zHhvjXVhyA2Bcd6D6Gf6IfJbMwGDQOk9/0Ok6VnfiV9GH8OfSjp13Za1e8W/
CHHvDxxFm92UQfa83RC9XAGAEuLXiWNxFbMXFoNe9Cskx4gbaPcJXj6Z4af2OzSr
/AfZdivoMdTGihyLQVByYF0nY4ZMWf+9r4q5eMKcBnqn0qOIaiG6BxMuZYIVvK5o
RtWQ9CL0PMWnI85Crcl263JFOd4efo5IOEa65LfX65o/ORe3nk1e5H2LTMDTpY3q
5SrNLph8wrGSnFImbq1JRyRNC9Tie/aScq6TvwJJxTitHDoaEpuP7mnw/gbQMtL1
fhyQWo8Uq9QBn4B5JTSv2lkyTT49mNedc5QnQgPqr2Ucgkm14DTtkfZrLrtLjfLQ
ZrBjQ696BdxB8fMwOWcI37y5DvJNbTDLCxQGRcvKObxHpgudnbCCXrJNfmtPmbdk
9SPRXUW3qbp2qFuwD/BDJ8kHyxCLjhu/770x3ycbTuzlD+Y79v4IdJhU+jSTLg7b
DwHMfPqVbNSLGnlD6vWfYmcaVMzhcGor71a1C4zA74umGWXIpy6zYm6L9XCeP+1c
lI2thPCmcP2sG6M5HZ3AYWYUnoN1bjzZ8qfjpuZYFTAcNweFIVpXIXsx/xuC3Qig
SvcJSfp4QhZhSTJlRK4+iJFLfZKa+SIUwqcDxBbqfEe6/W8qhQ43y6RrjGs8KRmg
x8iTKtodoEjyeIMkM77N6LnXnzbXNMZd6yteiTHcg+k1rZXygciqMukW+MmAkhbk
8nIDMQycQdZ/e4DpG/zSr8FzVUjsgnLHES+KdWMPwjdlWxhUxnUrUU5eofvtQbv+
CkamN0thuFLaMDDiGdUe+lpWOoN3Rn2AcZQZ9bIoGdeC8eqq79oxTqokk5gmeNDr
8GHrsNEtC+tXIOK19nuI0b2MDCviKFnvbYOzVPMNNOyHR3rvCm3ytmmVKjDws2XJ
Gl40TMzTuAlsqa0yVN6WrIeIlx6pMmH87gTwIpyryVam4IhnS5Zsw65UxxZ2W1aL
Hi0kCMVYuIm8UJ6B0T5iWHxMxVp5f8xZycXOgwTx3UbgJ0XFwGybBLVbbG+u3p3Q
cPzSt1JkclyMerWSlgPVrNH85VA30ImKMMYJpn8Ei2//iGCG92AhmSUBqe7wkNyG
BHWuaU8bQ5WdzBAj0wgBpgMfcs2hkHfbt0OXm6JLNtEEqrftrcrxLahcLbzRDyZy
ajuQQxziXIV+OvQuo9C18oJBx1ZDicQSQgvU9UnhM3QnmZmIn+KVSpFFb6vths3R
z9w8MXJCvTrBRKR2dXWm1aqvyqdYpFepZ8lmrwxNyb4RjEPkdlC6hss7vsvROKfk
2clA0Ar6mKP3bOGtjt7IUl8vy9tUfxZi+b+dOsBdJAEewIUYU2fqr52unaAB+jKR
J3lQSWfdIKCJ2hNDO2Kh7a+maLvg6qL59451czCOLEwbj4ZPZIVyfN7tv82oEOWQ
pdE4NVPQHlCz0KHpB/+6Foh0MPgq148sY9WHmj2W1KR93h+zO0wXiQ3UfUZQjTI2
BSwb5rCaelAohlgqrBJ69dL0jgHeVnLcrGblilama+aIZKnDP3fIMk3Kjw5mvbd/
0MqwgyDey9/vzAdo82fbdwrp8d+S6IgxoxsuyCHUzDBFOITq6bhHVRwm0b76nVv5
qZNwnR5+z5daw35KGVzT7S81bjjUUwjhSLRF68od1RK7ZMlLBlddFnZYe7RrgCLv
5gutFPoRiw3Y0fx60q/b0U+u0CITdNcdVBFUrWH7TZkyL5hmnSwMWzOAs10BKJPd
pKMLnKIMwlLKFIO6/CZTxA82U7ugA3o3qCPP9EpFiXxhywNY5Oy4Bu7XF6j9NT5d
c0phCzBVhq1zawQG+HJFLIndVgKmcFIvqkBZyuKMSAJowAN7NOq/kq4b08fj+FH6
dFawD+KHkxgNfhVy1XBRmsGS8VaQYCsqf2elVr/qX7xsGFBY20VA8wjtfvxscUfL
QMU+XNUbEfrLSUKskW89C+ptjJGvu8s2i7OlFQjBiIcGeNLBQbamnhFcG2cVPBkg
xL/oJshN1nFJjbc3IJlK5IUT4KOLASOG6cT/KEZalvmLXN5AKqGrfxgMsSm67XFQ
J2dHoVG+ZIjhb6v7ByWOBTk3ph1NhaBL/LNIIM8ZmwGiUS1+I/7GLS5Ngc2Shksv
55OYICkqF9Jbm8ervcafAigjIDQqkAiiT10kOGNY0M2fzF9N4UoVk25ZnAlDw+TO
aNNChw/LrnIjHTGmB7l/7FoXh9YMJGQgvHlFkDYKDzboAW+xUi2Y94xQ7pb6buux
e1ak0MEMiOZIIelwhk09DeSJL4GC60gnbfdZZkoj7qvvu4U5HV0vGmpns5s60xtp
UCuA7O/KD+duX976VhtHHojQ4N2NlDqCfeFyOpf1jFFJ2zWg46EfMDa7qgGo/IFk
kFxfN2zE/ZlhPwBFW+kuyDyOIuipaOSJ/ixtWkHyS+HAToL+7I6+ObCgVfCP9L8n
3e9PMZps52mJvLks/PXTmzZU71Tn2TZt/2bEKinDxhVGb3aqhs444W0mM4S8ajhK
WpIm+EIkGvuuj+UwgffKjYY2fPNMagH7Z3CwMzam8s5y3vEkcJbIKjAc9WPWQjcf
NxyxmOX56eFYLm+92wm0WxxO/jNuvTuFK/F7vPkN6w3Keimba2nk3yZSS6y6jidN
ESC2SddRbfiAushigXkEVOGyU2UedYgb3V8SvJL8CA+LVJ2gL1Y7gCESD4rST3tO
AlTmkrmZHJYj0je+QFakvGa6wOMFJ7WraFjJMfzna3NvE5I/i4f6O3PLdZJmNlNk
jyf8+CFG7s3mzE9iW5D4Ds2mE0TPqu7RNNY1kMQrlGHpn0gJNQJ/lWwRZpeTFQrj
GVo71oXiSyKkoJW+dbfxwb9POmuIb4QeERMacHePQUZZIGaJcYBMxBnjFcDZvVYN
CRMgRzhYNglwvcWonyK5zTfXk/fmC/ehnvE7hu81puD02lgBVSeQ9DKUeJ29sSHr
bcNB9Z8xBNfWVQowNxjKf3UV3zi8Sxh2ZNACD1IipWKJwbkre9G7uTDN6RDTQ8J4
KOODSl9fo8naPaibXTrrNbEY5PKO06n52SwVsJ/Q/1hOMB+78/Kw9cIVoMfuP/4/
1kGn+Mdttffr6JbbIV7lRqZ6aUBZI4bn79JQADHwWxCb5kAC34OXGFPF07OOKkZz
styQx2n3YOAPYxEWVlNehHrRKVDV3gft/Y+eBIVFxEcevrToIscY4ZAQnnF6XhoN
yXkSItI+o5uRKuFmJYCJFN4/3fu0GG7Rt1FMk4uV3uxd65ZBvaK0v7VNQvDhHSNN
5kCGrodpBitbxhtLCvqIFP+7Ejf+F6vkG+4w+t1KESTgAoFsqP/vfGQB2JJdRQni
nqoe7/rwkhmC6zDvtfrXQZRCKhYBvI8L3DdOg0bWhElCEMmKNH/dg+sSHA9krHLg
YvwonJrvfifKbrCRVyHBwLJ76uX8nwixnc49PiOYsmpD3+6KxeloZu2gUX6tNY5v
6dqwNmXY+EHuZjxBzcXIKEAoHt3851bCG4oOdEFiteRN1wfIBLFBoQL7H/Lw8+aL
VQEwNbZmRE2Q0Hto08qQsa8g63pHPt4w8NuvWFJONe8Mqr3tyMZ7kEQob2EptTX8
2Z6SoQOAZ1vkslw5lzI97j9+OW9H0GgYA07mFgvDIWLzR+NBIbvoQqZzCcoIZ50p
DDVxYeZ/hE9H0UyVSbltxKovpg36J/IxQvJiZjREID/7aDiPrHjbHou6lau13ueW
3xt0jaj53r503ZUUaWF0LeJANyYxVXWi2PrdMp/57bcv8lkdKujNG0BE6x60gL6b
E5/wg0UxNHvE0N9RMlEwJ52IefjE9uEPEKgXZtC0mLNu2gZzRBIQvv9iwYVQu+7T
nklbvz+M0n0nP+eDiyIuf8u3DOdcqqstv7gKWbsmm7yS9K24JWGn60xgIZhBjRPG
AmNY2CxdymZ/LSON3g1ANQH8/8H7+XEdl1Z9S3CJxAH2/1Q5Z7NQ1NYMcttKCOws
mhGbx5CVmsmSTmKsEEepsG1a7OyHMhqeaHnWrn7QB4cUJ6QvmvqnBniHjDtM1nTc
/LbkN/kCVLIeMgFcOTUK0/C1vQhCHXkg9hNLjv9uxfgtSwxnlS3PaNafELtYjKnj
cIZeklXGrBY8dtdZmiFu4sv7otn6Q3lToMBqiXdsIMR7SL3InXebkjsbGdXUcA6A
zXbeVQePrtd6KQYNUcrE8mld7s3yZG5yisUiT0VP337O9O+6jWTX9enVatVMWqFO
0RxfxzbMmNUBLr0M0ISH7kxjOz5czQbpR+iWXIcJMmZx3DpL81BxXHNt4lw2sVwZ
DzsMj00NibbX5MOK6D+54QMIzK/RHX6Xw8GfVXtydlwmcgW8DrBfN3o5AWWhK9J6
AhBx0Q5TxTC5/pGlrX/A6U/KbEA9r3MVQNCoCK6VvckEGzuSuFJeqTmFhDVqv85S
peCUhJtLJmbvIB79VTszoNJW672RhXkEF0WsAgxphXw+jo3c+ywbsBH6HJfMU1WI
u4ttkVktL5a2ZERWS85TGSlxCJxy6yxXIKzuuOE12ToUXxmOtiZFos81TI732HVV
3z3XWb6+wbKiOTeYw9KMtFxWyN2Er0kKJlk46nG/ELWPvLokGI6Kr6ZvwaaYds5K
mfLtWQl5ukF210+tRYNpyuMS4+Orca3RFXQPtpSKAhYkk74ARkQXG+TGD78fa0XR
2YLo8NvOZJB56Kjk5ygFfsz78rsslMIw2bBuPm2EYeOY2cEH3SFa3T3aHZHRfDtL
v/HaSUVSIZbOb6lvIJxcyPO2wu0XsQeAwxSaTt42GnwTlrgYhncdKcG02KWod/pf
E3MK0BihAkZFyJJEHYupWRxN1aCqmYF2IkU9BlTG+fyHyyPxztbe39GOeGCESL8h
okuqewGJpdMOOWrMohs5g0ip1/+jOooYyvQLkNhGFDJ+ELcY7isk3kbOfOwcmVya
D7jYXFgPCTZwcK8gNw5sFny+6PmOCw7zvLYtSy6fbt79b3vDnlPpH07Wbm5LTII0
knh2Mx2warQQz28PuvVHvbYdkULY+1y2H7B5qhbNTAn2gkSsyoeoF/QZbTgC3+RI
5MO0umcPwF6XhMB0M5cAkCkeVo0aZR0LqHJ0yHMzdqPgAj7xMxIgjzqe9grP6Ypm
OrkEE30Leb38PLr+1zj5extab7+ir8FpDMN2odI0PgQhli9mXQGqv1z7NNYv8eSj
Ikoe/7BYOjvm17ynD7netGOhcVwaFxbdYGfbG57aCXBvZCbY5hW2tp/6MkmobNKI
yYOpFmr/ZxB8wjGSTqRlAri2addWZSp/PGQonEMQd0yCfIFnNfvUc+FN7DDLcUDJ
3ke3dXkHL5up/7xJSAzlxvs7Zl5LEk7qwVyOFQzYjIrsYH18I5JmLscYTniSnqXj
j+yzgaDoSCS1PUp/g3K8FO36n93UFzzfzlYHP0HOMUxRM0PWbrJhwYwUmdXWfIru
6q8XTGp0qByBPQWSg6XbDd8wC+m63UWn8DmrKITELQ2pUH2QUO0gdA/lvj3J1oIU
bTi7TnBoyUI/05OqTb0Ps7QKvxYupvbJQzQ6n30FXAqhKtJW35og19MKJ8iEOrDO
RcMvvWIDPGiQr/4OwXJKmcuONzq+sdgzuJBrmCVfDRsIdfXgWdEmP1c48mX5yMje
o3AonO5fmgPIkdjffBHDpRs6SpjsxUG8N8fzpNBW4kYrqJXaCG7zJ8/NtD6V9qa5
+S+Q42PDgi8RL4GZeLZT4HCLM6CVK0f4nvIK3LHSbpQK4GwIiHa1Acv3hPLKgXv2
qmuJA23C+0aNytorAliZMPQrnDfGTv1QnEGmDbsYIagwY2tKpRfSlz4bYZmJ9Wbd
kEDoNkg1YFA5WS0nSTSxo4CiwAnrbnpwR4+sZQYvS7JsTHGQnG0fEUWhtv3D3QyJ
m6+pD5B6T+t3/Pifs+XPveCdGThIfUWj0sqOvh5vuVjDMsoFkhRotNFvJmi8sVzP
nLJGfZOsDVIvvdNrVRGU6hxgf9HU1oP4XjkF5LUCT5eCo0rr/tHIfSaibW5e2PV+
TlJo2H2Z+eD53i6GyoFW6gB2Hn91HZIiTTAID6ZgFmGp87SVQ4em7PeBAoyeCQGs
bpcA5j0cyvu2f7gAWcOTEDJf1qmxHHXYCkmwk5wXi9PMhuMdEJz9hN0EKANa6++h
Dwuz7nrbCFNoMnugrT2Vel5pu7Dok62hzbbUSJbtBpeuc+t63QCHZAMVYBtQptJ0
66ffQLzdMn6g9pIjlPliqwoCK26ogFLwNDEbfJk33L35FSDKAxuoJE/ps3EzbsgH
tH3kjo/jc5dnEPz0kaidnk5JDHzQVpuZpWAvlv7/FbT5sCK14yg5cMjHVWgDz9Dk
ktzGifysTLjWQqs9mp2SJdQGWu7YikQSLNrC9xfQkKqZRIkCYlgmtZ1f+s4s/RTs
VI7WxbQ2z4DQXZaezChRZpIPr4ohJPDBkIfAuX5xsWJRztY7J4XuCf2nVdyQHSuK
L0vYCb62z5n58Q37S/KVsJVEjhqOQLX3I3lmBmZpkA5BkUiUYJONBV+6XL0EdJuh
ilNEgI4PKQtyHV++FcYT5yOmMX7gnPrmlVXLlzIxjnakPK9HgKzbbIXk72e6L66H
k+yioaecQV0mTsTD2OIPyOxvCacdGO5omlYVse5IiGkIQrkDjqCLxZhfqZCPRQKm
aUONvZos2EpRzHa9WjvNhUVsJ1g+shqbSE3cgEFwP61zfNXnHgnYlMrpsE0ytqmX
lAW/fsQQ2cHnpce3ZxQMNZyne4z/sUkO1swTkj6e0dxgbN1v+t+EPNeQR3IaYHt5
DQah254VO+HjmeO0VGED1e/Vzqv6r8Fke1Ayyv9zmyz4t+Ob7fwArA/7uB32tinD
ToLdyF/vPOS06QlOXNXfT71oZpTdBTNOGTYYMMdXg9Kif7P/T31RCrSbyCA4rs3g
DSBHr8+0IsCLaiQnl80EMiHhBVPuAIpq8trNxHSforLMTTn1ABzx5MYAD4J2Oo5n
Cl/1uDp32FOD9Ju1mQy/xWkgw86XJCq/ZzJxGDYbhHUcS1lpfKcHyVaFcJ29Qyi+
JcqXnvykAkHbJcoTTb3QrlJd9H40LdT0tmbKfyqz3WzfaxlwNZjhzlVgd4QhOVB0
n+tBUqvUhX0Qjcyk4QG9eS/cFz/K/kfn9vSDV5k5WXbar1Ned5BD1Li6Riy4I78/
9OGy3ajtF+bf+PVAuLLzrBpZW5BR7ngG2rZvcbv1ppTcEqWcILoAa2hPNosly4ks
uJW44xaZ6V/ef9x1pP34bqrapZviyrSmq7GhHzZILLkh52yQ6aDfk1It2TINye8q
NKO5vvU1xbCSTh4mPjKtuKqZYLMnWWGh49dCqUtOQ2JMFIiUSpWon/Gl8s6tuQon
ht9m4BuJ4xCnD4buDKGraxhOJ0Dc3cxk3HkzrVic6rrTyeVFZxNZoTGiM8t8I+BV
lwpg4ur6iYEYfiD43B6D8jk/OXtf7VGJWUGZf3Ln9FZljTALkUkv38A2lapsWjsy
hzBEpVN6F19fgue+Aa2z4gI50PmRGcv4pIuKB/CyTTIZVTnLuczV49ZqRsLJKQ2h
0YcvnhLufZWFBxMGVulNFkBM4M2zpJYji7YgrNX6N4qaYPEKAi6F1IJ42kpFpXvD
BTSfUPFuAebY3YgzrO3lboc4Q9XRER7sTKEZEDcTXZlZOSB8sn9uv41Pb/LIsmm8
ioFiJnKL6D/Smpje1KHL1ITT2wOeq6DeC3VJvW0XXc8xMsjmqsZ3C2V4XF3CSFRY
jMTY+zBbeSrGDhuwW3HqsqttENmbkFF5ypS22dSfIxdDftMFIUR5LKdZ5k4EnaxE
nLSDyZW/yHc1mM/rfVj6WesJcVXATCBjdL8YE/ZWzY8MEuWQ64TdxnkWTkhfWKxb
q3ikJ18IQBlT5Oc4zZutIPJUZlcwTbqmrVwPg5Zo1l4aO/d6dp1adiXUaK69nTRO
iu/PSWHDWs/PcjRnzCNdrGaIPk/mwK0yfMNCvNPRGo0255Qtir19V69rHt6X3yW1
QjbNnQsSC++qdztSI6WqA00TctQyvyoOqh2wQMa337b6WaEQSaKDyXVp9ziXf6vf
zCQUsNxyWrvhiEHMcSl9vtYypBNrq/I4rzxbfo2NmGnEotBIyVi6mNxctsYOvnD+
RMELkMASQPF/uN/L/BKHYRv25KcueljMiY5dDMKma4enE4XzNPD8I3v0GPuOshSM
KS9VmioZCIJvLGT8gJ+cbtIXGSL5ATRXWYCsAt1jNEqzPNwr/w0KUZAQ7Pz7euZc
o5g/v/Vn0P2H4r1OgPpUA+z/zH428Pa90BNzM0TCFWlngI+8MMhelScb126zPT2X
BYxnrVl1aEBJyUAB/uq0lAczJl6SMywth9kNcLR9cJ2McFfO25riRHjUrvDtdd8i
EzvGsKz+sXeJ0TnG5AdJdm98moyHGfl1Zfdq+4O1CDknnKVA/KkBp3UgJN2Q9g0K
ZaMcjTYZxcrjG+kK/lxz5yCiysUyu3tcXu/leswqw+gdfB2/etRvvU44me1GrBJ7
UQUoftDg0vZPTQmDmSTbBdYo86jra5ypYb6+yIAcvoVyvpu6NbsFSdXS0JPO34wg
6pX7+QtWdqckfk/734Ys7WUIyRMnsNDR9r6Yhe9vG2KaDMPl9oqcua078+HyoCno
9V4/SR/RgFY9Bg/9c7xe6MGlpQvyPOjGKPK9zsmg1Cv/NVawvXBTEaadJtpMUPwo
5C2vMc6TDVubhArnx1suOqlfpmf9tynaRejEr5F+ft7jl9lfLapWDbb+DYCULKgB
o5W4zXZ5NxADbuy4oAzJ2wMIPTPPhQB5+pxo7AZyWSPnLhZXZn+3brpV5wzxCHTA
2UBhshbIKOo+R+bFpnLeGRIRRY6LxHhOOCMrVAv/c06mKCNQDKeKO/5CNynqltJ5
lYU6KQd+yLr6gmfi71jE04Pv4Jk1Hvs65ltCisCPXx63uwBCAzL5/5jeMAQM9KXH
UXeu8nHVedIOJCPgJCTtV5wA5JjwM+zQ2CNrnbBgHtzf4lhmtAaklJt1Jd91iRXu
dIH6xGA4nM1MPBvo5yngCuGa/XAdpHdeHLy/x4BrNGRNkRfbmOyBSRrlww6zlGFl
sAmsu60CK+S8y1VI5NhBN78NVycYA/n4FHkxuk1gTGSVk3TDUW5ZaoTTf11FcajD
MGABrS23JGm57XnNP59nwsAHJf1KQbPD9V0u0KAzGeEZwlk9l7NONCqPbWx5g8rB
Bx5nLj0lJAM7WGpt1bF/xrWiUL9IY04MtzKATc7z39JkTA24ShOcYjOMtko0C/aX
7wCEqJe+Mw/UeXXga/FRyKzLjk5TIR3K4YSg4ZJ+JcP5JO9CXzhgD5dChSqxvLHD
FLto+VMCHd54AnR0Qcr1IvMK2vQyGxUZeOVToOwJ79vUhs2M5qkLSV4RM1zm3P0z
W8ylg8EnHy2CSu5Pon4vIO0KXdePA7Tjm7AQagVo6bHfnkBwwzb6PXLm8aUIKJS0
7aQ3WHOUyzzu3KoPSQFGm40hExSyvXREO4MH2DUsxwhSQe6fmV9xLs44qMgM7ezz
hh+kUVSpxQ9+TCxnJBzR9MvEroD7xntRP6Ik73sa6sQ8jcYLpC1RoOEWeDiqXwJn
EgmpM1euoIqmYgf+JYhL+XwOexVW41uTmjCRnNEy9S6iNE6eBir1YxGStLH7+Yld
isFsnkHKglIbU8yZW7KYzojRVGfRSsr1jfcsJ0btNgH9OGQwNVRLFhYmgQ4o0IIS
cXmatZNhSrJwL890ISmv3DXrZxCSgNffF0wzxFgeCHb4a8Pm67NWxMrPaXLiD7NR
fb19m8byyLUTLRkq8bSL5h+3qxovR4o/dMqv8zPT3/XBLbeoeAuVX2qmjxkAacmL
ofTNwJ523jSM0jVHkJJ8ggpYHI206vpyXdNYqDz00F5PpkUfxyamXp6U0c8yT4Fy
qiv+PmipXGabpnXDLdYOfBFPmTWh2HkvfLly1wj9dJGEsO0QVDhhFA+kIm5qf7K5
wi8NHbT0CyFsCmVeY63d/190ejytU68AKk1w1Zqv7JPLVMfPPahA21cZ/Q+aUfwM
MIMTFWcr9szD72a+XNADaW7TbGas9hXvm+AeaLg4hRVoBQLgjokoThZKl/xkJw83
AHFT0f3lbNk2uPQkToisuuBT4Od4UKqTKKkjVkCjvYHO/n1JMau9F61RE9Y5M4u3
DMlZSsCC0CIIc07a+jTHq9VX6tk01Rp0crUtcdRCH+ucAq7wYxXCguNOXr/gRcxF
uG655H9sKlLK3m2rE1xw7zop/hRG0MYRWKs9sF3tUBEjeyJWpyL0CZJYzoDtKFHB
lHXrzulXNX7b6u7NLQMsCCx0Afj07sbEk0LlyxjTDyPuC8jdNdknRcWQDCYyIqZ+
qyiggUBJ3pEjZAKKHWEo8O37w/TodHlyL5rhUvbembK5T0AfGTHGcIqwRv+43OIy
Bwar6yVDdM6eOSUE8518feqP6/8SixK4SKq6IjJ0Sf7ryEuXseAovccPB6DMYor2
oA4eCVfLw8Zo7GLMHmZl0MT+zmzESAwLtSn/yopPojYrktrcbGRnjRp3u4Os3jEr
mxFKpzvFAshRHO8jhhT7PScechq/eUDLbIbfz15vMvNmj7nhbfmpzGOxLAFwAAQS
pTcvyVWFHrFHJE7CHxL9MvqYqpS1DOp6VFdsGncud2Aa+wTyyp/kwICgIetDLeaT
ELuE7yY4tfiWRmcimt0zYNUbxAIZ576++GTcktInokprYP2ZAqZAOst2FDu+N+aR
JpXVzMOMUbxqNT3D/4DmuJgNcBE8q02Z1amrcKh7hUx97rXYT6N2xykMTrip3E8l
F5ykoOGsbMRB1efJ84VsxF5dh7NNu5/8Je7xRoaxt7aeIBHb9254aVYssQJ7ssCP
KySjguo+CDw2Bo/61jxiSNzT/1d4e3LZh5kZkSBbD0Z6v83PHZgJ4+KQJt7sQvs9
Id81IkNWu1QZcjDwbPPZRSuOT56IreGhTVl6t216u3w4hXiEGqzvqCRQ0bXXFRt7
Cy9FUoQOUO50Am4eIEHVPVgf1RpNX79yxmgAJ3siCHKngK4zG/SIBoa5bqogKYXY
wTajdWjTK3KPzRMy8/9CKnNdN3A7VNmt71aPiE5FV6Zk0uuZVSuGnM2Ar7T0L13c
r7PJ4Dlcuy5hkVSok3c4Fcwpj8UlEnXYM5SWpvh2ykyrT/2FgyD5KE0UXWYVOev0
HgJP2GOMy0o3WOeLkD0pFqcbdWdPvgVYo4V3E9CmTfcTyg6v82N3VH0AGhEnT+Hx
OMHk89ga5STrQ7VhGbAbhRHJ01aF9bWfZW6R5iGDiHPhmYIkcqA9ds6vEwtO2cpq
lMom2XylOiouSSp7Nxs2+/ajhgM7WUnm5Dt7W0OMIEw4n+m3JWtPKb/66CyGYU2K
7ytkBywDj8DMTFOK1X1F1at9hoJnqXhFfdpIsvfeQF2jwMtIHsSAWxw/y0RY/CQI
g8jMUf6tcvaVuDiayn5Pz5G+9M50cOAUyRzT3p6Nz4EFs0rb9g1+bWz6SmrNXhDq
shLn5NS3n/Z2cEUTnxv70jGuwsYx27AIj/K2dbj5emaN46dNT+QtEc3qKVb4CQHM
BouXc7TFpwfjimZLtvewTbrcdhwLYtmqaXjepFqNaGFX6MwB5lxhGI85UyHccLp0
nT5sZQzGnnXcODX2Ngs25sLfljp9y/pwJPX9pmjGCMYcV9ftSAOjG6FMyfpGfUeW
AaTznrcdJRwYrVVkNZSnXli4g97iOKJHg6a7d+KbEOiVsnztNvi+AvaRVZKENJjb
EUMmvzVOvgagisWRtlKCbp0OnusaPQvm4iShcZWfajoSpv9+eBDQRzzMJ6Nz1Bnw
PYn8Dr2MzwmwDNj9iZwWj0XjeIvBmWD4f+6XtmMuOHD92XBjStrgT4jXuxBrRpld
u8DQdZ85Wz/p0eGqu7JyoywGfQltZfXwibwbeTD3+Ua5J+iBMwJ3PZ2UpNATKXcX
WiEeWzWcjjqmT9A9Y/BAkpZvRClx1cQG40f6YZBwig1Rm4tqmohCtHMQlg0UBRbj
KJvZii93CC8trTDIzRjA1dTe82LnOjIeeogksiiokCONGv+IJSkh3TdZ92jS0bAm
++E9mkgRhxw6tCt9WhNM7gBF9exVvPejWjl9ywsDyFdQ1P3ui+m1+xMKan8BueV4
Bn+hM8jrDMvu8VGA00B5o4klzPfEccw+Lmi2QLNxYiVK7NX95OZHRUmEGMF03JwG
DkPZNCQIqNU91bQePpcY6u5AfrIwvQ0DdyICTux2+jWyGYeak4Zvv857iVR7FV1U
On/uxSfxOfqQseThqk6w7iEToBRAy6494uvnOJPb7XBWS73zquOhZvts1OF4kW6w
VqoMfdFAr37HVoxKAlxTDas1fg3RMZkr+wpmJv4BsciCBKnZj1cqlfzUoZg5jUa6
fljFenQJUbbIyfVpOLzbvLQhR6HXzKOfQshzUcDkEei5zBFjT4YuPspwqqcpTiSY
Ig3Xz6u9KHp5mlYWzsxypKLVc8a+8YcdNtO/1pizJjazrYJpnylI9nVQOjeJvGKy
9ULj7iGgaupKDAuhfWoPBrmjXEwkmLSDd7lV2KXLyazsnzm0Ju0miwymCX4Ry0LV
PfZJG8r5VfNH3bQxqkUJ7g2hrydmmfxBA2Cg7Nid2JngUWH3txM+NuBFk0V0YPWE
tS6MsY2XTX0rT/nj7zCnV9iupBmzwiIwn4xRkJOqOf7bksw1hlmwgHkgqK/dsiS0
+Uce/cEzjDO80ggrzIwtZV0mE/idQdFc08+AMZzmCW1V7E2BWiGw+cYUbNsHnQ5t
IqNcolh964w7kcqonPXwENj0Q14P/ySSy4dCmdDyYuQrtpnD2sQia6uvGBJUFdLf
7MMI+YwS4ggIHNohTZryz2U/tP/miXfI9tOcapru6YfLPrWVLcMEiydkXT9C1SCe
azjlB2qt6QKH1OeEA/qA/W6aH+c/Uzdmss1TyEBcHEBQYD7jAGQ1YrFAT2Sw7DgB
vmFjN6OYYFy1CRQt1fKA62X2Oa9udGi8KlbMtzBuLFTCu93zlFDRmKDuMA4qHPhk
so5MCo+wk81phzOqomFyRIdbskg07i1fVRia9b6Cz6f+Dx+ynUxJGfMaecfPvFHt
hXJU1gpS85GJNZcg7zvhymhASyZ7gYDeQbjqEIWJsaBp9cUlQW89M+yfDztwWF+p
I0N75j5UHnaEiPUO7I1WrF6HWMBYyze/Rlu1uZqfXLD6lAXqhyBZA92ChaMcK2n+
wzwu9aj/fOQtBTD2Tz5vFeQC1cp8P9wWpXOSe/zSM4wTCd9YfuPExENd7oLiu5fD
y+qQA6yUbKNT3zChZqW1L8jFUSXhHY55tiWt+EsnkWL8LvR1BD2W0UmVUPBLCslJ
JKC3+jcWriLRORBpMOg5PtVYHBmcZfq/lATch6kd24aqk/Eg4UU/+uxU8pxgf52M
0p1ftrXDRu5Q/byu/pCcPpmN/rZB8ukgIa3uZ5MpZaJC6fZ6Hkgz9/EprRSa0wgP
WWX9l4mvtCAfitImvLXC55HW9BDKxcAPFkt4r5EXFubUS2zjtywiNCsso6FOm1+b
kahbWR4OO+8TJ78LQZOoTlbbpB17Rq7dYTIeRJF0nE/QB7y7VfScK8Mt5Ym7n91a
SCgLnBzQgS5uq4mErrxMy+o56ZxdefyAl/vf2Po2jad+zDa0Py5tkNIFbhFWFhWx
x9438M2yLkZiiAmqVd/6T2wYcoucR7JH2eUn5sCSmaAMQX6GrSsNxCGuKZBUIoom
61wXbIEkd2MYDIu6QTA5xdrtSdZwEf/0dwpEW7wRT6de8LflrltsFhdI9ukT381+
IlRf38Nb5xk8ZltC8cRRTzO+4j36X/GE+pe4b3Rme4fq2tDkHCcxDqiLcFvT1IRs
kG3M+D54f3Tvzlp/unQY/1ZXJGBE18cfgPKAKx/EwkqZysjwuKy+yADqhme2S1Nm
MOvD0u9SL35YQj8lWcw/lrKvPjgggtO0DOEwRo+Ac+x4Zg5j4uql7vGaCznCdEdG
qn5eQbFvDokhSAMs3Eb4xf41zecANt5r5s378ZhmO/u7/cj9dbTEE8S5yaxLICrW
kINiWFj4JyouQsES7lH9vAxqxSFkZmHlxMfaRHa0KICykMtWk0nQjnh6g7LrcHmC
3w+XzmSmY3b8XHYSn9G8Pv1MHHVGXTAIKJ65DzlFKoHPkBzBMIbkGGy3lcAQgCBa
AGrB+MkQh0nTHhXys+m5hLVW1y6Rc2LZL1V+Mhvho6Pndu9CnGbItEYRZl9uxUMy
JLNx8pigeGcsHcJijsm4MehLAFrkl4/Sd67FtsF94CRrV4y1nLDBCyaWeDJvIj0y
es/xcWoXC26Mqc/VZj20sqPDnVCvBH9XvzY1VPEwuQmYUBsEdzKkkOwMoS/Rcp2b
1uy8RqVTcpfHTIrJDEKFbv7FUeCZH8jH5KXmrnWfPjljl7r5w6T5ll1CjTeYvL2z
xjeBYa5eHMPeS+Y3RkkF5NMdAhkkqbEl9hCW6v3X3TEzxRrMn3LJHU+b+Dv5k078
vIziqjibkyADVhQWqocoO4biJIk5r3aJJuB67mZfq8PT9XcDTR8EaSqewRQZjlAD
U+0dzoo1KpZVOxgQxOBAWVweQESu1Fi0eeiZ4X3NQE6C38Q1r/rbBYJrahoxH3fk
8M02+VSny7rVwudUKZZDDVtLUueYiT8p/c7RePvE77+BWjLJXzaqLmo2gm9BxIPa
x5YFDa0uwA45sStyY01bx30r21mqJrdhswc2LSLZbI+fkrHzn25d5XjTWTj1Zwd/
G+tD9DLmL4Yj60NCOrZCxFTUm0GyuTAb+dvLOSj3cEccSQnGaxGyoq9ruoLjHTXt
hutFIqb9cd+a7S+2PAOMaFcgC4hrsiG/PYTHEPGmqp/vd2U8hRkF4FFtD8w6DN03
0Kw9s7TKp4aMqEDE84Q91K4VCoGA7rbhvkmwgQrjiPeF+KYT6B8Y7SMJxZNQmYJi
tm8LzW++gylXetJPJnBbhixBzrZkk+AXLiJW74cy+8D+yQziWEUR3ukv6QPXihxA
0hdvnWmplXJrptQtyXSZXwpH4n9rEqZjVa8G4p5UIf3uo3Q/NFsyvAn6McbM7Hf6
rrq/lEKe9zzEdQrz5UdnnzYErIyI7XbUCVweuvD7YZDFOxfA7ZzbdBLyYFypjcj0
MQbwkfUugB/+WJEyRhEyZ4WUDUfDZmQ+5v+x7MRJ/ay2oMRbr/NEyfxGERCfngAI
ubNyagj3MHODZSSYXQEHDFqveVl9GScu/XVOH8gZ2E1IWJYLVbzCKWVQPw7lHPs9
3dVEwY8dwlU5GLmYCueW42INa284Hj6w7O9TTfMAa6A8QDbYJaxqF48QiRPf7r47
RDQlYQABURol6eANtGqGMXSXCyP4ecYrvDS7E7MGsWHxHgyzii3ioNbEF5KKfHpb
2GN3hgnBgyR36VidaMOY9NrpwCwSrJ9zgQeygyVo+V5vnC/V7GgpVTbKeFyKHgjN
mbIIEcbX6Jw1w1mMzArMHFfnDc02TGwEy9C4Lb9sh6YZG2BxHLW8uQ4OKRvA1L9e
16813n7zgFKMiBW1FUxmzarBmyd9gCWy9rorlMJd/t2h9OxXJY/3K3V0YwWEjYE5
G/LAWu2upaDYcjotYpm1FaCODasJOD2w+J5Q3tSF85j5XEtBo9D/PkaL0+rj8/0J
BhyX9aEM4YR6eSnWYYQnT+rPcksY3+fAnCEpB/W/njqNJD36JlFKAYo/z0JCJqqa
Xh7Zv3zEHpzyzj3qGS/nVWfDn6hONiW0yB4s6sTViMC6g8M/LZz9zSmote2UZDrx
efl7Oz4MkPvikZfTX9aQ9yHTqxN0B9/HwdTIeldOsnEdVOGJ7CLnBX3aDNTfTQJ2
dL4ckzRKwFD4dZ43H6r+fOnbhkorqVp2ZWobmxyuDZQXbZlPr1laIBScAd6j8udC
JQZAIExS8S8OEiFlHi3e9IjUVEnLNMVSkNhYK15wKDbX1qe8syOsDLam30EZ+s1p
FEL5H++4c+l38jAA9KxhdwlOyN5wbGX9QFaTnjPL+uIkylMX9twQi2WsZzR4ZWnc
PN/C9WsKKNiXPx4tLW7KiZS1zixvFFkl8k2RCW/J62vHGGnmi1/OTDVAVlzOrpcv
B31IXT+SnEArl5wNtb/zooAq+07P19k1lE2LBr3m8m3ExEOr4Fqp/ZbtA0jth46Z
aK3YehQD9hbf7rrOCBH0AV6F6P176J2okerTQdf+jsRD7NcgUFQng/l3KhQlUPcC
oByAL9fSCKU2CmRQzkJrFwWlRsF+s5bfw2wCL+bL1/QzXj6y6SPodOV/ibfenvEW
ChJcXpo4yKSd1X3IW/XueHflyUXfELplrU5MatsPv7kRxDbDjbW/qgONAqM9tye5
YjpcMHY78y3O2EBhn5SqvxRZuLLymj5ucHcjBdBUQfyXyCeH1noC/lHc3u7DfqyY
4a+6Ii3IJD1CEmPcNPwsrIMvydmR9n/45G+QNBcj2PVHwxpM4T5hPYdx22ftytsF
Ahuwtrw3+HfKIgwZqJeXIs4MG5o7Hac4K/P861hvvBvYxGpkqWptbP6e3OYFhofC
13UGnBpH5+/iKvgTdriVTSZc74WJivF6Ow4R8FBYZqsMQpZWDkEgZ8isdy1HlL8P
Q4QA8pVwF6mFBRf2lfdMyke51KIfRoctULqN8hk6FY4rxetohF2DsTcEAyUQda+0
YVRa0g+0XLWzBinsRcj5u0qmNfoHi5V+Y8FEangaeGawGouNXZypEOk532Zb8SDe
x23FiYZsaVZs8I7IXg8fWt++ECZwk2VNNlDiisq3zWCrXaNn9Y/KvO9igsTEF+AS
XgSO/dK3nHIVDy171MSDKBnkWEPVGBGQ5wMp94Bq7jVQfXL8lbiI3ggFkZYMOBo0
Xp5tAanvbRhYZeftqVgYZDPxHJ3xE0CHzcsMfIq8NawWiEsfW/v4ohnqhz6795Vp
mpEs0HjbiFBj82S3usSG9Evnp8Mu9jyH8oZSkgdKB5qvqi8tyJpZh0hr+4uY5Lf0
TG0EzhITTteNS9d6JOgJOm6JmdxRWSLkpQOFYnM8J73ZYs7bttXB8GAFvSsFcRHh
EuB+GTUVnu3RW4KXA+bQriZF0RMJ9s5ILeMFQjeB18+FHO7bMbSIZTiIgETDnXF0
K4Osh8ZBfyl1CSl4cgWftpS7d5Xs4BH4BASQA36mQd1crnUW0C2AOrQAfq6DZGSG
WfuJQDjsYYjZRH9I6HBKQbBHeZJ9V8g/R5N1Kpuv9UL9UOnB1d6YFyd9RfirmaZQ
qmfsjBjidPc3XFkQyhi+0m3hvdOYasQvXbG8hYAbwfI0uWTC/HxmS+2jx+/n4fa5
pugRdPuzCQUEGK677oQuv/UHlG+QG0vdnOyycEvbQXq+Fdd0vwrqH5VySmBJBiBl
b0+OBe/vQxf0GNZsJr1megdgQaDm7sS89/FIAUAShFBUmBVrJM9LrL98GMY7AbY2
lGgenqoVYWwAIpbCtphrcXPDI3S38clfAb74HGHQw/dGrZU9ZUAMq64Lqw20nUQN
rV3QpMwfhmmk/7T5VimovGxKvMuFTgPSqQ+zU7jTh8MS3haYVbTGnHStyoBv6MnI
QOV4WMq8Y+FqFzXNQLzGnLVFSXzKRsDBe/smnenZ3+DeQhQ/u0hqT5v1yNMYCIiq
AIpUU1WSJ3SkA42jr4tYevZpZqqDKLTVTp62dVfm88yvDnoAsV+ql4Lt1nzi0oB+
kB1Ez2k3TObCYhv8nSTSFNr8+Sw3LHJWifVrluyGq5R9vddxpIAAOgZFi2rvG/dg
S6wTsYYytu3NYgttmPM0yJDRy7RuNKs5NxtL2vzOblUj7FFBsOynlqCVJeitrGFf
uHimvNpC5nMvpwW77bPCe7BndkzwFS6Sq6wFwcZTlK3gsKT2fZ5Mh/XPnTtiBZQL
1fx/HkG7AF20nD09cF1OD4c4JWfwk3k1T0gmm2DEPVrTRPrLHQ9bRtG68MBM6bzV
Ztp/o8LviF36goDMkb2YntHAsEAOBcwRjsVUK9AU3QKuHOhUwd6Ayjhj/mTxfjhj
4KVu59OlsmAoUrxnakEhv8oZtC3IyIdm6GHbdxs4hLypSVHtrY4kY0/Rov/7F8fs
xkEgTUM/A5Ul+c97zkKjyvlA/xJK2OomewmQX3bvuZfU8/eyENXbkRJ69KdFnCMi
rSFchkpzVeNOgBmVXMHgD6L4h+kScUUjjpkuz7beoPcU6Mwc6lNemEz/ImhX7lUQ
LuUjFS9WsYUWVFPlxwBjsOBCFpMSH5SqXMcZhmsNOm3LS0tvmLH38nZlijDOaWHV
uqMb8eVEy7PkCA9fZ4+w0Rf6ZrlZlZhlvLtffcXjuYB1rHTb1xy/k1zyKzgXg84/
h9W9FgZ4ZzbHguQbLjymt7dFACzWEb0eNs8UpJE/nsTyrcI++fp0Yi+pFOhDgC4g
UunPcl9vZk9cEpyaVt/QtZxX890kqk4FLdQRik8lqyJSXgQLhLi9kaVwCA9djS83
R02y12YOa8gBPBddmzQfmY3DaBrjAdgSmX2XS50GLgjR1nd4oZq777EENhoXW/dh
Rs+HTsf+VEgYm416Wizk6NCmltEWIj5fhByPV6uO3qBzUMFSlkc+iaHmXO0tW7H6
b4+R9+AH2MsJvzG4HibxyKL/x7EtB72UuzNnY6pKU9SGRn4/EWajT/iOMJUrEHhZ
uITHy2c9AcOkr9E5/oMAnhg2VRcpo/I8KwUd2jOYuTY1ftXtcSUEJzO0UyM0LrHE
UW2U5bFOIPw36rD4KPQm9XmbKOICHReseY7ARRteXW4nzpQ1vpTu3jHchPxEsK5L
0d68yzzUS3f7M4osSo2nCJB+jhaKenH2NiNtq+C3JgVACRC4M6zxk9Lhq+vSRLfC
3ipnQHdRfJMYJUHY6W9TBydczvQZEoyfu+0S/80uFVnqWESb5UdW89umgUutB3mJ
U+C7T6iaGQgTLawX9lrVBECbvCkPfmyTEzT5AgV776fWljWeTpQgaf1DBcEQX9VT
0gytGcDMseQQ6nL4uBEpfc7FUl0+VV2UbQqZXve9kSn8QHcle24pR98PfDD+ocD9
jgKutw7HcSVmu0UtXZNx9ZZ++/qgTljzkXqvCcE4shmScsj/XyWeVm45H5l+svYV
y+bPyjW2Y29fRkjP+3VT00+V+tAebkK8CQOr8zOEzIIdhi5IJIL1aFHinocWHO8h
bDSDcJxWXO1WYKeT6Ju7/jlchO9iucGMvc3z0Cew1shWwpjmzXYgPp8BdxWjwHbu
6FPpUrumr/I/M0JRHk4n9xS0mn+4HzrIJQfLQA9MUthIGdsN+kJyoOFePHm1d3s+
GD95NUn7GTEbVN7ZBeB42I6sKX5Dl/wWuRV52BznXkeBUdxXuty9S+ixH9+blFhp
QMKTntYH7hdmFRgZd71Xey2+51GysuSvxV7B8ZcRolF1hHGzBrDAidb8yOvMEmDD
ZGy4rHETfRVW1k7hTtbRUPagkaxERIL+Q64m12iebeVzGYsiuR7+hhSoN3C2g5tn
RTobLHPjr1/mq4fuAlBM/7zCJo6hFd8bcgeeU7IaHjcfBRqoN2Y727d41BHl0d/9
+Pi0r61WaZnujWgAVhsU8HpzWeMNLRr002WEDfZI3cnHUubTGBYnsrVUfrAf1q0V
e8gjVc+8UuW2Heaf9MA/+ovafqiodHYuSrOA8KaBuSZyorAYEdCS0TRCFXtnJvQh
H/rLwmmcLVySUjVbBPyIPAxZ9mJVbqS+d6Ssw/E7wqMBc9vSsKEuvxSZ6P8xjzhW
p18yb9qaoeoo9Ll5gHxNLkvl0cHb8P9WlLXQPy3Gas0fNnAOa5vZiRJDXyuVI5Dq
npT2mpal1wyFHY1hfMsxe59wZuDLMsxSaN20C+eldGT0RRNQx48GjVUjCjMhUrSn
pJUwWV0dPOpDX9pzs7V/T2COh6Du3OQ5ZxUVcL57Gcalb3i0F0d/77TkqWl3uI5E
j1mYOJ8JiPdnAuNjk/YehMNpd/4AyjO5fPmE/QfMSFpxzP5Y1T1yJTdS8zC1Wch7
PorcKV8Ebwj7dQ3D7tEZOzJES+Azut9PgKAajYrvuRuFfA0I6UEnpzWr1sKqKXCs
YziJs1z3eecUp676K9ZpoGRGi+ZVqLn5/vfnf61cXVpcHoa7Xy6QiqVCzrVRfMEs
KWCaGEiDY4+o+tAMvflunAeFbY8y71nNas4YZS2W7UcO6uTCzCC9ogM+iApRsFlg
Tcys2+GeUpI1vycY5VIWeVp66WZ+xoWQvqnU5CpEM6c9nWO9iupNLjRHjjfP2HrM
DDPTXcP6RyG7Ihgiz3S0g58I3+RE2tSbfIpjNRpAKn0OY5uHz9kSHkOtx1djJ83K
jorz2q8Pe3J67GK9byI4/PYqt/PEBAsxgVK6rRJdcDyLYhu2ai8q1AT9SVAXIHm9
A5JmtM+DPJvz1YvjdzfvR6mMrWkxceAQPNR07C0krZJolRSI5xqge0tn+TI+6qaE
WkyEMpl4Qu6e/guw7lUg/B/RTK12s8ncy9o2N3wKOm8=
`protect END_PROTECTED

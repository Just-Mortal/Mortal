`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Za/IxKnzW9FYBYoqy+NkSWpPeK0kDLoY1vwY/WAgHrnvXFdPtAQGyYGiHjLBZ4+O
vhaYT/6VxaRAMms74adoi6Tsi+sU8qd/8ZZyt9negy/V3CGOz0zCL0ZVUhhVXkBL
aLbxYNNTi0pYjJaK/BDyslfKllodWazSy99cUtIlFcjWra12Qt+WiZJ1dVXWsSSH
hre2GpxFTCJymQBSlZvItOEL+B8knEsjGfSGKmBihShFcmkB12nNvYpEabVcfl4g
OAYekx/LfzUM/yx5BPs5//UvQ2krCZ5oZJ9I4tkYEVYe4YNQnVanBClT3kYJnKlG
Nz940MjzB/XrK2+9xYag+MuxrF/gleAL5l5cyZntX/azKG00SthWwNJhBgqbopPl
GrCHjGRL2rcdFIBMj1RjuMCejsZouyQhLkeHKXUErhJDYEn34XvZsKJqoUKdkf0e
lHUI0bU7SUxEK/z9JYFOjXriV3nVH+I554x4AVTrp97f7T8JQphDo5/DBGAg61bZ
XBTW+WmrJUgscpppN9iwZwdQVdA/M6LkM7Bd0wMba29RWMGxVbCWupLR8MapoFBh
4t/LuWNB39WW2zdX2yxWyEYOl8KoA/NK06UGfSAKMeNRNL9wv5T3eGFeCy8FH/do
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYBhtluUPOP1gkXJHWxmwghE5zxdtv+LSCI8U6cBWZV31vjJFp6wKlzQ8wiiS4ba
xrmM3KEXkII/AAIb6wm315J8FgkVsBAPFbIzbsJdY5YW3QgGDvlQU8c69AccGQy8
P+hidywUQhlzFfc/ntcc6LNSY4wHL/QNHsXLAbrk1Md69oQg+vvsPA4nN6s+H8Gk
++9CkhBaDvdr7GY6GQbYwWDI8h1EVFZ8v9llKaHoN5FU//QkYGxLp/lL9hORR8I2
j9EFCNlSI2+1U+CaQ5lSiMzYPmbhLMWJ236cwKn0oG3/uyW0hXVTOJQrJlAY8GtR
hNxbkqP4bcc28NvcwZabJu5NkrqCz60CxGjpnnaiOkaeeMa7OocqP0Jvy/VU3o7m
/mZ4XDxU3z7lmdJSUQFJUYSgez1bzFDgkNtmWwbbNSLAdukNBVFJE/pN4n5phHl7
I6OsuzxUaW4tkVH090xXFftYhRjE/T8VgNhWs8qWrIe/GPc4DS3PRfpvpDYIpYNX
YZZfvhZZTsbCdO9CU92a+gyO3YR8cMsJLJCocuNcnTc=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eL8qaBUjdYm/Wk+qDqTcdbe337Qyzh5Q54a3d+pjn6Yk01bSEuH9baM/nT5YYkbZ
IxUi3c4ae1LQbatAmPDAEqsw0QkHSZmFpdgQQ1L/65D7Sjiee+50d5h0xRg9UNE+
+Z2330kszWjcbg7mTs+OXtnJ2rcpry8ezgupT3pIfnZaKFkqoNuaD6ixpBI0Ho5k
Ichq/WHC4qqkAigB2Sh/VuxZHF5wuAVJREahLK7H9B5rrK/tbsa6OsTLdbcSm26B
vw1+X1oIWB6dledFG7fpea0Yyn+wOGgLMG732kWhQ1pkkHz9MB0XSSWDD+0KnrXT
bf9pdil8pVNh8X8rld6UuGcWeEGLORv7D0wyN4d9jNaspN4CHSpTfB6umCsY/kNL
y84pIw+Af6SH8/bMSdyM/IfD/N5bk/0/XEj74cdI4hkY8iWKkATyYa6ykl6web85
ZBamHY5ULhuIY1iWwoKpeg1loFF7wZVKqR/aEBABWYCBed1/Ycg2KqrB5l3dvLC+
2n9pLclwVcdNgrlG2tGFuO2i+XupydLY1xXQf/SQcA2NL1u/XtM7wDjg+MYGkPoV
FAvkmNQmWY3f/RHm204DfxcXqJU+2MqtD9pbaicpY+ilSbdyEOTW0asAZMksipU7
KnkIBMPRUFmpTgXDd34NVRLDqELItmRf9hXXYEErrz4ZHvpJmgGzzW2ez1s3ovN6
GNNtTeTLEydDiVHaRf5izhYBcId2IW9HtjTNAjfsJTB05mBdF76aYl7kLvQe2F3h
WzzHK4qjL8WBGOViZuA2wNtV1CIAIt+ro2JohDhfmQ/rJtfO47oC5EPfVusV1S1/
45NnnTwueOCLxptqHCF5QLbpYr+QkAxo+lnQ6VeMg5yxvS6nfmpa2Xmi56NOxi8W
79mz7ZEYoV6/WjmsSWpG3obuFBdIXaLeN/qSJpH2pSSgTbOXilC2Y/Sl3JrlZSdU
8UOr60AGU5XYbYqpiS2TsmV+bwGJlYp1WGbiANN51kzro9BTN0zkGDKS39a/VPNh
z9dgTX/oN5Q8Yhl2pizVoPxhi7W2BuXLcYpUpOUrNwaEWtHsr37Qc6B0RXioy840
m8NtAwuRI2SIj3xUu1Ic6eFrYeEanORvCoeqKBucMsDptlEhQ5CCrqbchAoOeHm+
7vdnKNcAodrHZ4lJCdNkvDspYVdmJQFGL1F5PClh+lI+t6uulBX+zn/N2mW81W83
IbhYLGkdZiv4hICKdEn6A6oj7DUtqT5t6bc+vnH+SW1wPwo4P95/URe4tRRB320t
3fAlzyT2rluaaoj04D+vMkOndNdwBj14xpv0n8H84yeBCBSIeDB2Y6pnAPihyl/S
cDhPtGiVgPxBjAiwghQsk9VaXh8pWVxDxTHVpKW2Mw5kmuD6qeVGjblqmqzunKZb
Gpdy9KATZt/q53YI/0lV0GEx4w3FlsqWVjBDkl8K4oDjf6s/eezjn+OKVqUWRLWo
Nri0NQ9ozdjg4OvNSuuQ2Z1cT+2OBnxiZZue4JAxw+5qUKHehKfuZmI/cLf6O3mw
WZVQsumOvQIsRnonkurl3B8H4SL4pxbdfsGNHzmONLiwhHH54yTjT8VY7sz4FzCL
TS4ve4b/n6xyC2DojqLJ8jo5riQlD+ZFThgYqTY0CLncI2JIBNQVYGh99Yjfw8Js
ne/drMiD5S7ou1sqhf9AkQ+nCIu7A0HXVkwqkgKnBItjDxP9ph6GioO/TuB3eI/v
Al8xTcE2cmGdtwZNmDQmmE5b41cQdfpdHgX9VpVtqEfCdMNtGiWSoxCPO133rrJr
l/t/2uTq5ERNLCoo+AV6ZbbT1OSAtV4rS+8CY1n291ZfCqY+9ZJSJAXJIWpXqLaB
iNSLT57qVEtAiIGfd8dHgLzWQyDqhg7Jnh20jn1WoNfsKJ+T52T0nAbdJ4LoNuHZ
Qtfk1nZGlWc3lYTEaB/TEf47yekVomNBing1tvhYGQnr/Gx4CEAhZ5Rt3PqpynHI
t49KtJwuTACuf4uECTFL6GF0Trjpom5XTtYJ5OjHHu3J3bc+OEwGDQ4vEY6N8AHR
vUSwPaeUUcCpsjexa9yV5sAc74ViuBfczxCTxDJPj7uepR8AZ/oAZQLhdE7VKnbq
V8qT2G3+N8X6Y8VtH+6wz/WQjLdz5Xg/D363Vw0m8wWBSem1Xe5NhrUYgLDdGBHl
NxBKMbGBFkM3cnlIS32wUxfLd4S3c4oo3SJvyomFQQ9pMALtrTv2FOQy7mLeAMOa
vTlPGbroUFpXL9ZMh08c/t3zpyw0NV6Af1OIlCGAsYIxiFGRKGoNPlcUtCWTJdMp
tUp+JWeoctHH2voDYFoa99qYO6MVy2jniS2kWens/Vg5Q0Luvq01CKpO9u7QDaVl
ZfIe7uTzvecGQuRLzmDYEXCX6+22hYc24hlLdsiejo37MmsDzjUfvyTm5knBiLzs
H3HEACNSUCei/Wu9WsinD/NCSBzh93tlJ515tKZMJ9cFjQ0zmiRKXwrB81XmpRwx
PvDFUqn+Q1N6BZJh19gYxl+GtQ1X+3kD5hBph5lgj4in5Z40hPf0HhHtIQjbZif/
JxtDCDME6G5BiWMP5KQmEnsDLAOGwQFA9k8CpjvexRXJRIsYZB9I69zYIivn7hNm
K5n7vovRULFHNCLp0IPwj3YVSWIFO3YJJondyohdKbvj+b9ddltpLmn8h6E2t5dw
6Nz/ddKDVdfVvRqNsVzytXJTyPE3ZTRmudqY50evVR/vcju5D1QLVeedAL7I3aAJ
HBoGhECvdd2RhZC/gQUbq2T4MyqjjvXOmCF0bS7YwrZC8EKLoUh4ZMQsncy7WK1W
Vp0Uj7yZMs5pivnwiqoLiMJDV0aD471VYHFmNwXKjZcsHgzKzmgMZhuxjdw5hdTX
epsRh+8yOSC5Mqt2sPc9sl3uhISSxY6hE8mZGTHBUNzL666C5uk+6QPaYz4z/ir6
KZonvRMiUZ7L+eyM6pOowlm/XfuprqYOtpSyUPl2VKKka5nPAVcyHdSAacWpdiOI
2b8oMSujgdQ4MTAj11wC15gaGHSWnEj+mE2beCC4wyXtvzY2vrtrI5KmFnx+pY0g
Ps/m2rTSq0HoHW5P8pftw7ZOprso53vf42spk0PwGE9u+ZRxl8+qEEdqjvNNRttF
Q+EjZ4xZ54yYbvsp+gVJaVWO1sUc8eEKzQU3o23J+rGl1sXN4bmnai3nZrhr3QtL
4v91+fJsIrDc8SfWEZDTnynqOVr0enSa4dyAIuObx2xlaMMKlO+O4YwnafDqR5p5
xAbGkGYIyurItttODlGFDbBhcw6Y0Wa+qub9/HS6KgfbhNr2hbxtELElMBd20IIR
YJzh5AQCBeiVDqs/zoycEweSyv+xRZN8N+WAM76SSqiROeluKUnlHqD7o3MU1xgr
fh4uDA1tqvwBntVvC9Qn03TUCWN+8ZxZY0T+DjBJZR0YDTYqw42zWrw7kaqkweaX
F7QPfQpd83hmSgvyrCfFV67FT9hBax1iy9vqoxh0QncnNOg8UlC8EJhHKd/51tkJ
+pMvHqgS9Rh1j/21B44NKdHijc+SudAMUZ7SBCupitl8O/bxfgbW6/SWzy9N/eVg
VY4TdyMcREAPJWPdURbnIBxtxLU0fh7g7q4lDCRqzFpcBOZ2mkrEKXuZdX2f9N98
ZDLsncORKe+UrcRXpS8Y08Iq0bxnunvPAU8oqsDqXMD86SlMXMz+fcOWaLgurQqG
Y+kO8H/pz5S69sSRGd6rN9+b8lL29lx5xXhWt095c2ChkU0FF3kKMxXZ8dqz4AMB
ZLwlpYyIguEaJmGv6xKEwHXh6U0huCdOO4L6HJaEjuCs6uoiTg86bhACuVl4hL8K
XmCw9eYskSJrEiatnjdbW/yCu5HbdzGApZg8LgHQuw7p3AlRvpMgZ7QMzcUMnGCv
1wY8c0Fa2STAcrOCbK2qfmnoLNLLBmpsGyBJtAH2TTXZE3kn7oXdYsbQxljCb/N7
xteip1cOwXgHU79cJxkqaKJTWiUkL4zelyw29XaooKqeKZ3qO1L7VYjdibfleuDy
aHFJ/si0vqdeRPxvDSLbGO4amRgCzs/8MR/9cvtz1gHv5y/QxdMxJ7fmM/QGrbGb
qnSPxDf/QI014WErqcReVV1iJoPiNRtj6fjKsbT034yRzBP/9WvVjQKXYnhtgYOT
XZRLjNwaPz2ZH20dXJFQ5Aj6mAX+W8PHizqdLcaPMNvGJNE1QQDWb/ewM6q+axBX
KUKNvU+tiHIDrpG7bUFa0Qm5ww2i/J0j7ceyHHlucLE/4v06HhXrCl0wkUo2YcST
cPc4gVRMx21rgRf3axXc9bH8Pabq3WVRv4ZMa5i8ocNZb5+kSiVFlOBQ3Ss/TdVa
UwMbUgxhb/dOP+JYi9f0CaUe0Ck8zj0e1pUDxz9SPwiB12vxc5Cij8Ap3Q+tJRkT
oyEgH54RnW/2xdWjC55Jg9sw4Hyd7PAr4RH8Xwm7F3Rss2iquVO5BAV0BFVXSwLM
vQvsUdpSTV2SZPoGqorzCzwqyQ1Q1HL1eK6l4jFLtuSogzTYPRlsG8eHlN8wodS5
cnWgEzc+T9c5DTALTph3aQr+4v0y761AHWk+Xdpup3uW4OAaqJnrtCdK20GD0fPq
LkfohKxhg37j0K7kayxzE9smv5MZZY9ExGuF8MnP6z42YcYWTusNiZb+iiQvvaSf
FuTLv7DwDHpUEckhWfGyinYBnNuP3/NtNFPw3Cpf8NIU+XegcZrJ+hO5MArj9WA8
fpEPbAKGtYbfIBxoT+ejPisOT9KzXFPMUffHhsF2T7RFV2a6i8UXDYTz6D+fBTX7
bYzmoF7i7LjLQnJ97rniIISZ+nkckVYF6+QAabLOk/r9NG1sih7SvMJrFkNBZjfV
S/5M41ZzuCehOcHp5D+shJSLN4lBHp11CYyf1R81oNw39DpI8cPTg163C0Hjvihn
7MiheYfwvPAF1yAFV6Ytcf1xafHFEi7wku/p5kv2dQpzMMWTvb88l/q68w+W0cDy
kpzcVACdbb1FnCxa+zBYi2GABIDWlIr89f0avFiI+q0yneRnxUbq5qcXjriU7fMF
uCFMsFteHd7qxJqYx6gnxnRLCcuxx4jEJTogHTIyf4qvNy6CrG/zR+VlPP3aHj3i
oZ5yCvZ9HmMZI8NCZem8M6gKpQaP/+po5BVSx+MlhvpzjSePquj9nGRZ1i/386mx
QK3FFh6i9CGoh8jjAL3xQPe9elJoyq+XHA444NHl+7XA+YX9zj24GMAiJ/RZG5xY
0zYmwSfnYQaWL8J/mVVaXv50OOGziUrm9qj9QPK/AaPj2U3nJOZXUqRBg++26ZdT
YakRds6q+IVQ/64HsRY/8x1M3P/ydsOlMKKlwAA5l77eCV7Lw5zSEFn/CFyTJOQC
qy+wN5CedXFRUaBzqSlY3mramComDkw/dd2C2x+MDfUGtMmtG+HuMEFF3DitH8JR
6XyXfdF/sIO+oS5nbLrdQhEFnMesSzOzA5k/WTVOlKNUjJygqVvxzmaZAHbpP/6J
ika1AcGzJsx4EtGgexGrcLwq5TRGUymeeqsiDc2KwYV6jwxN29CTOZ8SfkK2nTYG
zEictaePix3xECRKxai4v7wXJ/rfORD36v9vuGaBgfoEYduJe5d+FbScnPrUN79C
jAS9iGwEwCQCfIlPPRPMz3c1U8BTpKzXX3YsWh00mi0c1oIAM4sDDJ3DsVOAKZQh
vRRYUWp/wwUDlSrUfHiQ1e0x/2b5+v4cKPLYcc82aALfshOtGCvBNkx413UUtFBi
uj3yxo+/Hl3eUE3DXtTDuaaHk2KZeQ9T8dT5SPOrfYrU0P5BdR+KHwtXT1++Mf+2
p4JM+/7S0OtuPoGKQujimlZv5sCOVVpy4VGziK2uxegw66+gVb22YupvbJWbZ8AJ
Cc7vlLCqK/3x45hE1KNvFng4g6KlL9nshKM9lQSCHFsZsr5a7y9OhSHgAA3SaYBx
4aaEtCfRfU+NYeuxwpz6WmbzZabGdP7H34YSBUHCzFG8Gqk50FMfCj3F4YQXjyWY
lC8TPMvIJJ7vBnCW8h1OHrvSXDXQgvNK5F4VLXV+NhuG/VOvTNFE7dWo40sbP4xN
8DADv6s5VHYjI3pg6SkZdpuzjuvcnTIOxdEOf/J9Ku9bQr1HunX2YwIiKxfLKguA
ZikzttzcEWT+sbCkQiDLoZjeC/PW44TxWxEfWt40JtVCOe0VvlKvmmhFwEcTSaqN
Am87bAoID5yF3ICzGOBRQ0TbOxk92e6b+JO6ECt128zuWl9VbmxjTDeoyfzvlmDS
yo4Y1Frn/u8tH8oe/U4ofrCr6Fjzbko+4AdbNC47Jca2XcLesrUc+oX9YIcrMHtG
eB6NNauc5rlZiqnpVqraDG0dwAEXHQQu7rCwRRXa0BpM+4g7rNeitnN+daacNjT1
GPhKOLHzVJ8xz1JH/QIuBWVvPddEODTIan0eFPJyN8R7d0L1gLZgEevZAq246Xxx
brkRmubmquqlRExEKVASyWWD3PFdbk/PqY0BFG+NrlMrU4IQY66HN28Z+YrfKXaA
r4Z93hooN6mdBbeKG1wHAD2ok87qK4TF1Jl2uILfrN54Qu6GCCmqom4Af/LrAzx0
0VT8NhJq+xHOchZttAfO2FUdVV7/z0mLBK23Fy6H6E2dXkcW1lHg0VDJvDzAHyQD
7w8staXQ8vU/Ysrg9c3qEcFvnVp748N8/CYOkez42/J0MRSHhg6gb2EL2cB1/ell
uuQSuAKjBgjlhfTkCfFvUkLnOnVyGO0eTp0vziuMMmE2MWmOzhAbkDfs89sp138j
OrDf3Vf0Xz8ezz8QpOGKq2dDxdfY5qHINKPF/2gnleFDLc68Vnj+wUmRKPcOx0HU
cZZYqXlVX5vjPNYJhir2xG85c4ZZH+HZflFbkMx8RKrPadqIMOUlfDhmEwqojXGg
74p11IvPQN54y79mIlkwtAEI/Mae7Ey+3W/m1DXrDaWFen3U6AeSZrsuX8WoHPHd
V8Lh0uNzl1M57byb7CZafGiPNK6FKzow8u+8WO9uHnhkJznb6Qj6QEGWcRAWD5jt
MHBa7/qIpM9ZYjgVdlHJ+vfjc8SosfG1NxDuZMu7T2Z7/xuex1qQjR3sFkpgH7t9
1DUPw+N4HhzHs9UyTIo4iXJxk13UtLSpAU/0CH9f7doTdZ8aBcXFGfpc77uMJYm8
0bkYCdg6xNq2Mb/G46Ott++NhFfQD2rVFo7dNVDVTa9dcF60QcBZEzszgg6zolqj
sAEqbf1ZNy4epzV7D44JCKI5ny0bv6ReWin6XVImGRjvGQ/tnkTpqmh2GugdizuU
1w7h3ULBEm1bThrJ9GkWkTvjgT/bcZSWGiP97YXa7UYi5fBI50qSFmFVWx64IY76
xAGoZEQpUV9SX+YUogwp5ZLGvrIwEpBlsnt9HbRAucO8pt908H7uLpmkDUwSF2Mf
sOge0pq7VrCi5XErPdqA0lgKCqsbtcVB0HcnHp7S+U4n5CapcBdfmZPcimC5mhIV
2jTh6ulq6P/2i4j72Bdug1g89YVrjZ2DvqPt/1gVSj1xXq35e2QoNlZg6oAz67Ys
lv4h7tyDpTLfpxWoVDCD5GSxwnvuVy47MbwOorZko6KTAEyHvxGrdKQU6V4b6uI8
t+FAerTFjAfxyh9XpjoZUxvE8l9X5KMaV7s+8lgDSZOVBDvK5C7noIv58m3JRco4
dxSbNS7XRTewtW5eQxrk4a4hYPbEBx18TnEc3HmMtTI9h9zdkRaNyJnukKpy3CYx
e61ukGUXyqegcxbWC5Y9vkE+HVu5eWwkzRpqOnAR/I+C+xuR6auqM4n0wxgffpSH
CMFIa4CN+mFNXwCB1J9WxxKLpK/zfZW4vOZhqgJ7SbJxHiREAcoPnytM7huUNB8W
tmzEdxoOsr/DW68QRy3LWw8hhsfqJ7qeN4Zy6+wvBOKAEOfv4cd0K45cF6xZCjJm
mWiVbPF/cjlc/sCpB3ArBjw3UpfdhKS3SLQYiKIjw8Rxqqyv1ygr0EVAqsGZlKcG
MfknV/sz/LZSK2fu9Ncd6Cwt7L9GPGCF1BDCbP5fC98DzjTAQlM6JR0D0PjDUl7U
mkAExK2h6Ht0S35Ct60SfYckg4rxhewaJejHm54Iw2JtvuxGrw0r9SJ8kdpf4bci
WLW4aO0O65nRhkLRUq5B4Mmua0aTo+FMWskmjpAMbZNNCieED3ROCPd6feUh7uWo
KF9cta3H27xVANNMh/bU3q2kObnv/nB6omOJCB8cjG0tBnK5frcuTpOn8fPBEYEj
dkS36C/rBXgYDLWIwlgYDKAJqq+ORFjTizXFvAVFv8Ce2Pg3uBH8sOn142hqFX97
v9zf4kVDBKyggE//uZqJxjsfmlv+PCLW04H+VCPv4M5ndlmfdT2V8DxlkGYg3pGW
7druBv5yVJ161YKfJz7sIxefopsBSjbDIqM/WYvqxTXJqhfzaJrJfn47s9WlVQqx
zXK2EY6osE56AvSnMXF9JeXek9qmaRkd3roqYCWeI50nCScuVMXZppRv/bdCFKyN
7yQfjHY5VNG3rRY6pRywMTMk3l3qO9XS9UU40KuotpaP3ltCf1qqNQNAFO67D3zS
F0TLHLZLriOw8B6aa13p6MAzpx7LE7hpi7kv+Bw4b8oC6L/TO9Pd+cTSlE65IHd5
xzbqbDRERB0dB9lPX3dODJHmGyXHhJ/iCYcVdqkbjZGw2qSdKbsxyVDSUSf9mSd7
t2n/qJ3LUBGhEcwWVl2Y9YRZdmiLRvI/JPLSlV2TG678uE+Zpw4WiN7GH1lyCZfP
RdJUOjL+z405NJ9k+Fd+IEB6eN60U6zw5zJIc8bhiLT5K0WX4RQRc3Npi29ZtRV4
ra498CYLSAy/t7Z7ZEWxENdawC6LK2Yar5mP85Pgd3Ye6I3/Tbytk5dy+e+Aw9HX
nKYhgKJKlDiwToq1vGmJ22RY8GYkJkziJ3nBGf//JMTXPuv5to/quwj+oxwZ+xk7
XkZXWk3iwXSkKOtEMefTigUH4VUbBLs5kdHzWB/4/4CCDn+A1I8RX9AJElAh29eo
bCaht04jMLBlSVe3w6fBXop9WMg5b8WpwHSJ3eDGj3YDyXxNqPXQlkgidgyZhWha
rY+udqJD5nlCUWTfNPEALLLR4Vj6U8rwnmHFkRcscKV6HQlGEtYNzsL4fsEfz4mD
BXV8/BY8k9MG3Otj/udif5vVlpu0ZUKcEw70bGQs9BhiC0EtJjrUYWwt6jtcWOeI
2YaJczCNM86d+pj3dS8BqRT5VaDUOgNemwZQLUrMXj25/FagZZ5SOJgurhw0nxkS
uNHnJZjrWomebOT4rp2xYjd08ce3/xfYQxZoj0St/6rKbHnAwdQJYhxSSoKFP6Zs
QKpkRio2kFbLVar744VGbXTI8qE7eItDWeoj0KKdCd/ng1hFZUl20MBMdk77qJ/j
eK2GRZGmPQL60Ll98tfTwRUtaF4VVYqwUJW70cfoom3cqdFHLKdl77+GPdkSpGnV
6VHbTI14p5C0c+9DMqLuWHO8e5MAzNE9NaJg2kWW9KilPQ4s/kzJnGCcaBNF/8BB
d5UNXs28uzOY6OwDhiw2eNtSnWathLCUVp7EoA39fLhWAq4NVxxVdjtnHIUdY2vm
ITdYHCyDE1BXcgCodl71Divucke/ryWTMmws/VazWrcbkko1dQrjv/KlMoJmD9Xc
lrOk5bzUmBEJP6huWe8uyhZzRueIfePyJEzIc8oVF+DSXk009WnGyhl60DsRFCRE
WnjD9LggoQ8UpGZnrtVoJw3L+66IL7TTXErJPHJt/4h4QYJlFM6hfpaK6Il/KjJQ
mI4oKakEkoWyQCJXzxwclUMxHmdzJoVzSV2/RLIlr6VRbZwWed4bGTE+BT9IIK0F
Z0f6H48uprxeqgT0RNBxZsjqXj5AhLcnhL0coc7nRsk4OHKJg6jnfyBKLBIvgBW6
yv223SIcf4xeXamOqpPkMiS6NJQgUkz9LJ87ChPoSYxmCa55BjlUXu9Ygybe156m
W2F+b1H/igyPUJJZ3GHsBjP0MXtf22Nx2vj5DpOXReTm79Mn0i0KM/HE5OZl6P13
7IIOsCtG8sLOuaTPTLio6WuIgyqHFDauYAaLUzgd2TUgRZvAwIp5pk1oPkspoRLe
NMVA/Qf6vAlfR7v7F7h15OeVeGsB7/fe3DuVhbprSdRpnRWNSag93iH1PEYDHhxm
lwkJgGxjJ94uCHotq+/authhTHLGfA6sSPLUXk0/J/SdSmHCHkF3yZ6LhPqPaBbH
l82PINVcZLk8sO4FHEejTP8Z5GrgdWH6Ywba3F/c/wDSAln9kuxPWjdtdQjk20VI
LfAFASuO/ajmncY8JIFT1QE/BR8umC946uqH1jl4Oxk5yiHa6U9rJLnsywCoBzGk
wBrLFlKU6vvGkVOh/a0z17sTBnTmKw0J51yXgVDO9yWiHyzFpl9FWn8nc1fID9rx
VUamW5ExcMtZ7GywV/CL04wJqhHNFnKKib/xP+pR8FXOe39zuRj02G72/cqkCTPb
7yzztNQLeMkiAJwKEEZiEMbjt6RUA8yec/zNAXrfIZBlWU4d0lQAPvk+yXXbkKK7
CEMv2y7agqSHd89+swvwVQGoTJUCA6Fcy9HnOdMtVKRsI4d10N/yobcAws/6S5AU
m6YKMQzrHPgELJ+fLrLGpyVfTQiFUlQRbnrfcrqk/8tULBmKxRci9yvmW6FDPo0T
Jnqgyk6lK2eyDcVr4PzB5pRQI8WomSOIct696zjoftQFWT0tqPWP717SKzn37i8u
IhhZomZSQRpgNhxquwV61TVHIjQ0wWsSFdaiTZyfNRvgi/X7FUtmaLrrFvNyzv9K
whYCJvye1j9BFOYqi/F5+A247eEM31aE1HbreCb9/y0IEoz2touMvPyi/fDr/aKj
ZdVTsRyunWQc5NT3j6A0dQfjy9MQmXK517ZM2bcg9+39PbJgftHdFo2UOyaJl/hO
M1F3NSblXght9yI+mH/tXvikFpxdh7AGqTROFR/3zoApe+9eTfdm2RfltsDisxBf
i25J98kwuKK/CnUDFZCtcGj0JQ/aWbPJvxWyJwcV8gOlZHWZG8r64/EayZcW/w3F
pG4t54XRiXVpLwXdcr+MDoYkF6E6PpE+A6mCvUX2v/sA4p1pyhfZlItvyYmYM2AB
KVF1QFU8DI6p+vJfNkKY8a1+PuF0j2ezhlgo+LD9fjD/JZLz5GvN/E1imCUTksOq
rSEap0YUEt8M+knXGzPm1g1YDdtEB/z5vTD/m6hWwDHi2kkm8Eyx/bS5vZCVFzOR
wCDUdaY0mi2aKbgCqMdebPo9eizG05CPrMXzdJrPzZq2EUVDC+jIs5kj9paNDp9n
TqWMjF93IrYQ6PiTyx1ucomL2A65Rytc4wLjAvUEqnhSzrQ4hQz+9emUzVGxO+7T
qhgoggL1PqbcynQIMu7ZVWqNJNIqsjGD2OrRClKrF8o9L3pwhIe2cwicVCu7pxoT
N4IVE7qC6QmN37OGxaidFYAP9Jaq30MYfs7EMAFOrKfZr9ZPdwKwNXWY4gQcilSm
O2Guf5AHnxmJc+Uep7oakS9ocom3xLbh2mbVl06yEGWi+kVS43Lg9HkCRPjV2zn2
F8jTaQ4zNdYD5RCIBlX+Y+wSRIwkHWKNP7UR46fN8/sN7Pm2F+1dU7g/2Hci5PfG
FovO26WEqsRqwkfquqSBFDpA46S8aN4OwTj7W6HayRvlYWZbMNw/A5P/QOX6Eo+J
OW4oMl6oOCf8bRKUyCr2s3dY8jb6RAViRlbzZMZ0RospAHlisp/j5bdPEvOeDMyI
ntfl8dDNLH1TjLDEtZaeGmrrjSeepW7DYQWCEdlybYn/3iOPNdXjClF0P0QNB5Z8
pMfNO8Sf9tZl0f3PFvLKs3thAsebf/fdOKXlKYrOsqpMeHK/KgSzOtCvcpJQPdA0
aCHoKPGk7hpP9spB9Z7nwvO5rIw+UI21dRarRjNd/jEG/51r0rZQUl6wzSkJwBQC
0st7duMrJkyHtIQsftXcHPkzynx70/5vKzSUUvRDCB59bn5xXxMW6uF72N/ddGGQ
qd8nV69RpdPGOuqyr03HqkSEjHJufI1/58rO3DsnZEkF0TY4sGr8NiwfItSbgJSL
GwjRWNifcHaTdaGUzdUjK8KFYdlf49JTnecFfo76pQRKtWvYaUerrGEBkoE9H0kC
wQbFutZOPcqmDEwvfh4JujzR8870a3nsnnBDDioOzwWFi50x86mEw1u/BDsFt+B4
iBeorqnxOs1QM27m+0q3B/9lvVsI1OQHd/zwcA7nmvjmnm7SttPktcNe4K00fVJH
JMQW5gU7XwvaLFrefvMQvS+ciJ3JdKMAjB4zmatZUG3lKHBezrRsfzivjT8HNoN4
w5R3px8Kc5UL58gua/Ir1dCCBotNdYVhdldyCoHsMclpYjqtCauuMeIls1dfsVTn
rZ7qx0EEbnqkjdink/jriRPoZAh1GUm9/krUlHDK/7xYnp7iNTYlOK+iPLaawKqq
C39CIkKm5eOA+lGXj1NEiTcTRwoVcKNBK23O6VYMOfbIyrv7iHi/5EwK3ByN1T0O
I0nztZR2jMppL1pN+Oo+EdO9i6di+jsomd27THhOiL7Feh6P8xzLu2ho5SkNY83F
+puOHl2fx6HiPY46db/lHOWJ+L/unuhYvQsJEePx5T11zlurklIVivO/a8QIyQdT
3umIClPqYfsJM9tmY2Nz2ItRtX8qRD34rvylvTNRX1h2Ka3gvmm90AQC/+n19aLY
AZCALilPTtxKPUgwqpOxrGtFqSEOhkq1Zosm0rGncqZBHY4woJC3BGgNBQVTb+ag
m2cyCNG5B9IeQviYT/cYSmWemtpHsLTC4nzAfLMpNZVikygMotJBz/DsjO/IiRE2
v9zI50F74zZ9Z7StbGLhyBzqwKXPFcOat//hmpX1R/wcVU12XeS2+2Dmybpsdsr7
DaegtSvSyotv7tDu3STgyFfsuRdE2xlQH78+hGCgr+YIYIcWj/KvOvQHZZWbE6is
v7r1iYanc5xaGum4KafFTqYnPyPFrpQdZq0eK1IovxB3Z5pajfHKXk48j/Lm6SMW
iJdjDjoB7NeAdG4ayUcGYhJ+eTBOIofaOcptXeiBSvQ0rHNaiYOBVw/MTw5mI40a
IeloCpLLoyylnPJ8srl2iVi5RPhfWA3Q1oDmKcGRKJE2aZBphrrK/1E78gTJShl6
RjwvxozWiBtgcL/JfS3Crlf8Azdjrpm1CMrK9ypKXR/xJMOiZds/XUb7lCulK8w4
RtWd78xMAPURcPPtwiNL4GnliFINPneGsIiU88U1d7to2NrzhpDzRHHvY2reYXWu
Pkp4W7rkFFrjb6HgRvAB5Ftj0HO+zqMiM1mUu2dOEL8p4rgY+9Ky2yUJxWuraTcF
NezxAM1f/OoKGgrXtK2SEoYMZ2YMQzQiNlFef0/vtfOvXC5oOo69ljbGEJ9t3IjK
KcmGsebnmsO/tNkfstJPn4cnD2umOC4KyVhJ8lqSW5wV7un9AS998hkuVxD1uS4w
pSUpIRO+zLo5sqhAInXZ3R1oOvMvzsnUcsEuytVOZwo4BvcMYbOlx8v/eo4VL1cu
jnJV4ri4aIsjwfj3GDSM19etARDXHNH/m5oRFgv1SR0SMhvUjZYX8Q/S5pisz+h5
VNNytrRIawxBv5Gv6YdnZJ431P2BplacXMe2uGurfJWiR4hllyeNonyiBhwefPnV
EtvqjX2GM7NnaivGiEliRNRSCAx69Z6hwjmfFWalsP92zBTZUk1OTTiKub7NXL2n
XtSup3r74dApQ0hxTy74I+AjoHQg2F64qDzC/vwHu1V6r9IwuRERwlSuSffpsHY5
Tezwn1nYTfXFaYNjFmGivNgadfcoeZCPdHkpIALFQ+hKPzvAw1NdYz+jxaa5iDc/
azawZb7bCJVU+0Ce9ZIZDCnmcFyT1FDnyDvN1gfupA8gc1+iHrUBEgpTwIQqXcwu
leVdhtW4vlXZceDSfefkm2ERT1UsVsWZiXH2lsGuouLG0nwjeXR97MxofokFPf0J
saE042wIChzbJPnoHwKiURND6y7Oyaz9+b8oshPt0BfYwTwuN7gt0llUnRPHHJBV
SS7zTX0BHOu4pM1bBwIGQrStiA4MLK6kWJj5nw4mKW3ItS5RdKU2yBJcDu5m6CQd
uh64e/nF807+wqTjteLY5qB/SScDicWoDfenspv2TWCwEQ0b23yCUrwMnLhPXQhG
DYwnbAjcgtCm0gTEP8Kb0KvDiGFXuQcpkNdL9aYcG3InuWDYt2nGpWthCJo703C0
kq3mulf84CKTXfJnbQmYvDYVmuGjJirfORjp3sbsYSvnJtNVhHF+nH3LWmKClceq
sIq0i5lEBP5GCz7Qieju8LhTBKD2CZSqB1xt2U5nF9zYFLkUhSjUTMyzqIThKMS8
uod9NJdAfR4mBqsIZGyaSSCRVlfX7WzC1deiKDpq1Kqt6tKUqxbIXDNc9+XD9DeW
NTffQEgDObN8HwvOpInbrX8Cbp1yEcPeqIpZ+sM3q0ugghTXO4QFAhfQsNKpKiha
XO9CJ57AnOyl7GVyUx+xkBQoPPNk5HD1K/T2VOuVLoGu74kns4V2c4R7GScS+VCg
aJLynTu8vpDEu7U9387ZV5F1T3lKw7E+MFlSmaxKU2yrOrPq4FBs1HRlgu5GBhSn
+2iE2oBOkhBbWKcHw0fTx002OjkkIzkBs/1jgg+lTBT3vgNJuPn0CTrzc/Mm1b2r
7ysGGnDQv+f8fu6XAcl+nUO0G1Mn6VYsQr0c3Zl771XNBVawnD1UdpG0W/eE3/yW
aVIkyqZpN8ZzNfYVH8PaiBlKFRWhQtaNb4HhAiq9Rk0tioVioidbMxOExpYj8Mb7
txAvqm09SlePxqjFCyNWseoUaABN/xh2OZznpGp8vsJA29YVGkZsqr+lnzuRtzJH
bjiyN0SGKEaFUdKezqVQgQa7RVOe7Jaenx5s7kVqePpmVeuS1GRaqcektkycPNv6
G/twhIaTSfUJbw48kUQFr0J0dJjy1Y15zdL82C4TVDUOmmk1Ew+Z2KN5nUWZbfsG
vRCmsG2OvME0TAxUTNnRbMoNTSf7jOue6amvjMOOQPcj9oCVq1ljlnOQn6Se0WoO
deZedp54ajPVBpwZ49fZlPC9JMuvyTPPnaehS1i/0YsJI8HgUAX0s8Xwxuv6T6D+
0UqYvA4YjZtyOie8ilhpfnt71Ta1yYN1/Nf+IdSM79iszSbn2HpbvIOKun2wJnyL
+hjgiyGe/WAPOQMWEwJ+C0wtjPxHRM2Z61yAIxqSzGKt3REwITnxxNPLk7xnGqOu
BHtMCwtn3mn1CJFyqFdpBgJTFq96XQ8lEOgkh7YZ9+mLIOWtIiBZo69t4UIQBhQo
Pz4PQ1m8eMQqWHn85GCYFPlBNvlZe3Q2R6XTEe56/FkU6quQDetO+KJE76cypgSL
+uz0QaGFDTp75ajeL2TaLJIjQG9shoZH5/AYxim7h3uA+qhe3h+EKV7rUdz3UhuY
8knXA8q15ynVGNeKUVASEFEYydzcmiJWbY5QPPi20gi9zFl14AnxFA4l+4BRUoaw
WtalEAS3bw5Hsi5Jv3dKu73kLOlv9k9kMlTVrTbXFbEBLSsNU4Zgqh7h0UyP93Y/
gYU7YAldSEXWxumwbW244PXB6rhGpIlEQOiOUfND0IDD2dBCeN76knFZNd0sKpxE
LckZRhxASMOGlC7800wFv5X0ylUrIF23a45G74j04mq77bpnB2fg95mJlqwbZG9A
vU+FgUCLDEh53Z3PrRgTTJk4XuMxOOCI6xdqLe9P0geVrQSLzg3LHClIlhVPHAFN
50zmZ4DGZeNgS27VzVpuICKitcR5Ga0a03ZqHHw2FEjwM9ffKSRDcAj4lj2gFxpM
L6GkOpm+z+FFIrNeJEIYUwJluhye8zyAXOwWhNzUfcnkLZYKGSme4gfGAHWMB4WX
c3+6e2z9Gl1gRUC4ZvNshAb67+o1Z9vx4pJ9o9/Z5C5qsKNjsFCa7ceuU0wrOvIs
Fm7iM06vpn8V9ZBDddmHZeWBppIGPB7wtUGNzqKcMZjYyVdN3cgEG3g2RteJ75+O
dB4Wbt3XtRRx2TCBmLU/bp9XRIgQyt1/S6nKe71ttex/o01jbAXe5J+JRvW99GJs
Mm1V2IbVaAObO7GUArkjazpkvFUwLBSWobBSilJVDvgpZGvmIdnfMUeKHDmbO6n0
v2B//VIlRDAlVTxc8dM7CpEjwnnkssdLR7QCwSXWj0quD2E9qChRUKuPlY8A4mky
bSABaniMtjgBbN1C5H1pl6DRVVFl1OxrbpbTB5IBUcT8l93dciy+HXPNeN2MXUD0
qY+dpKaYTAQZejuWirmd+b9p2dpxscITCYD9KsrqX6UrhDTRRDHHr6VCnYXRNVZx
MXsGSebeWgdFwvOLJq468dIuJtXpY838zaSxkeGmJqmnQzi5lUqBFNjNkq6oUZTt
gF/MU1lvsSHmB6CXSqy5wwD363624N6ScEYzdM9QtT4N3rMoeT++iERvLgr2oSa6
V+9dbHFVK/of9N39N29U3aGywJsXzmsnY1jmifGovZ8xCK1xAAs4nrGwn6Qbcn6k
xKUTPoD+MH6yiHDCjT9wz0gV8CztgO1nE1I/LmUEH5FI9ueNp/32yP39Nb6z79wP
yZL9J6dFP/CgVPtampDNfclbgSdE7VDTgqUPKEReqYzcVH1z3+gMl5lfVOg/6bRj
kbq+OudY+1bpwZb6jkUjWYI6E/E1lAMWManR2Adl2mGnF+8Bxsab4Zni2BH6jmGG
mCeJDMWdFx6kYmmOS29caV5ZytLZezXQURbAITP3lp0XyhWIhRnpQyovdLiin73e
QNn6tfA8VXaE4GQ3z9G6rIiDOE7ZtYnuIFF1tR4DN4BDvmMFMbQ+68PH7KdXQXt9
voJisZKvTIEG8O1HxtrYBuJrKmMJXomiwlpm4UG+KKl/2EMT0SgwSe24E6EGFMiw
mYt2q6ccE/qiFOF6nWijTbnpYVnFackZWj6KDQVHTAB/DFCXpx9rv7k+lDyS7vEu
nvSm3dPc5ExR9RB8QMKnIxCOnxUYJGSuBdxhfLoTjOz66d37RnYw0BEomhKKLKc9
/htbDgFX6gdOjfzIsxA0Bp5ScdL6TQkB3ifvodiO4H94NLdUAQcXQ3sefMJy5DQU
r4knBfFasnYue7KDQ55slkbJsrAC1J8ME3Pr4zwjJxR8FHwjlXYvDqumCuhMVeNE
PZx/fBW+Mu4vKVDDsHBfgt4ZzFZuggCQ2JbyLQzUjkR3IgxSoLZZo1rTJ0V02LAv
VMVHaJ1IH1WIs1gylPNHzUU44o4ylXQC2pS1m8sHrrOSNbpgdcM4sCfejADwGnCI
1JVX3l8gMCwZM96u1/tmvBnKeI1E6GMeTPJmWrM9XgITQC8aHoO+rXvri2U1d44g
20ErKk7g+V8XxFQxBfOA+wxGxHJ06a0UXVQGUiaf4bXgMtIUCI7GhxJNypPMthoI
C4giuKV6oBIZG/6/XyHWSJc8LYPlQFieHVWD9v/KlB60xGllXJZ3hmKENeRHLCVH
+2+UdJxxMI51emb0IO3r7eF08pSV79aVQEt3QPqja7r0SFZ4rs2gebKP1CVPAjh2
uBdH6SklXz2NbGuFNJV6Omcd9jIGC34PwWcxBdLbeCXqehygU41VJ+7J9kULmqc1
Kc86Kt3sCc0i50baGSMUOUm1A2sWDVPV9QsSRDQt3OPMD/E4nUnpweVYOGR0e+yL
/T+MacDk6C/h5L4nT4gHpAVSQY5S0MILohCz4VG1nsQeuPEIiettu/r3NA7LtfK8
9fnu9NE/DzQxJXsnzKRKz4Z0+knwyzahIolalTRhvSHW0tMGqehY76H+MS++yeDr
VKwUTk6BDY5x80mlEXsNFWxRjPQJsZp4BTLJj1uf4D3bc7uxT13muIXM75AC4CEU
vpBXWs+zUrc08KTEK6JPUqg/VaRzvsLTme07kFXkAr3Cb96ec5jsvZ68Lz46eSb+
4/lwbwhKRPM+O+Xq9ofS60GRcnJyGw6UNFYJTAX/wJLZyju9RkTECSLwx5vN3KIj
BOHQ7AbIy+AICszjuKPlFuJEpYOIGj3R27RS9XkV4lUq0Qzfx/R7UVF8eD6ZkE4a
tR+eAd5iIWKyCMlRFY/xneY/lvwX7uGmHWT+6Qiz2zjuULhAyRWD8XduHAJJvill
muZ+VQaBzIAvg5BvWvGgcOClxps2TVI3ejrg2ZeWX3w5rVqWBUfDtVByQMA2eRlR
auS3Uh+jiTn1Aalxro99vXUvcVpcLlQouR+QwTUNknA5A2m3gCPlqDRo4/mkCObz
5eLbW4ojwiG4p/yfVOkKIclNi2d7vwltrJ2RshqbQaYtdNrchwTHM6zRyOj+TeUC
1CGtP3wRKbkw9C2whvEp/MJdTgop4XofAS3vo1c4wNlRWG7MzoewU+WwIEc5Q/HZ
UMSLDGnxZc8Q4rpiUGIbuR8q7M8Mq1id90qrRHZ69hCg7B4jHF/9Q4ADBxfPJRxJ
ASNkIpbEmLFJrTTvY8UoK1/HhBFrEx+iZ1rFbYemWvItkiVAZaB/ubw3l6B/SXV1
iGAm0iZTyMf2HbPGcbQBQg76NFSoMBBPw5gqhd2HKBI8r9QQgxM5IxdDdERcm6B+
VgpMl02s08eqhv2hhOzYpVrJnPi7jb4xw3yyo+S+LpLk8I8KoxFXXGCJIO3cy2pp
RLiM8wLGXIOyH9mkcWPdY/lQvQtxcnTG0WCSCoUNK9M8d3OaNKsopjoYLQTSVoa8
+eojjoil1FT98XC/4SItWLQ8Gt+CJPKUOfkITEYivCEACnL9S2pnFbn/pfi4OHC9
+1s/wB9Kk45QDcxh/dCkpt7VMDWLKVh8OLLhabzPiOl+UtlcSSIyqBtZGshaZR6G
7wXqoEOD3y2uXU4SfFNYu304y4dAWSSvIXBpwZ020t9Yv14bKRm+hykW1ofFax8W
eD/A0/vlrfKUyeSb6TKD6wVZdRxZ89sMnRVyoxHarVKVhBKaUAsY2JwL14VGers3
+8E8/aCAfqFPHRuMs3mB6NDkPoLWHdHFnmn6JDJVBUoh+CFed3DKtU1fDrbvoiYN
Uv2ZXnyd5c8IJD/bX6n/8mdgL+ZNXTpYQECMq/Jup4vX7LYstft9x0lcFhzAbnwf
SFlBdSBAMHoF5zXXHgbrzAlSZXvJqDFWSa/Qw9rquIA7R6JE5pn+hp873IxXteS0
1RgRL8kYVk7pvUPRzEzsFA2fFERGxQWUPCPxYS0dZd7M+2+MpDJCG/2V+fIK7H4y
KgBVecD2lsqpjn6lG06H9+vv6Njo+f7pzP6jNpcgGgMOKwChx7AWd7uG93x/FDuy
lu0ShjpYLcw7NA4Do76XJQe1sO3kLeXu1frLC9SapNdNl9PMlB/4bxc3zQJASK0e
vXNedH9ap90v2mX3altXXvuGmKwK9HVZRrm66ZTZKGR+Be8Z0WusylNVKUacqLSq
8ghKBHLl5Nu6RgQCQ2sF8328SB3uJPJgYtt7qjxtMlvGeMXkDa1gCy2QTaaS1j7c
I+LdHHyuLWRNuaCYF6+YWwosVB0rNfoe1Ew+Mjx/Kb+mNHIAffTedKXCEfeDmQsi
XjhiZ74NIydGJg9dlwGuprQ9NwNNVOHFUWBgsisAxDcNxfVCm+0O4P65V1JDxvlQ
f5QXOdQeiI+eMCsEo1LkSbmv/TeU7UnZFTSNa7o5JqxZgSUvy9Tv3qhOj+uyET80
5LEr34mppcgSdAO+6ycRbcokgaHxVu/AtjFi69LLppLA0e7Acj8pOk1yXRkgv3GF
rSSvhr8Lwt93IK+r+zgtyeYcpqhVuA5IB3ED1x0hJymg5oQR4wIAnvK7faG05Eg+
9BjvFKMFisTFl17JFAUwb8sJpGMnIepE0C/4s6OQTERTUaRU0D3x9x9aLIWNcnFZ
Tr95867HtCIdIfAzGKMLuVsuKywchm8c6k1t+Cp+Y3TvhV63ieg5nuJmebtzpuIG
rLeuagPhx92V2D2qUNKgICmPOiN8OUqtNWAka7cqV4Z1RkZ47sb48qBXy3kmb9yH
8DcfD+nXnk0qH67hUZ0eiWNF4v7i0wjSHkWZ6unlK2PhSVeAD7hsmlPXHI2Pjvk9
pTk+74OinNZLnUy7iA/ImGh6gqn7axSXmaFUmUQyEI1TxG4cQwfa9oIYBl2n5Ag9
WghNOpyihail7W+b7N3xaHbaFKEuiWC5LvKqVDC0XMGe0EwZ3eJ7BWLFc9qdUz69
yAcSae3t9ceUgL+gRxfZf/nhuTG4QoxCK4vI2+Q69KFiiS56guY6UDBxStIgvLjT
Zd09SLkY+DJKf0URnRhB0GlpSDcgOoKEzuyJvuuTClilVKZ1Fpcv/96YFzSGb3pG
f5YqEjES8CALbxVUKdHzOXovYzCFCE98AKmijpglgJ9ueyvrPUKFs1st1g2zgHEO
DW6vyZoV19TPbOTp7C55bPT90Q/6MjMOZhp9tshVQBL8fIjGiGh6Qv3Kda1xZifG
jetiOyzTTlbiYp34yNzhDRS7lErKCv/LbbO6KkRhAr0D6zCDBhc/7w9Id7qxhi5x
fSCvwzNtwqAgWaPbaeKpY00KMZMjYBp9fd5BZVieZOXsTcxx6jwoeCSwYHtJPCGW
3cdd3jIHe4crA4RC9hRZciW5D/umNpk3LWwTq8PiiQsunU9V0vyBvkqD4ojv84CI
jcAwTA2Ol+yC87Sc/7cgZQBQhD1rTsm513hrlk9Bqvn1LVAmGx3eWoCC1wcJxuCP
0Lw+q2hY9gYiRV3SLDsLb4mQwvgpR9ROmd49jAMeOMLJPcaQpVqXkMbCE7dFiXXh
euvBQG5oZx6FGaxCA0QYmtAaZQ5p67BZ2d6Q1bgs9i9c4WY4o+7aan98NwUHaoIs
LNeJzbkz3qPWs5U2ryavKunMY7FUGu2og8Hvbvz0hOTbc/jSBw3MIZPSp7LwaP7Q
rLhiS4QgBA7/jgldzcIp/ZgRk2wkjz8BjYUyQuodRK+Drrtx5SemtYNTj6S089C7
8HSqm98fNZfgJe4fNZKFPK1M+nxqRM5PDsYyEYlHJOhN17MM7Coh3kBrZoUL6FID
nAPcUK8urG9j4X2PuRocbWFsF95q/Iv0ipxjeoEt/N3s8M54PYPjUUSIzo4ozbXt
c5EEGg5F0tLSK1U5ihMiZkefoa67B+0rRAkLXK02D2Dqd3qKclr2S/I2YUSddUGK
zH8LNQiaoXRdPWsej52+PRzA5BUmZYi8GAG4HjeDPbDmmlinUOo7liRvXeswpAzG
qiDZpW3TtmEnM2cv2iG2t622Pr0z+2cHIQst4xUoLIFyHi5wmavUe1m/od/ExZkd
sLgK4dZp4JCcFwanto05ebWxo79aIMuHxligp7435Kbjrn/NdZtt3/qNYfoZ9uFu
SwLpeFXQ09ZEYn9YxKJIgC4RjQJeOkr8TDsfsZ/Z63HdOH/mk8LDxs2kwEwL697Q
NIFOMLTmH/Bq+Db7McinMW11Rhsi4L3gWgsMVBzX900qzJ2R+Qee/zaofLkDfcY3
cZtlWnKlOn0r40XtkamI3V0zwZ8+WoSobj1KQ+82XaA/Qu2WcoGiRpugOhd/dKF8
/MackDh38iDVR0fD/vpd/XCZYfPjNKXLe+6LCbGjjD5Ne/IKtLGBC+4c982EkcZJ
PUTiAaHRlNQGnGEdcQY49PJlCwgvZRnF1UzU7VNnLMzQeIVuAO8xXlBcDG+onlwR
iWexyyyrfZAxuLV/D/502BRiaCXLw3c3q6tAHDImmxJV3koH3nMtV+84kAHhtlzu
tuSQWQ6aV+tW+ujw7van6ocvmHL01t3r9xFhhe9VivhqbyJzchqHZ8WDGVyV9Tt8
a1b5sYfaQly0LGmfcQaM0AbUcXOkuqLmgzOD/z7TARWStSyANMalrJwJkhxZPR5p
BQEdigFX46GdTwQ/0tRk9864Uaq2qnMBIcprQzfu3wFlHjzXlHL6RdrAOEoD/jXZ
AN4l0V8jpzOb2hPYDNL9hF47zuSttdElLdnV1BqpgQZ/u+pY365GM/G1LMALIN9t
pZ23zYvl3qGDDe0CDWKZoFTgX315XKj60H6VroDI0HkY91u66J0XbXl92eL4Y+bW
KsGTyf+ceuJrrEuxr7Tfo3ixyOFzXgdRZVI0Fp2DG5Yu0jM8phXkvL6U0NGUqoP/
fmlvIqWtOSu3fh7E2QWc8LTAhS2h7R7HUuUN04z1tpnbBexFMPdqgBvVKydhj6rV
1VDDfGHMxjpChajVN7TrxH9IWGFy9mjeweZK+vqK6GT8sbKL/i5iQVZZfFDc5HH3
DOUFPvfRbh2Gqj5EjIwUXbm/xmcE/GLt6qNm8ELwpTDtP0lq1PPnV4lN/1thHHnr
SFgmBlmDYRCj/KTDK2z6t0bl/Jh3UyIXj1pc2RJGme5bxJt5JHRnlCzlnFYvLH8N
is8brPC08BPC0GUB78p7HScoWlYbH6ni6Oe6LIjcn2lyeOA/Sy79JTdz2eSYYr0G
CPYchDi0ggQ9K4WAwI+SwZwCnJPtzlKlTIVhphPlDZt6hD7hkvJYJI3msLn1I8KA
tGprW0a3/GQTMFajKqILHxFGNbLWKd2k7eEXTsnZOYEU9LtyCG1z6D8EmqBGj+bH
gvCBs5+vtmapGOtWgnpzkYKz6Yen18CDMYEazFJS2GHBEfTm8AjEZxD62O6sBIzN
qKj6bfr9blyXWCTY3VLNJjXKgJpYz1KGCnkCM2g0GtxKgooBnRa45lF4j1cLqvSn
/4YKeJW4oMz8mK2lJ6UgHQ4BnC31MYrh8gIooMFFkFZOon31N52JgLhb9sne7mVC
KmhapOSdbIcl04YSynI0lO4+q4oSl4uonRLcwftPOwrvlhZ43Na33vn3UU6vKe+i
nBANEn9xYwIXKe71t0QlavyAc5Qs5B7AskCfx1fg/PIFJorg1Bang7cJxouvVDRk
8Woj1Nixce79KeHxEVsLUXJ2KimeHyYKmlXXvTgwQyRZYPa6gL1vdAdNtndy100/
MY9V7F5V/knXJ+pUj6vso8FVNyhiCNK/1JRYpe8XNfEcWuWqC7WJDt+Sa3Lqwllc
/CponQkZS69ovLYs38TT/c5CmUV3CQyo7T2XtAqNZIMD+2UWgBPfKISIG+5sRKGg
S8iHVeop5uUdFuMfr9UgPkcNAb+3PAWKtcQ2we/6uJor+0COZVPzB3a6PcqK2Rjk
g5EjUQL72LwY6ctInmEtW8525b3o2amOxVSls8TpGhgCvXOajSTZOSUd54/TKG/C
6dXmdOyByIykLqCmyizsGtwAosn4BiD+8Z/tW+82MruhPRyBCEI3AoLJe0hNU4tF
i+Kq0DbVVgnTpB3v0sbT9+aZrDYzLYjxlpd1aSYIUlcX8oyVUal5Ff86GWLDvdN5
IZwi5D62OWwDT/uyyzqmtuw/RMj6GnmjK9trA3DmbsDM2WQH8zOdmNtGWRcXRNLC
QvpMP6qlsQDyZZnZL2WGFo5zm9+TrxxYz/aYACod1M6LqvFU2/Jro2fZ4k3PUNks
MsyriWV+nagXmHPLihewF8qTMmUFvWPkXAMpDYvMg0W73EwqW3ChxVxGkK4Pf1rf
VFWJ5NQwgQYSdVraacoeQj1wQX7+IwbW9mbXztIgVvBmrzjGQ0+zC2MPorEhw/OG
bPy2BVPrPkn/v/HxoF6Qjws5MGSBebmyvIvhtXgDYLxRrGAqdVm9d/x8wu6KB5jK
wc07ExNz5qohHQx8aoT+amsawc6q1KiOFmJyZ4r6nHsuEG0koK6EjveqhAgoubh3
hdEFtPGVOuKEuBphAY8vuNWp68sGax9x59VAhswN8dMyn8FOFM6d3zeG9JJUgS/v
uQaNPvPXasd6zFekJ6B0bIwp5qXx+In1MRqYge4xHQSNqP8aCDNYKKHlRIemQvdR
GJomre9Q/SM5Ceg5+xU/Bi4lQZfIMrygUJHPTkuPjtEpsgBfrvB24GXkFPvVb2UW
d1g2irpODl/PCglQj9uffXUZdP6NLC3BVJha+scQs8D+Eg2xgMk7gGBHxiHwfpgD
QsU/Yk1x8Xc0EvNfw85jHgSMQDY8d+1+64rTrLcVHcADfdFFGspOlFPaOoBb6oOV
tSuzy1/Zd2tWxDhScndut3XV78adxHAb1hHokMpLyAe3asNkch7hifvjyDSWXXTY
fGKKYeRcusH3diKlwMnzvOMu9Z+DVThk3bvvP+kwsOXPUI2jyVbQBRnIr7LeqMxx
uoi0Jub/izqzqW2fje3ICtm5KjRFEjBwDVdnlimdvYrGTIMctrTmLiRl9WpMkEZo
nlxFHJQNl/2Da3pQZN+Kxl955fyJznA8BmnMwwU1Ja1D/iir8gaarfMjTTaz7j/l
0oET9cbIscmD/WULb2RHyUoaLJm18IELFdX9oecEYmEQXoQ7ERcP4+Bmj/bBb5GP
5m384EXMCM0yjsE5Zvhy66a+RPnvTb+ichQGTSc94xHW/WhwpErY08U/02/uhkRo
Z0kt4Z4DMYaZFgFd0jjeJentHJi88j2NX0FZv5uzN0/6oII3ZNsPzsnm2E17KMge
OuqPMdXd9C+v0+jbzjKRIu03ullb+SEzXhOXnl1bX9ZF2bdeCKH7cAocBSI5bxYu
jb4sPDJrE3egEdcSDzmlKUV9kCc51ASijbunKvYKUZcfV3XiD4o614V6+Y966I95
z7HYtphv/e3U6RPtNAiYGklksNAA6LJdg/7HesNgOJ4v9bxGmZwih5QkIiL1ZJg8
rl6H2ZuA2H/Vic2euwa5oys9KlhTvIAxW5n0fF4bhseHtRITaVASx5A2irs8FW8J
F6AF9fOz/uHWMWex/tAAwrNI11LB8DDaas96w5vG5LrsaTDRxAvNeN3MN1ZWpW0A
UHpeqtkE75bP1CiBTH8X5p1CvGq/6XR6XKlnhrM4fPe78hrgoFxIG023A+Evp10v
SUD1OjYrUphmKXATNAmPR2IM92SvI8A312oM7RSYQhEl1Gb0oCbC+t8fpP9O+KbG
k5GFtSQ3dFff95W6KiyMHZtvBQEcpZunI/6/psi8yX+0tWVnteitxn+vUT8og9Gv
DGyVrYzLKJCcxaadw+ofM4R9tfX5vpYuKOkjOGG29H9nX+1YqjuCBPyN2S7wMguj
KA/a+qiVgjfhzUUAfN3AP2rkOzgnOFWAHbL845zN/vIxVLQLO7sKQUbqRmsNMdAU
kG9PMIC9GhtUQdebkduiXaG7jEGBf7+1nehV5dQhJct9uWO16X2R1SXPNDdyk9zr
t8qHI3H9I0+K57gy2yHw3sIwA8DMREMhSPjS+78d6BxsuEFTG/TEfekWkQZPNGyX
ZFqZ+Z0CiPlAijLZtCtfI7umlqKpiobMzH82HA4CMzWdMVGkI18ak2IRYtzLNLA8
G9ZXfqRW4eQuKyqDASrYTXbBCHDGh5QJzG/6zhmZaWAwMh9g5NTYY4ij9QgEyY8G
eln9xehPpx8Kuu3Q6kj4jSpjf95qacxL9+8SxzaBXH4pEckQjgcke6F2zMO1COYP
05MzoiD5nLn7MUa93xmQrPIOzKVgLKELO83t8kKoUq56lmZvTXohJZOUP/WVaBCg
jzlkYGouTZEVh/QJdTUqJNjY6k1M6fKBmRmDQx/SZUl7ngvkMpBl4PCB92nsIEYw
X9RnELTvE4AtEuBhgbK8jpJv4CKOOThZ/hUMtz6rrcKE3Pb2y0CDTQPSt2WWwaxF
T9LiOXmHdKzCMXPzXU+eDftbBgOYue0QpicxC1KjMMI2hktcdubWN2FmOadaAVZ2
oYe8VJ5+qscfiS0v1hMYuI6qqsmksCAraLt6B6/0GuEEHnqorD2tDbHIrlE2GTWW
JnvFJYJzU8pWM/lToLlyoGXynSK7HHVx9Cf1BjgKSwC+jnZsrEN46ZkWqYephCzR
/pc7QAqeaprCFI/aLoQKF0B6xgUAmPV9WIoAjG+ue/q9Fkwq05DCm6hgjiEN1Wqf
8UkuzVJbnarHFX3HkPeCjCZYSZEsbSWMgJ99JrHFE9DeodF5Q9yoESBcJfbyJ4Hv
1sGCtHhMIJpjlI9FSLMbhE26bnl1BbmpBdccyoz2VsRGWW7fhc2siAiOKlmMBgpf
HAShtD9sTrWeI69ZPb55M8HZ+KaAKb6PzT9rD/W+TOf4MbBKqe7ayCTZrOCY0HK2
aJOuBpjba1mFUAgJSoB+PHncurgsj0AmAvOH4YlJPN06xrizdSYvB9KljhV+LiHP
Hu3rlOOhh3GX9Sd0CqGCtEl05FAPaoZTVhvoivLg1AwxiXgT+Zu3bMvQO4t9aCMP
sawv7WNWocns7qAqBL/lhlnHc0PJ88p5qxfMOAjk/Jsp1W7cRPp+mg36p/oIR+c/
hlrIimQbMq66zMBlbZuRF6VH7GWos3hygQxo2E+mVITQgLZXm6ue7jcXgfCLXXD/
osAPWCEaW/6+jRuDaWBntiG0G1lNfVu6shKQpDLu32uFaNjLcspJRLIfWNaqTBeN
oZEhb13dJ0cFBYwGMLrbT27SJKA52481onQeb3Wl2+CjjlCn3yyltDL2hSfluWZ9
V27NrkRYMUFbwPKe05G53g7xxXHXbM4/ilGL8SgKMZcA/CD2I4bn41kM/j0yPwsR
AJYAZLF278U2/HSiaNBJPkDCYr6NKNtgn+/p7ytEX3GGjx592SS2Bp+YruIL6dNb
FzFlPLOn/moHWI7mpWENTXto33Mp6ShDlYv46q8kiyIhijJKyCs5u7TP56QiMUsW
IXB0fE9I27ELYi0N1gbqEn726q1fv98tHYyujKMIVjeRjRdYXYyOODY2Pti8nKe9
QZSs5E6pimePkH890t5GtXDKBWv2rUTK8buWvm5ysSkI1TtQ9o68uuRUCb7JQR34
zV6jKioX9UhuDlX9eltHtvHwEBzj3Ry+BMYNkD19qi0JJ8qWrloap0a3kQ7rdXNU
Rgp4Aov3Mhfz6M5DlsKNDVgVcTfgtdv5znJ8zCsfIpxSPzrt8PZr/bH86qIFGloc
Fgbmw2GagIvY+y4v14PnFevcnOQ9AUUcKH6J9bqooW+1Pvtne8u30ifDuK9vxxT4
nfahlEmt2b7D3OdXX+eF575KU8Md5rUvq0awe7TH6w/s1hv+RPjaoLI/C1bg1kKb
gc1INarbZ1Ll4WWcPjz2Kg+SC0EXboWZLdfTIifZlEHWTUw69SViMlTiD3T0zq65
0BhSV4nTnb/vCj+NOu6UQk6/258Jhyoo7ypAZPtXqjnmBXPOYoDkAaddYRu21N62
IA8KDtiXznT1hOXJx9thASA64moJTI6HGucYUaFG1aVGGRwEFWC8rw9E4jzkWBHM
I9I+tfJKH9kv/wpqdUGG6hqbP3mWI/RaLkRbkXhyiXcVQ6DOnQwOlp4DYTyVhG7G
qoDOKHGPQne73znCLFqVwDUgCHZC0ibHFIB8cCx28tNaRDN1xr3eCMkLMDvjanVZ
k5X3M1kACE4Q8T2PwJi4Xj3t/IPpcotcdAzKxfkE8ki94dYMp2eV1il1nID12lh1
OFe3Y7Fd152Ace7jwlNtsdri6cRYw/hV4DkuiO4xzWxDVU8gSOQiEaeS83p0MBJY
et0NBZ5lgEWjBNH1CHPheSBxYDCErfrOAbrJnxFCirV5LQ+51FU6NzM+uDjxtrmd
V5W4R1PFDCZetG+4ZoDiNNz3rC02xYVjxyAdrvM3oWNMwbvAQCJyKJmcTgBXu5w6
me6qRr5yVS9qiW3E+QnbAUsba4Nz11hRZzN36Rz2kkQ2IZ5mBmerg3KTfG4kT/m2
1GWGE+TWAq1QorCY5aUHQid9PfBje0rnsboP+8ibque0Cv33uzRkNcRfjZw4FdE2
YhkFl3DsglUeEDTGLAgiCBh5pwreXAEYXbe+LuHmZfs5v7cMBeJjXkA/LnGA0j/o
6yQYEPi7000nHeTA0ASqo8C933MlIbs+9iIKwfZnZwoPmLqCASeAvYSTtI71vFE3
cnj0Zn/KUYFxekH7GMZ1cekqTefKxpiR4jMvKPXL9DKQnyMsDEeTQRXKUitlzRed
ng7t+P5qhNj1a+90nIJ9/PY65fuW2aFHwmy84GMNr4wIxNJlc1w289QdHFbNudP5
gijD4C0rhbPZM497LoCWBCjtImMq91gFT3AQhydYMgnqyKvn238avP8Sa5Lz52Kj
h7L/zjtwSgMjsq/xUM3wMeLriZyz3puWGN9KuA+Nxby7+xh8f7JbYJEPkvviCMWN
fyw9ZYsrMJF4z1Z44S013R6pJRCHHdszVAstuObTbHPCO1BWUNTq+kEn6JCZtVI0
o9l5T84BGbBImTlOPHVLKAxzzNYT1r6aQs0x0PzcnHwMTvjmOORa5YxSNZPU74bt
IiXr+ibK3EPQwzaBn+lUZYMvumEigVvyCtX5xpM5iLFRj0VdgCzqL9XJyN7vodY1
ywTPxj/9Lwe8PiJ5i3UyutvYZaCezhQ3iXlFlHPDldW/Cc3+KGQix0vJLPanFMIY
XrnuoI96x7fmVSWpojX+nw9RrNGtBaFnb5mtJlV+7jHBF1fJ3BMb9RMFATFK/yya
EmtwP35XxmT+cFV3FZE4miwyk8xRYX0PJkcepTp4ODQs8Z6buE8SkCEAVFfqXAK6
eAGi3sbHfy8/2pp2nSKsKpZIqxU78+6xJEFd/e5iyPfxMW5hwnaB3pnktlWPphkN
xgQWfi8rGFGtGxxsCFdMZzf7UkvCOPDxEV4bnKz1ytexN5f8mY9nW7KMMj7sgmtj
Lv3Yr92MZZfWy9x51HyDLUq5sl7Iu7EWtC9CLLWagtxGwt/SctIDM2YDqBkKSMV9
1PggKFHzyuUpuM5ffrly9Zr4q9iA1APk+9p6Z6hCnNBL8HqMUSFW4D6nixPo/n8w
gqnXtuX9juzYT/swPTW7UccBWVovL9KNZwbJ5TMbQhotN1aCmw9iRVTLrqwv5Bth
gVnAdSfZL/8ahzcM5PWmjvj2i9NIcglGqm/ebgaMsFaHHfvtmId5u7CSghVqZGFC
KvFOwtGlH6nkyHkDgHpQV8On74NpUUeFGGPiyzaQxp8XEY9fwK9bft6H5YaMw9YW
kBQaGUEIj3WnTL+z9UKl62TXZs9E8/sfGc2XAZhHZknKAMRU8Tn/xX4QnirJIqCe
JWqX6Zy3cLK3u/YXVV4md/i6Cy+U5KIiRliajbD8Bb0MQIDBtnuo3BqChoH55t/1
yP4QPCAFxV146YBeXdQxL6aBNA982W2VcYrGE/XxJJGE6OZdIUY1R1DNNQdLiMYa
xDvJbq3/fz+rIBXUnkebXx33tcBYBPjK7lX8BhKjvj/6WhTJiX2Xxhkp/EpnufZ0
0CK4hg4P2G8sO8DhfK+26+szytfEwFqvrTClo7e/EAy5voCqUoVsQ079D1WfmVwi
euicfxTq5r7/pgvm17lh17Utat91PkFd5LXg/4rCo+Wr+RD/0aAMlXM/GmWsbJdD
3WcZicsSwDPwqjXxY5MKIszcnnqFfGm6hPe+aN4FiropyKbYZLuSEcYxUWFnYz6n
EbYUpvku7vLFw/FNKsAgonKmWJury+uIcC8QFtlsyaqOPiM5fKw0nAjSF0Ofp6eK
LPWf6HU0DqQhUb5dRvE4ezpT5TDfcamZISeaASSRJl56zCM3CGWyKWu/L+zOoHPU
1Wfo5LrbquasmVgW3DziLETYwKerw7N8M3hvwu36FQG5asIVrV/TOmCa64juG+Mr
e/AkItVyxWbWLkq72LZcDlB7TFzZ+QgWk7b1kl1n5uPe0oiy0mWbYTrkOinvJb3r
KS0EpC4ygnNGMqszPoiBt1m/1puGOLhJ11RbWw5JCelPd5v+tSt8ormSHrC/O/+Z
USHwgMsiDuIlr8P5ch0iI1OS2yYlXDXOW3gR1RsShWH1FMk/AfE1IE2rEW4DoU91
AQ3LqsWn6l4TyBaA3grTFzxZEwcO9+OyjhZp1vhd3YfC8uTmHEmj6hZPLCRtXKVu
eA+rW02APhsgwDHL7gr98eLaMUyoRIkY7QZLfscrfccNFRdyE+X6R4Az+Bc1qNkn
7IyFoR/MNGdkBWbJve+18tPZf48dUB05OVkx+LZPHIyeFb9tLnNkSC75OXweXPWg
tOm+0U/s+4UhnukMtAxDs2DmFzOBW3C3aMett1r6RIORKyd6mpXTPOavrxCEB2NX
ElafU1rSGZtZn6RQxNIUgRBT+CGzrSoFTqP/Ju23uBrOhrBoOvpPzEJas2XmNzw7
Msw/rzSZLeGifmBKorQtkv3qg4lpCdwyKncdLOZaPbARsWXgAihqcDOSVEIQpXDo
Lyd9IF1Uvi5P6QMW6wayeD3elwcj9OZLTLqD6NFwbfsRNAtlV8/j5T22aJD+niGV
Eyc0JHu5KBSvc5bZVf0ZwOVHzYYYhONYaEk6Gk/VrVFsMsXUhe//VlE3DanutYbI
GofjMYi+5txC93c093E98COS8gTUpfeu76vb+aMgfI6Ie90YicQTsKkAfbg0zyhW
XGYb7C3McU6l0RyzrKC/sw8TSbEeJjima23g1l7C0xQtOxA48SjBFQp/iJs6dpng
D0rHkHtkhd4JCk9XRrtobW/G3XlnGaYdoaiNbksnivbXJ+ony6fvag2Gw1li0dsz
F1YQLJrFiWaAnRtK4GEvkqURP/2Xe26xTwrK7zrfGYEwHk/bZJ/b7Ho5EKYeohLk
ePm+8TlGkbD/MAbCr5Oeg8m+v902EejcB5oTFTWZkpbScWJTNCl9Cy9sQF1LHHXl
2uYVl5h2XYZW8j7mu58hfWvc+dE4VopDaUFgpPKp4TFlrkhDTrdzOBMGtdMbVP2V
dhN/b96APkKsUtlJg0Ozbkfa4tHSNtbhBvo9XjMjCLpewpJpIro1mqDCqX0gAOzH
A0pZkr9oCJgSVJ2JgRoycMqjfa9mFvR4O0lj2fXacJgPPY/T9VBkE9ckg0DJ7eA+
rLcSzE/siyvnKqoux3MJjhMTYLJYjnd+P02REKJjG0fDCyWSIE3Uf1xFCMwtQny+
1JPSXSQYauadjKSSktP8sybzqkt4LZwNzgdWUMqYm10RvNDlzsgSKS/OnNnRxEUx
+zlON2UF//cE/qyS6rgDlfPfQk3SV/bacHxVndqT4TkOzZqn34I79q48LnI89CXl
vJot0EPLnjmJQOHp9lsaUS/9DYxTjEUaxzFaWIYwNuYLKhPSWGYPBM+KpXahInBG
5vrOmJ4ONgZFdW4RwjmwgT46W5LT/Q+jr1fewS04DJYkrHykbBM+JU1S5SK+Ewug
Dyv0ywwFB/7orWpLZS6euFFF6H+X1AiLc7sMiPdf73frLpw/oaZHhfzBPS/eASdo
ewLrtJb5mdLjBX2sQxYXi8QxuGKQzeSTdw02q5IhL208jIDPvhmKtENqASBmR51I
ygGmhsfppE683rCj4hPn7aL9f1WTCFJRxolVT/upbBKWzo6iWPaJyEfdPbkI+MsJ
WLCVb/iVZuRo8TAudxYtkaFc/ZjjFIsv/SyyulzC/tJ+zUs23VIL8Bve+5VOF8GJ
98mCL+AjVMaDDb450dlqH5WKOIvZ8EvcpGZteGamOSZLVSp8rpnlzPAAK3KFLJW0
1xEepo1vkuEZ2IOWlk0T/XvHORBAjV3uYBhRWG5Qr2HUqjoRg60OpFosw9DIr8uU
/N0AvImwkf8kFntY0J+mfPdb26tItqOUMAazWCoxC8+mqcbgy5BhirCki6Uzjeje
QtqfJMaiR3qkBKnNAIv7nkw/JWlI9MhTnzTRg6zXBHPHpRxXN2EaMRj2U1YvM8Xz
1LaTkvCIS4zU4tV4RnrDvOdxaKpAYe4d0CzOONAQ8N0WFIzAfHz/wsJUVA0oN5c3
8cSv5zdJgr6tqv/lxP2IKpN0oEeVFDHEL9QqpO3KiFCJVU9z6hNpRgc0nXkm21gq
yGnTA5nIthfzq9GD/UuTmbvFOUoMR532g4J9carUWIMnV47uezmeCDKBDwI82h8O
h3QftegneEXSuJh2SCOGOPSeTc545qKTkmSS2rp+o0dwQ+/m38Vwf/UBbOB2UejO
aWllf/UpTTDJIt+VDhAqMiJVmAFzIFGljry0yqkkMc0v7wQcLVzmqhbFB5S8xJks
ho/ata76ObnAOF8N3hT07WD+Gh6p8LYRIfNr+RefY+8sjFzE/rAuZO1stiZv1HLg
UjJSUYI4LHcy2PweUW62tftcFr7NXaFCaeWJ3c0aBxsBCOMZLw+wdA10/88gJKMU
IYJj1QHZzAa+pO1gXJDzUQBaI1c4x3RDEz26A5c64wDo60MLk8AtLgXnwRCO3xTE
KO6lxX2zv9Aeb6qnMljlSfvqzwKBUUpn/txNOz63aF1hw41STYofDZVS1eUgByD6
gd0RFLTTg3EMBnGNqy0M/F3T3d9HWm0ABYJQ/2yF6MUvI/dDAkQ19kg2AZjSnz/W
1XDAx1x88Adwk13ZUCuG80xlHBMnqaoB9W6VKircnCoZCfhnSHLwtMVnTEHGG90l
7Y73tEdVTvHJT8xGFzLhOvp7ff63XSxvTeOnQoP2j0JN13u0RHIxUJakt8J1Aetu
xrRyjW3IPV2CfAG8pyd6px8/IcPv5B535SYnQo98fumuwO3gGV5lBqEg6W6Du8SB
aGqW8Wqd9Kmd5FVfJJUY0FzPQnJYjmlsLKiDLnRODg6RPsu8Db0TM+Xk1VshUTbj
Vzv6+rytFzQSULzeCdVhXYFkTyk5zlMVOYdJujypmwXTqyYlaWj6pd+RQkH77Ft4
jQN/sDl1vnnGVjjtlo/g2oskaZ/QgJQFL5lsqeMtWcePtsILJPr2CJ4Tr8NWOPiD
xIOGZjk/WKWACVDYiRBmLQnKns0ugRbg15K89C6esL78EwOEb2ZaP5Ung8dDRFYx
jgMHqZ5keB5irhXEklVdT7Kap+TKvF6KW9VygN8X9j2Va8c5a53H+G0r7di36tss
Gtaz8gsl8mxUxxnTAZcmK0CfgH9IjSJIbnrIdzXEG38sGjQg6phTbzI9ubqcMA2p
mUhn/iGhY2d91PsYqTX4NDcoAWQXE1y0T+YnfIquG3v43UiDt+JxrKfUNDSzhSlz
KQLTByL6ffWYDYHeHGPTDCcIhGyahOFvZt33mcQG507/67/VdpZRpMf0po50czqa
fsGFBrHRtKoD7+JhoRx1GrStUSz5tZ4rhhGn984VQF5D2yT4eAL1PhK/Ev8uaVHO
erFAR77VMRe66IAufhsoqPsbGwHRhi18lfNkrFHrPExuHKlHEU5rdaUW8nKXmOML
KmSreRGWj1oz9CAINSJTsmW0y/fGXcJXN4rTiLoh8PWaY2z6thPeXt7zWKTU005O
F8Tg5vN4nb0a8Q451OceFtdrjsgMVVmk6elm39zQLZwdvou9UPGHi/1DKZnSB0DH
UiFbOPT9f5PuHbmNAV7z6+Nl3zGy4IO3Y79AeU4M0mGdlLIZGDTlvpnANPXggmRJ
dDeHfgUP3XBo1jbV9BcrODRKIvZdn62v3k/uYnl33XRhKQBqABkmarPZq4A25pya
T/tKywcx7B8dWsJtx7ORPE4U+Uiru7e+MuNANym0hP+2Fyr2gKV/1J+uhjaFoV+I
JOh+zmz6Ta/nHq1KLq1QxfcFSVoEpaF7vcyFG+zF1p1TyX+BQDPxX8WMFDJiiLq2
8OGyffW7zlmmOZUrPSr5S3pi6STYUBORFV+RCqRuA9r8kO1TsOhX8DiLGq2OvxsH
3YX6GVZvrnsmcIeEcUSzMxbPNEHnciVw2O0fhC2jxl/uFyBuTs/y1ZB/kbAv9mq8
Ev0Yeei8FE2X3bM+gGnoYNYueo8OYQdnc+FVbMt0mj5sysNOzn+utbQ4c9yTmZ9n
N6htGBT5PZqxfZYgp1eOYpznU6w6Wq03z9wxZWDZK2T9USs8aHi6aYdIsie6PimU
dMnhaPyLUWyHTrPR+JCwXP9Jhi24rfitS6YgI8aTw7kC+nV1og4WvWAaYIKe2aUS
TPzhn0iIkyp9V0yeQbJKJmt5zB2OY7ELha3XrnymNqioJrLySdVSsSxoLJmHzJcX
jDTsctWFzWpxskB31K5sUIS4bF5SxDnM0sN7VPZmEvky0ZcJU89lT4Pf7ehNvirl
cx+zMudxBYrwFxboXseePMxY7270G2Z/B1+guA6UVfQzNmVjcsFeHpFDzqK0FqsV
IvODYOCN/oGupt9BBWtRMApZz800/ycsZ8JHzO7Z77e6ks0YO8sJgE44vyExrYqY
7rwCcdq8026qYQrAnYFV4PrTFPJ2AQk8nXwSSMqtHUbFlW2+WJh+RybDUSXOp6Wr
68Gqd7hzlNfWywi3wjtezCXlz15t1iPERsKu7v5i5RAUxm8Q5na/MNNc9sHkE0YI
dMXPvW/h0QJhf6NhPBHkV3sqzZi98xYxNtVfqvhWXqmke1cO5UwgkNDVQeZ4AiOg
S/zFsYN/rPOOTeZJG2au65z9Mja9+QHJv81djsTSsHSD6FTxjX2xh0HGeKr3u3SK
5gai2dhWBxf67hhzLZ/vd9pjL3voodPmoMJc0nS682FVTC2/6elPniOkma/MaTcO
l/COq5oNQJV6en9+5Q75gaNAQRITQVALqlKWB0weQ7fjovu77vLjRbJT1zMLaY5j
6wqkV57g42HGs0Jf8FVzaQxB4YB08T66V2Pl5TEs4Ib09fFp89Cg64GU0JbIyF2V
iitRX7MfHiBcHKHNu3gC12r2yROpuBFuq6fIfiCb/3qX9Dmi+JOEctxi5ZZSFdQj
iU9LOte9gwmV0kPV1S4eUcLKGXq5V3/tIAgSrqMrRbA2Y+MGMAUKcfvcvN6a2Gkp
ukHvIfZdT5wN1mHLS4wHAEfNYVIrQ20h6+SJ6emMJBTQ2C/Mt73gYNicr3UQcKjA
Y/8mT0fpv3LH8A+SWEjIzj5FOx4X64UjqGJVh3+wpYB7unj/AkOxF3RRxZJTmnlY
q6bZ5FkvkkwsGe23WCzXkiqhw90dvAR7IV9ZQ31yTGiNv//d8R4b4sbqXh1mdNlr
oPjGd+GFrtbZdfF5jPjSQQSHdovz79DRra3ewj8notdjbYH8NNU7wBQEmHftee4S
OklSLUvfQo7BiXYMYkv+z7MWZiIrY5+sxLI7NeDccQAAFtdovigE755hyJdO7qAe
Q3aKy7nyZ7Tlu6/doxDG6kMQlsZY+y5AfxVNk5bwk5MxcdO3sv1C8XOJxPHeD0Vy
Pq7RM7YgpnlTvxSx0onf8rmgZtknQsGHfqQhbP2/5TnDvaX2TgA3FFrbww44hxrG
5Fn/11rpqlrCfTffNnkMUudp+qFzrqeipkPfQ0E22z2W/EQeD2dK176Sn+qB0uZV
WfoDM+dgknnP7UQTaBCKl2in5QpfR1HGE+kFJmL+vFyqsYAG7OWCwYjXxsFtuft8
EjrmVUK59ZuQkEkWOVAQCCneTlJR17I/xh6C5zYCT+082YgIuxxkVOpNnC4jqG6k
zCfyZxnRmCS5J9pkKSaPia21rrDnd08XotgFEGJyrHJJsikyJgvb348SRfcvQ3Ob
xUKeOm+DqaFQwD0GvlYwsc2iiyY3a+JIwigbib1zw4oGIq8uM+obBZ+38uyrHHl4
vVXTS4G6If6xHXq3ehhiiNhjXyePGylVTRAkFLhjbkXFTwl+HLGN488940mYfIXO
ZoK3zMEg3zs89w1zTrWANfgsUbZ+19aE7q8gcWSljEIRVfT2fFEh5i3LzA+A05sK
UMs8nzSzVO2UxvVY5zv+Vnit+JaIs83jxFFbyE/FCND35Hlkz6PoMr4FmvCoW/0J
fl4P5Cln9l2bq3tatpLe4dWVesll6QCBEJe8tAL2ztEQtWVDrxfxJzT5pJnEQEcZ
Xe5NgMLolrdM5GvXevfCqZ87YzK9RGDCU1W0MLxTBkbaWu2JHggrtE7ztIViGCcZ
pmgCDkxzxvrwMx0hCxJuR8eep0+DzDIo27eYAQdaBSqkaDejr1myXjFcb91zjnD5
skAzU6/bb75ac7kS0rOOwF/HpWGjXaMPJrub0LwORBQoXYq1gIvL7gRIk7DHzAKd
fj02ofJJH+pHYdlaDLliKyrV4K+ssIe1Cyy2d5BQS5+KTeRijz1fah0ecEtNUpfQ
kknpwS0kMpPLADufkJUZ7EMSg+ehVOnHBcvib4qzg9haA6jZbWsAUAmIoZ5aAO2X
pkHqPpuFzt1q2NLGM5Z2afCjf+glniVHdlNQqtPSGvMrMKJLypIn/gawr2VOZ6vY
paz9hXEwbli+pXGHB6x3o/BPtWpcmZ2fd+JvArAxNWePKHsiMuuhT4WxL0GpJleA
LSU9s/vCcLiHEDVbYUWL7U+4SRtZ++evaNmoq43NkclUe/9fbDviRVs7Xtrw/F4s
te95DTgWdd/WF/wZhMSbzWxwTjGqzKlo4jpA1nM5peoIiVzNJqrlx4aY887rpTGV
AQUOJ4LjgQFYcedPGXuPcN+tGniG3wgdvAAXlflMLaguyRFcoU57lABj5gAfD0JO
cmqEvV43CB8KEC9QMaCj6ydlu0Ublq1nHCcG+wBNglAY3x9t0rV1KPRL/6rKz0vW
dm6PHNSL6HTDCYZLIu3FOcQw4t0j6MA5iG2SfzJmCR7zjaBCifgMg0Uy0erQ2TqK
a8at7OsG3me61d83DIz7YrIv/a34RpgnUwi6UYgGoyMOToEhacAzGPKPqDuBit9b
kmdxO6YeszZsQ2wR6HMnteFksVWgYL+6fPpTOG46ADFxhFDZzGdwxX/jojGUVkt/
Fi9Wh9UPFPVCmjxhaWcC3goObkqXg34JiDWEbE2lc1DLyjYdRsz9HR3GYxKc+h+t
CCFqVSr/H+jEDX/wge4tA4mqzYDv0Cnu9x/YJNu2uhAkWQzz+aFOTfB58X4MoFzi
VGV7VpNkTeNaXjEhlA0HzwduWyvlOoNWIRMM6XAa/ppZGU/Syh36z1x2MazUxsfT
Nt1AMphLHfiPS2FtQL4KNj0bp4nOZewMeqVOEGieIPaLatBAxXucI8B9zl/H/umX
DOGxvZJ27csQKwp6TBanRajS3jsWncKU9IDRS9k28izkMTT3Ib0/IvPARcEjmq3j
7anNbDbO7o1Tl2xT5or8mn4Z8IgyZO55aEE2f26/ClGowwARTJfialfMLXYK+WwC
56Oe8IKWKgvUAwuLsqfF+SSvn0qdJ51dMJLBwkdhXehqjHCfAAcDnmX2iWheUJ4F
mFNVx5W1rGqvF4lW+S/GXo7REpz4mWbr+kGkVu5k6853TBXfQWL/vlA5eX8y7nWc
G0FU3s9ZsAw95IuRx5j1C+/m4TcoXTYzRpJvxBu0Vf4xIwJNRwy+nh26DwjNbQqo
KM2dPm1X6oxCQKCOTfwwIasUkm9QgwU4PuZ7nXGTgjxHc2m0LuxIpUgfSb6a198L
8gRnSSuAP+u+BFxAuUdFAA1SbAKkJnVZbilYM/siZQRmlcDOKXNtlYm1Zuvn6hqn
ALPrzYDp6lRR8C/nt1STwj3n3KkIMvQxP3yYMltvuSu6cda22d6Ot7eNABdZ72SG
rT3sKPSvH93X2Rp0YXjNaXF/ZkFSkRRYu8gUyuooQ0k+xAGxVfeVnKvJc3To7tMh
5k3NR1/qfUVXoxuwO2xYqwW1+PxvHyhi5UDOwdTyQZUaauFm8HXrq+cMEnhisaal
JpUcQioA5AJVTvW0MV54MninpeiQX6iLT4JYxlM1dwxis56nhj3EUjL7dbuy2nGX
XzWRxk3vilv/ycma/oTacveNJMI5J+U5RioquhiY9WaCK8f8ujg/XCrKDznPyp6O
olRGjhO0j+KWpK1jBDSO2mTU3qFM4PATDY2+2KGvO4Bsk42uNvoVSt/yzh2G3KCN
Umzgjo2+aMVVMIiQqur131mCcN7SQi7TVPP6vWtajCXAy650EPErUozLX56BKr6m
Uzs65ihqotWHx6FtvIxbJ+s1+UbO99SHxesKUTac8Db8yYk3yKq4gqKs+zCCsC6w
selHArlKDzPgL9JAsRm2VSJg/T+DUWMTI4nlJZKtOW7dwsOLdots560Ah4ruBESO
1yjjvTo8woKDyRi6NXfxCKuEaGeVfIykuya87q7SxgfcACGVPmdemWv7is67vFoR
86WgjAoNFSJ1dX6qP/t2YzYz71k9WN4695A6sHghQ4qhbGQ0MXTDOEkVEau0/ppG
7q7XosbloKkgCx0OUc56Io7T4MbOh6l59A4i1Kgf76rqPrsmWANdXKv5wLiTyMpM
eWq8hKdcvfq7CG96Nbg6tExyIAUaHKxuQjwiQ1McDI0Db/PhN3/x/oIpNmr+gmY6
XTBsGEsHBHzP8FJM4443p6bh6sDcnME2eZCmfN0+qm4b9XFFuwIK4DMnRcGyaHxr
eQ6fJ3cAPzooi4uTx3DJi73LLiX3gdQEaF1gO6N1OKY+zzV/SkdyxDrfi22nS/3j
TJ2UnW6/N4XKE5trFKSXZEgqrhrKrJh5DOJvwsgMZ+knLxFvsRXtCpdyV7cxhKG2
tUqGw3tvKDj3nIuJ0aBAAPe/SISwaKZPnkK17ULB1xCGTvXTN2hglLdDXt1eWM1R
HDP+6hMuNDcX1Hk37we7Oh6ZhUyVQsIrzR6+QkC6hyrKvx6eyMLuv9mLY1ga16CE
ZX7jybdOPdY13YrHlIBc8qI5dZ1UVgY525YCt766NLPfnhf2PMHlE5LUhF61eIeu
ZHqTMTdjOrMrQfvty1GZLciTPEAByl/tWXfXPgnWnllGSG56zGC1BwjLH8Km9lTq
SZ5uYbV7J7OBjISwIiaK4wQYEJYUftcXZXQUQ2u9s6ydRUYiBVw7dTtPKIJZGHR+
3+neCZMj+8rUl49XGJUiTqQNTXJp69LZBCTq5GHgoeQ6Zdid4FUJRwuN1gTMtccC
gtbq5QCyJIu8IgY3ISuk3UEDyWARqHdPSb3zg38wmlMrnlZqm/iiXPgY4El+FXyS
Sl+95TwLxJkqhKv70/B/GR63MIGyRXONk1UBDluSVAMoJG4aIkLcYXmnpgk4PwDn
aoRITd7tKx9zUbyNX5GzKqCofV835TF6YQW6+mghqioUOkz9S5SMM3F+FPG3gX1x
aDOj48AS05TF3gRQoJakhY//PSs5dMZ/Nw0Z4CsLVblqnvLGzSzbk307LgPzy/TF
au9ZempQJZFV8FNV5CqKSPTn2b0Uiu5u+6M01WvJ3+JtTCWhxlIytEZWCwoH+SXF
ffRlBC9YzATqlhJY7pdvZWPFPymccJlsj1tx7kpjBRNPSaJLxpx7dmF7v54gsSCq
5pxakXFdwf0Q4Sp0Vu4gCscUrGmXPre3ADB46xrSCeR979AF5AFByTYdjFsa/ms4
9VZtowzGCh1J1XHNM6M2zpRN3JK4aI9U1MRv0F5l+almmvYvHimCmRf/TzlAuXi2
/QbAg24ehQurgjRFo9oG+grTRCQpI6EOm0ibIAZIY1dqlt4RN5D9xEb6wEtoFjCf
VsgNwH/e8LHoPQ2i1mmCuoOkjPP8lh4XUg+isOAauKkzpYNvBScmxRPlywim/TPx
tVeMzero/lqYXPqelGX4GPlE4gYxh3FDSgwS0/atZLz+CNzQ+ycxG9cUVT1bd+P6
IkGkjXS+w4982ch3KExJZDjCKxH9MOmV53ql3XAdqX2KI7kme8M3j5611WiPPdUc
7Y5u7t5PyrWDs7eUhGmcuwIGgXdiKnU4QIQ9BZHuaFKX3OUfkHDFpSrQMlO68TqL
vwt7c3bVDZ++MXZUfvLaSNzGWA3lJqxQq+etDlaxbfbyOjaFZN/w8fGh+XdrwiyG
xt6vKZ+7yfbMeY/Pq+nGh+xr0pdWFDadF2ENsYalb3kWxm75k8pDm+pSjVBsWQ2m
aMfmt0DwyTQCaixtUepsvBFgvpgYI76mCopVsFXyBJoBZcIrzGh0xNyDmtI+iNnX
5WZ1UTusOte3K2KJHlEfun591Ze6oWdZQRoo+4lM4wDNE1UIxLo/R1IftsFauqf7
Z2k6kpueuHutQ/zzmpopiftF5YsCU1OCRU2CIL2hLIXuGXdhITyh3Q8eoDTGsBhE
enp6IaqeLSz5LlDvMyB3Mu5xBoaTHBFbMtv5GHD536nhijqg2tZ3V5GVVDKI92u8
p6XEx8yfsBdVXhGbh4rGGWW3bgA1VTpa3XygH2qLrU0fizqEukgQXaTgNX6AdvM4
rYVwI5a68N6ldev321ZRZfNq6jKu6B70J6D0OmHMUJ1PUbxIpLOyX0KytExcrW4l
8z3tStM6zPOxy3wwiqSOjqz2UeXtxynDq9D6X45qsGeVRn0INfJ0BYPD36V1HTyS
0XRX1crimMCqY1i1vQgWWZhlUj+lptxHQk/4Mj72hu+qXwleg7WDYB14Ss4P93av
M5sNr3I3jM6sZ+G8zxiufuIic0yHllnesqjiS34F9cdUwByiltTfJEBzkf9nAUtr
ZR+C0hejNLks5U3CMH2Ovwedahy32gir1n5ZPiTXljONFRhp9DKaXW0XEg/nPvwz
p7aRCOohScJvthrdINgqQevBUJwhVKG+3a4bWgLjOLNQTuheClzh23WZnCq5ShiS
xZxvBnQI/HIdbdvGu3BB97iJKNO7vg00wM636034AgZn/XYDvV/u/2KMGs22zsQs
s/uaqElc5+p+zdBOmHbI4zCWsXT8JXJjcXrk+6WnnxgGHKND97woGXcatyYhXmsn
8JiYJQE3atLhh8euFHMvCzsvh4wahkLnbaO5P6rMi0aUcLUgKM6ridkd8SIudnvn
/Er1NxwYVwHQdbKVS0o5TQ9P24taHYx2Zpmdr1XhOtN2IjZfpK/10/RU6eCLVllv
MvUP+lQf2CTOeKxM9tW1wUO8pA7GTPIb8e9a+5R/jufvnmWz+CYhIW9fLlyg3/yn
i2g/GgKbWI91BHrRgdHKNEbpXzHj7Tl3BVdt3x8hFacU295qsLr2BXMDW4FkTBnE
+sgmzQ3MgnAiiNpZqCpWpOuCeeYVbra+ZACicVvBdxc7YemHhxmUZq4YYm4oxDuF
zEXiDlP3XjwDaikC7l56/3Bp14cDj37SuoM1gubht8L7TTt2WxPTCQZ2gxCHZQce
wp/KlzgH8nBRFvsgDZYUj26AV9OtMKXYAY6v4fnq4DTh64TCBcGHG6VjBYBDudOj
zK5nPTmdQcc5jaUa++BQ3C3veX9HvM4eIl5SA0XZIbKI4RvhFWU0rQrhi792FgQV
yxMCL9HnhvwGRbkhfZnj7zdj3zF1mIzveSRXgOE/woxnlV6H/3DyjiTv8i3HIrbP
i01A/iSYP/N8d+Le44yT6P4Oc2AsgEMMeoQb7e0oxrybPErD7MNsCUqCdXi6dNRB
wVr0yKyf3gjTF6Jg/TS29YC8rL7xi9uFeoAARGFA5gC4OcbELp95ZxweyldxK4ks
JwUkcBev62JGZq1hNpMWG7Lxza37vddwq0xTpzBPPDrw0L6rKhSBZmVUnbnxR0uf
yUgxc7nVWY1ireeI5BGAyQHK7+18Cib/iTblD91/+vbakF+ZgyXqutXOYzeF2OCR
WjX2GYdqo7LkKZ1jBAY9VimRDRpvFytadUf2hcP4PqC1Mez3+oYX2ph3qcpXMYMn
Pfh/e+L408P7HiU1zo13HRiyGEkvOaS1okglmfHm3biKU9cXFbjUGO3S4I8kkeX+
+HcSVOCGLh2/BqHGmojsgBCaMVq73sgKdegJs/nEURQQX9sojC7NNAYTW3eWGCLE
qss2y+URcTpRt2uBRpMm2ujSQHXM+FBZAOdFRj7j8jF9NZ8g48hAo26558arCIrp
l9/aphejlA3Z8zmcsAOgcz6NkcrCKwQsXgxJn8MlkmXHe9V+2jpeKQIUN6NCHjfo
fhZV5aUprl3pxvCB95FCoc6jvCft0y2O7PnBA7eRCiu/hlUifYr7PmWA/NKI78aG
0NMaKeVzYNNXisJsGVDPA2mGSJrz9iyB4Rirkrm7FBL671WNF9dhKZWQ3EBNTpGb
hGxQ5eJYo8XFmlf2GCdXinkol+tSqZRNcBvQ75rLEQbzktO6ICKx4zzsvFX82XVV
MkQi/fMfF0tQsGII1RSC75t3voiB3+ODMn0s2D+65WTT3Gsj3QcIFHJ8D3lYZ4M1
VTk5WNGtXM3l3nwHDyDJ4uL5CclfPek+DF9BgXlM9c/6Nh800wsqOXYlUt7lmGdD
eQJUf1sK7ig/CtrgaYO9noSiO+lNHGH8DiOFeffTSZQej54HU6j3Jyty+tCZdFiI
J8LgTrmTEla2rluQQ0+u816e7nsVK4+Um3/ENnPOly5nxUbHXYUORbkC72fw5xox
DN7TG+0sT9skIODMbs2oiniAOudW4ZLeW31AnOBZCyk3uqCn+Yub9uqoIEbVwT32
RnWgj3oGbzNb/wqCTXsWTcQfiksKDPAQxlrwL7Ukq/nr27r9l/fM+FL5jWQwbLNT
+C61yaImzn2NG+k45ze/5Au14NknWNmgjJVcuP8LZ3ZPxCPqn1qDHd/0TaIioniT
mmQLKy5jOXror1RU82MLcIo3QwWdD82KbQgfgTlHMSxuZArT9IU+bAjsN5JNG2Sd
RChmTeZSExrdZq9b2G7PbHk+D+9QBRAv3rGn0DfYvURyYXXD79A6rQM9gksEQRG6
7EwcmqM+RGk7wGvReu3qt+Hql6WXdW9JGRv6sj58qhiw6AFK/F9jlO0ud9IQCFQe
Bvm9nPzAChtmISw0iMNNde+ZDJXusKfWbYC1Uc7G3G6PZSUg/HUkwCcbd8+58FPy
EFE/p87NNmQoAxQ6xB9DIYS4W7iqyUR/cNcs882dOS2xBaCINALJ4eXPh7rdI6X6
jV0Dc4Th6RGm96ZjqaIDMiSmYkFZvHlEuOkv5Onvz4wshOU6NyFAlkuJ+FHYDDB/
18K8w/yPoDLMsjluH10D00ihlQhr8Lp81aisIMW9FNDR/HyhVF0X9w6XBQbjWyPP
/XIyYFFnWH7UTOPmycIZ4thTXCbRD71QZtUmaUVUOnyg8KLBYd7utFUPeeTkF4Z/
iJS+KBXqi/yXGZzPefciDEs2sjIove8IKLNYbHTgDbDnoh60RU2GCRo96Lf79M/a
vMfVLWgTb2l9ZIVo1WvAvw8L6u033jYfEMAsNkbrRgoFzevk3RtR3kTMb2YoqTMC
AwPujLAUIz4V2KJ6favC7XDqknz6bDq1DCXbjgiZ3v0UOLMu3oL4Ih5k+uwsErnZ
z/EdrgxaLLsmVjjb/pifVn1p5/n1g61p49iJiW/uYsrRUwxRocMq8IgAxs9P8IWJ
g1t6FpUVu/N+G2XLTnpSTSWKsR84EB6uGMx199ynlmwsTlpZwWjor17oMfcWaVsn
SyQ9wA/1ZEsMeTShSH6cvzlDAT3wraZym9Hqwbl7VRJaDCYLJyHqjwmAh/bbehOt
V/0VwfjBfMjyHNA0DT9MoCx4oHD1VItfpiF+eh3NkWWdchKuaWfFK1o7iIGLA4bJ
wdHE0QxRdAlSfBOf4tikb11RdhJrAfozdZgES4bhRS+V54Zs6fCixbPP19SAx7sO
cgVr1SorCw5EwBHGuq/NCqFUJhUyPYlhrbxC7Uz1OjeRSZMW+PrwOUoMzdKX4hq2
me8kMXzI/areXGAPlVOpI00l6R4ga4DrmY4++uOTQdWmw0V9YgWMufQ2BBPnfEcL
jQEZcJkZX7q+NmJkbPbWu6hGe5ioEt+8Qb8KZPL36jYh2DiZWKVjEQlv6zf34eM1
dB5SAKzk28wTF27PcOg5CDp89+cf4W+O7q9YFvBA9GbQ9wuq1+778Phh3gLnRAPZ
42+J030oDgB2TEe6nDaVsJg636nsSD/zmc2BgYlHFWPoXoD2Y7R8ljKdPJOv5CyU
YwaoeEwBKeXkogePQEt6I0Ww2C3D7H01RxAMM+bpo/pc+rGs4EOBkLyCHzrbHnuF
BQfAjtb0Cu6Y+OkMyDTnKpcctv11WWi8me3vBbJuZBudnl8rF+YV51fVmvNAl1mU
XPs3ffx9GSiVhUOjcAQQ6BPKGsOyIFn9vfHypCuo5GBYi/OpwEsHdgjFxh8APaUv
c7h4vKO/2K/4LShjYvf8i5O9QFGnhIMbvwfgI/h4Ead1Dy7TuW64sRFXDOvKyGqb
dMR0CivSWfRPr1kGOZxWJgs4pBdwalpCepk7KN5qz7vLQ+NvbwATQtt9FqVUxV+f
3+4I9+oRo2+IwA/cKb6i6Zzqers9uZudPWBf6Fz3HyhJnfL3nEfkgEEF1sEES/Zc
aFRSoo7Cg3ZY+LIBGFH/QXzKgSU3+D/J0m33bn8+fsW+oSM8cHq13EGe1ivLTj3+
0Ffz8lRATCgCy9TLZ/bdFFoYdjcBRZ/mqAIVEBW3fs62lmtqyIjyhcshms2jK4Bi
Htn0Wck2W54irSrhwfwjeSR8k2KkVYaYxxn0KgCDP+kvN26iEemO4kO4T55glpKh
03l6BnDFTvnX4Iv/m36/yQ4bSjvJ2Qqr1IyznOwwpsZ5LDvvtPqHo2HdA3PUUXq8
RZJ2OO53HYciyfoaZTalHPggfo3BuYpZ7Td1qLeHSAYCsVi3Pk/pzMMjQBGMf145
Ecav29ZlncOByUkhFbsxN0vw+jlySLoFPAKtPQ61GwVcJBFAshjXgyUbtqAKzHPK
7eMTExkWdOdOC9svVDEianJxpsRdpqB2ZAcOSuWleu6NPPi6B7n1Y9XV5UCvRzqi
2llB0diBU2eWjNeLUv9WeQk3tjz9JSQ2Z0kCB+92K29ZuKGpkTWBP4BUomBSBvQG
Qx/k8Ghb/610uMHXeU3NOaPmeR6/WZ67N/AwgExpz0pqWjV1kRzzyykkvBTTNkdU
oh6k5SdK2GQ/LjhGUez+zrErWSWhcZOjJOtRrIndYVYyV3lKEsBSK7Ojzr0s7dOH
9zna+cKaBhp+Z4gqX2UkmLvqcRdeqEgQledq2QZ/vJF1FbxzSFQonYLzOq51sUK6
04OteQ+31zw5HYmzaJOJ2GqfNyJmX24vTYnoeySlH9NDzFSl2JmfGKGFuWo9DSUU
KG9YchWufuz0QSOud3ZAGraaazg+0dXNxX2nyOY//kW/dkiM7E4uEEvTJG65NMUC
+j/sYkKqmmo2bEkr0bChJsEN5Uk98hODHxkscs7+EF4dkKMDn7/hOGzi/gtBI7xv
aKrC5fCacAI28Xnedvlo/xDTRzPfppYIMVX6L5nNAF9nIBfeEsOz9dW02DWTSzKi
nkR3DSRyAHxwLsDsTpVxJqUAb6FQY7XP5ty4H4zJCBZcbv676ZEcNlEHQVJPzm5X
pCBU7p7efQmfzVA2UtZdhxp9fvR3TwmBXlTAa0RxDhz1iWOkWAQ5r78Ze4hB/ERC
tcDE0TN+wayUawKNUSW9eqhSiuMgWAn5RZCiq1+XuIBQDCMFooYArg14nunFG+n1
mtk72VRgMY55jEmkiDVKSLDrr4URRbl0THeurg8t2N8xb6MD8XM/nt/e9D5Dmrzm
opkkcFKnisD6k3oiAb/6Gdoi+BSvobFOCKHF4bpaMfFQxknLIhBeoyImz2GVW3fu
br8obdWttR+0+Ld5yzUCHeB9IHaTrAH+WRgphanrKM5pJvNVuFpg/mafgCkpVFTu
jMqwFf74753V6xExq8zNCL/GOikhQf0Z4Q4LJeku1hRRlM1keXNZEnw3tj3NXzIV
zyf2gjVO7Nqx8RvFy3wzE+YdNNuR6u57qUjUqqdYF2EShoUYzpyjIiE1obAeoJER
OqMt05rfa4l2c9YLT+BT6GmtTC+BX9ZB2qKBfWR/skVbptpgGtT1YN5npYuCzDbP
oqZu83/CVb3vIjPuF9cqM/T6FMddNdCKOQvRP4P5PTiVO2DCaKi4zFxj+j8HtScj
cay6UbgK9CKre8tRfjLkW0QxH2JBect4s1D/YIV8ibZkRddX/4IrteigSMh7Nl2H
yMA7U+jK/qlXWIhUpb9l9q+32NdMcUYEe6DiICY8YiMRoH8EsETNOGYIUV49crKI
B6DqVNtQPDiUNBYwnVm0jWDX9tRlnDXtuiHzLylkDqzY5MayJsqGrvYgfFIMSiJ4
WYNb3MqNSdjphYDh4unyLBd40G/EKDeVOCgAhIyxd8GUb2k29o8wqA3/kU1Q/7O0
V8LNJ9418UszjHElKlsHjtpNC84RPMewiFfosEkFnYrj07neXjrEZXG8HWxkaZf5
0ZbrFyKYcYLV7V5nKI7AbHb1fpv3Rxpr8o5VbC/rq8asJg3N1UQbsOcGa/nrNuBT
mYvXMSiT+Ac4rBZfsui1pAQqQ4XX1SFuAcwQFb6+Hv81Gbx9C3oKU/zrbrv05WlI
gT6Ssbeieiz7bI0sHepB1QumrgWvD5A512KMYXspkanndkGsZ47ccHPiPTIs6NGA
/LuaBl/ehupVIwrobBYQRHP3PbIZBRGYcgnA37Zdv5Oe1UU/OTSyqYlyUyn1eEtl
RiwN0Dd6zpss1R5a1oaco1/mCnYKN/RGExToaKRAzsBABViMPhGoRqjZ8RKgBqeJ
x9RtKxUEC+hr9K3wXfyEKLXYTg0ApkBDdkJ3Ri1UbRxKrj7r7LKwuSkVFBGGtc5p
PVHtxIFLE71eGg7TwUl5RhxNaSJcS96BVMWPXUNbnFeiTOr6Mr1TQ4YX20MS0+Uu
rqm5cZisDd4NevImwOEfzNzCLzbtL9aLj8pVxIY3QADQjbgrd4lGrEkIBgukfLoq
NnBORrKD2gnx3cxSD7jJYrA1ST+zi4+b9XRfmvo6E+5XWJkVcVDA1PGDkpV4mTCL
KWP+vS0+q+Pm20y1cLwxKlOWWRbStob+v4VxXMAigjD+Th8G2etfcQUX5wooOtH1
GI7W0ymQhHxyBns2kC2WKEYwzxQ7nmKbn08jhRky4wFebU4aoIBwMpfU6fUX3giT
7CD7M/UyFk5b5YckYb/OphvZ3n72XE2MxTkK/LKyrD1Sv0RNYZDU3ErQDYgy3xVb
8eB7t0008Y4IQ39E1RYFNhyjQ+LBdb7caRvOGFVH7f9Hk8uHKY8AE9Js0P3L3uNf
hz7QteUR+mjaq5sp3AETgX4lHiXcg0HaD+xzpfuSZkuaLpPaBO2X4NDRQRkt0DE+
0DR2XmPYNa95y53Mb+6bC8uyKb8kV8Z5qXdH/781GywADVzsNj+CYaof/bj2uis/
lH7I/imJufc+aN2jVVMTuHm+S7JEpwPu25pjxWlAw1aUiXLJC0klYxc0tkbAFozR
UIxg0MnhzpVY5+cTL/pnfsdnBYptF+4V+Tr11SM61JYMYLCywG+0LlECrcgB1PRj
zxW0JDUsw56QUoO6+XfvSSqJmQro3xBCk1zl63eRSkt0HmhSx2iazgsM8R9CXrHV
4JwZZA9zA+nBnB4IOtt+3VlZ82sV+jWSMqnefSmAeL51z5wRNIcmq9ZnNC20slvR
CMOwtKAef9iVV8dUlVvrBeF7pXIdIUVFPG9i/GlNDg9fPbZ9emFtg045oi7ha7N+
xe4IRyQXc4vrc0YRvx1BRPKMQ2Bvmk3cLI9bcpkfwCcJ+qWhw/DBrcArPMe0QPzM
+9W8Rf7YUPjFE37IJyk8u6RSoZjH1GwANFJZWgHqK3aMFReOpn0s3mHsIKa2l8ws
dH4H7D3owKxAh8cK4UwEs4GKrJEj5kkaQZaa5U39vx3HTLwHM/uzS1PAb0ZbvHmc
Nru7EdGxzR5UqNbUM4S3IFVVi9rxoqh7xZ3N8fqQgqdA9Eod2Y7yVg+lgZDrCKzM
06rTSnFdUECnXh4tqfwLtGP8cau+UTsSllizOagJAhS6DwB3j9h0/IMKokRHNdEC
YYlKDzz+f1xRdASOdOPt2hdHhMjprQTrKU/j7Y4szFyNga/s9Vn2HItf1fvjuAY3
3Q6lgtcQW6gFpJyiCwgsNcOI1v7TDvs/0dFNLtZSaWsR6owSK4f4v34uW+anNadY
jwcID6MdpVJi8OYpc3W9t0jf3vVjSBz27HatJs0QgwRz372qMlKaFJhKMToqTNuo
zCmR7OldKf8DBIYdRLYLeaUcq4i7/UZ+gzX5MxUCFg14V5top+7Kkd7Gnhna8gKO
FcZoYnTJULq9V3n1gT8ASyRR/pFSgjSRUok2vq9vXJKgfvy78J3elNmHSce8Zcvy
J47VBozuoaXgvIi0legerVSRPFVl4lJQL+6Y6PxxaVJxrm1iPigdsfKJQ+0BLsAh
3c2+Y73slyFdSHQSCmSk1R0diWf1DLNy+9qz17ggFhtVysMKkHRhuc2vv6qMUodO
wjMYM+B1kriby76hIsmyZPOdqth8zYoCm0ZBri4G13FSZkuIJtalGWX3rYBZ5FnG
/lDGz7zwNwQouWzuEy9et1/LG+b7OlthbclApi4w+reYV6gYWqOOQswOvT/J2vsF
KthzAR5HSNxQx5mZ1fFo6gWamIxJv7sF5E/dWdYDqkk5dDLRKxIqZ1IZrCKC8Hc+
7niQ6oIQfB75EiOsiigiXImF9Sz+wp64Yffn+1JAwRolJTyLgXqJDpEAlcXwjzaB
5X90BUtKluozkXcrYIIByCcQtYHpmQj43zPG4VVNfGTZHHJ8oz+rYsUvu58RxlcZ
z54RJWvnN44/Ezotlv+CxWR9Bbme4TbG1mQuQavb/SkEGyaHStIC4404CssC7xqi
A7ajE1MwoVdRriPE5KhslAC5oAcCU7yTXTVX7ViKsvU9dKPjieLMZaTxLMSEMFt2
aCLhBs0S7uPYeGl4z3U1Y5RdvIUgizqo3AkW1ePxblgIVs52QgcN2qsXClUa8FnH
I0yKywakeIT7N5d+K+6D2F0Xq8qTdoFdiryKJiwH6+lQ1avxxFddFS1Of2pyJ97j
b6hKpr+ectMhq/WON3eZMBPUI1a4s8ZjxF9ivCqhpSyzcIqOVN670dM6A5+Tf6Y9
01wK+XNIqbAQZ9keseKeLxn5Dlpbn57xtv1EM65ZEoA7YmlOcd8bJcB8Ro9r9zyP
ZLjBwbaFrrS60BeYTMaZRj+jePEr7pMShGVuhtHcbt94G53WpFZmaJ6n48tjXari
XX6qPUNUcBWDySrgfrn0SrNEzafq5gmRkyW93a7cRrjO1ri31YnXBsusdAfmd5Ej
gzsltckPYuZGWEMLRUZzpKnLfVM9pH9yu/ju7bKH/M9EwChUyPtxRh+OP4C9wgHR
rhAEhEs55mxaBS21hWMHO+kNwLWRxG2cx4VhMW7ms80fZLXny1E8dUqZqL7UCVM1
/rQ5tpuyLgYoAdwdU4lEsgMbkRGuk0Hie+nIeAOep2LzqJ/zlMV/MM+uaIcT39GQ
0118TBQ6VsQ8C3U7fNuGdGs8ci//eVn4Y5laWQ9fRNm/F4AgWt0qUjtU3sY6iEp5
AJ1EOMSPUCDOzY3xyJTq6dX6+Ibkx6ctIFcwsVLHiqjbyyvvsE4rFmWHyyga72RO
zcxW9jiKrtiny5HnjUgHAg6wwaNfeCS/lXDe3/oXIF8dZwo5aS7ldjhH7FoONtBi
PSdE+0ybGsx/S1N2iqBNgfIhpLOwoXuwB8BMjT+OPw4AF3c56/9DD+1BZDxKH0pt
rBPdbqbY2UMImpWqnBjlGmRtHUIzB2KC6BYsXytiQxQ9Zjd+brWcy3v9Ul758wTw
IDWdy7vEzHoj2vRiKOwQhVEZ45Pp+jrlY4ZeSi4MZO5ZmpvofggOgoXRMYaOo2VG
1zyJoK3xA082rCRqRRjYcjCj2onxbuy2a90wViNFL5QDw0Z5cBcwGU8vnTlNGA8f
R1nm6jBKSwVr4M/VqTWujxdd37+FhEHSm/3GweaEMpeFLhoIXDD6gAeJKtmHY9kE
159ZzEUvEyo1Dr3pjQCA4OkagAaszze04u8BtJwLf0oaXVVu9UJG5khMis+vJI50
DglRQjHIqvzh2DtsVeSbVkO7dUzbOJay0TeAAkk333IG31TDZ9tbGibmq5xH+nrP
dsNKknYyGATH7dbmY1VWFuHS9XmCU0rAO0d8Y5CNQfF3NEVhjh76aJpicqz05Qtv
jOUDBJ7HuQ0z6PrLiLftEbKhC7A9M/FHnjfrkW0yoKow+SpeMmtgl0K9mre2SxKH
ajb2agu9R9wMvf9tOcnP/QuYA8Gg5QFdG9C6VyY+NktJ3Kn6EClJfoOfRL7fsv0V
FcAD42m9a8RiC4Ou7yHyHClsmiOPilTphWGff7r5jtmf+5UC4jQ7tPdwaiZt4jzJ
r+PUjEVMj5W9FRWhMQ4qZWHMooQwaR4Omw/U4BXq6hHMYEX6mcAnKquLFJjdNMl+
ZKXmwYf3mR4FcdSRBn7TywNwD5oMLxMJcZwXnzzAJzrxqOVPRKrUT4khIgDAGfm+
KlK9TZguAadyvXFRWgJcyoihdSoSoJP5kuUNe2yCRikQnDbViTjlJsSiPLTwe5fB
d6C6m59bDiW3cDYhyYV1DKy9bZsYaV0Fuzrt6bOZXomHF4YxKfeLkFyHKWI9CBeP
+QzaPGHLhaFKRunz8DeqerdcwPofmF+kCWsSZ0CoDbWdgtMGD0aYJHtLbnm6ZYmo
1wXV0vk3leaTUR0GYjaAWChopkIL51jBEuQDz0pFFpL35F0LhTYcvwEFlAa0idmi
/KIPN31WGumR5HDrt9+fMCQaY24rrzH0eOPP694JOmd2t/jeiFWtYHYp9EmHq15M
9duQV6/4UCdpvmgiXQp15cKftjzNERe7uxESDTppFnCua2ZhPrWc14fnCqww1WmW
Fs2v2wrxJtlSbTNCUSwLfNAP5mFfxUHbVHKIC6oaEXag5zzepG1CGBqvrxu+8lUw
8aSeRrSzGcNHIWeMxoL0LsC1cMA8Mb/sN6GfMM+1TesciV98uKJF2KGPZV2HJV47
Shcv7Bb/TKG3FqxJTPaLUumBAc0wyOvBfcr4XVivaBUyRiqw8e+I3WuCEr52hbas
11csjM8XX2W6HyIapHEXbWS2YGTmEAgLIsq+sut6XnHP5eph6k0dDrvl4/b8FwZX
RhhXu+8afVcSqB+0lyx8YRnjgTTsuJfzSK+Wg6DP0MAtq+kQUhx5mJge+RKZAFDU
4AWdMOWLzu1NKb9sytW+GdQvnkRcSfH8EHFgW4TrOO0feaiIccJrAruoiAij0lcm
nhyoRtQfTv7Y9lm/Z9O2TzC/iOxpizfocaHXJom49QGspzkfOvaXhdhdBeo6vPvP
719IqbOMK8qVY0toaEMt6DXoPkzR8dBUyft4JASZveAoiyDYELZ6JEFeBqfV5qnq
VbBadLVWT1sHhlh5WiLBIUunrfWgkyJMDxLcK0A2uE/YTW9Q2Dhad0VWYg9tt0HT
iVJY2ySSW75eM23sq6o7sqSCcAqKu7Gl4ArqrI/6j5AXIuGev7Jndu8fy6Gsu88R
Cd2PIPWTs7uoKy3YKw9WKWMxI+cqkZszl30Z585rzRxDN9odJI5HZqR1VsjGHNDO
WGW6kLpHEZA6SkeEKJJok6fKEpCVS7CLh7aTOgi50sfe/39xb1jjGzbxu8BdZvLo
x5qGMSXjxKNHvf6Ay9cIFyRwK5j3GMW7pou0BUqPuw0TfccSr4Fex5gX2GjYlwc6
O0Lek0o/GaG25KSQi5R6GZkHug259GiUJI8CYBwyrYPo5h8mcw9ZIEumHmDWeByb
EVV1ZMW7nKNDVMD/WPvwA0r5TPZzzAZZzxAl8nKzx+C2cJLsjLF5SWJkyz5kybAf
7Ec8SOHBDdTE1y353j4gZ1ziF1EOmxVyx5deVTFyBM2+IxkRZEZ6Vn4Jgpwqjz0y
Ps1dUV04W24DGzJe0e/6rX6lGUZ5EeuJ7S9DYEtI55XfdS00m1ubfdV0mQPKAwaR
jPA6SFCnSP4XZ2OxPbuaG8zq+wGtTqwcwIj3fbzA69kJ+kpPVVk1QWtiL/6vr9q5
2O278ji6vUYapLTrqINhKaqkF6Uw7jihy48+oW1YMaJ7SDmSMWmvQ6J35QyRMPxD
khjetnAG8X6oAuUYMVUyEtRR53XDVjZkEzMrtKR0+Ac18rp4K6mNkm0n5/tkW25I
yseMoZbOWz7zdoUoa8QYIw8wUM1RUCsxoa3BD1MKSIOjasQ9rbNKltjTDZqgvGk8
yFzdXY2BDjOXg8QoYVP4JRTbuVwv3sGDTh+XlkcFczLgzEUsXA0b58CHLxK1Teqo
c4QY8o7LcQ1MME8/20YgoggCuW8TbxZA2nbAbtgS2e0z+RfkF8scym4FqtPRaa+h
vI49UhCSIJTK8Q+6m6EMTvzlQiANiplCBNBUClg5Fg57csX/mt0H11OB22DkHcEt
ACfBiraVQRGCp4GFpZCjbj2IUURHVxRdiFnfixAid9w7n0PN4AuxbYJYKk5O1fSW
FjsZfja5WfVeyYf2SxnL4qtllwUthwmixqvsPvP9i+G3RRn3MoxI/m8FF5mGVvb3
bI30gMgIaag9ZPdC/C5be2TDDmmgKE8k95ThoVMsgLXq+qWYwLAe8jvzbhI0zFd0
CsifxgvGc5ldCAdP6WHrS8eJmNBcp3Xb1VbPkTScfvNtqjFJNUg4e7oDP5K0PzUW
YLMwo+tVa7kFYChDa4O0G3BrgMK1HxUzpZ0UCkU5meM24eqHJtswhKxWICtFoE1B
ZFMEs2nh7nj1pg9EhMq2C2U2swj9IhEtHt45tLhsZcbeynueDbgFjrbWEvARp1hn
oghjbdSUtaDYaJJVMtlhH16a3HOzQlbDryzXYo1C1h0xoUBYJXgLRkgpqYd83pBa
CTvrl2pZGI4DPBGUxSM+tVKOy1rgpgT3U23IRpKcgEx/7ockCVXyOeaO4KLUP4MY
CTkPYS3zTdy/o9xz7+J+UO6HZNgkwrkp31sRyChlQL7n+hjXXnU+qOu0pbXtsDPK
O7FvLYEEFLp3QpOMGMHgkN1Ul+3UbOIzOZ0W7YJjDSMum5IiioaTrikOnH32ALXr
Y9JnNWuj3c2s4+IvBMLxGMgA4noMfck2CO+ZYCVi+13tNO7iIQgwCXWAY5uoFBTE
pfvc1WIWrLvYPm1p/CX6fPX62m3lcltuAXqqvWXZ5Viqi07NgcF+Cyxz30opwAh9
/DZ/PdGAwA5W1CEKNgEqAcOSjlyRcsKm4KZHxF/2QOi64hTm15L+SLT2rgSsyF4R
OjJeZciYKDwItYQahapNKplxotswJWGaVHk/XEft3gEP6KeBVuvhk7NM60jD9tjl
MrFCKNXQbrCrw4ZIruq9Ju3BemBCMsYiqP1pWBgfxU2/FQAOMZRdlI0QIWaZQ0+a
UV1cXXP3NJA8/qMINSZ77bE8VpaEEkpad2ZxMOrsGosHxhU0yVswdOCDxf8oooSd
9OVjukMqmsIXyh+K3uUaDKv33vMic1mbiB6/XCEvgi3jLjSqZw2w5efHXos9RLV1
nxMkIIJjZCpvmjCx7JRASj1PNATyFvR/CsE3kRRB1v6a6n2OEkPqHt+vujJAA4a4
Cc6EAMC93nMRwS831aih/EneuLvJIE4HxXpmkhortkm2wh52yciZDy0lOCFTu6Ci
8EJO8617Be+VLfWCa4yVPJMfZsiqW1a5SwpmyQd3TPsZaFYitaGk0yIjHrI14FHk
NhX6KgK0wxImqmoHQn8T6Q9yX32KJs1cvjqjd5CRtTB5GRgeUSPpQoH5YkeML2R8
hVppZgNU+4SHU2ABDbqWgG1UBqRTzlktAMmRNYlyhIetn59kgm/dOq8rDpQhnn4U
ZH+oFk29vApz0XsMUQO4mYsDAvfiJ8v+D9KtsWQhnen43Q53ZNAVaoLFoOIxCpDQ
TUm3o5zE+SCQVqofue2tfJmuXPDZjXxPZyKghPVBwomEYBbU5TIv/Rja5WEbmSsp
rpK2gBXbvmyyBVRmqaobDIDOtGYk/Yot0CbDxXlI9uibiglR1PeM0sNivu/QhWrh
8iFIuuVcrE+sUZj4+YYAw/dFkqxLduGyqUvZedOVS5bLvMua/uN5YKHKfivvx5xn
OiOwRCwsypDyww00iQctQF1JnqtoXgI7fyPSXfwtfUcpu1TA2bwGK8FLnI3wDH/2
x5EQLbCSbcRB6TZ7/8Kf5TRCZjOG0RldTidSswOfSomtLnu2jqqR5qObgYcw/mji
HVQnY+o4qi3/sv2IeQwaPDUZQoxdDqfaoZGnqqgcjwTYibPcEvFeCYWHSn99Nx37
u/mu+1JvXDlWooiNWf9k1ObaXPmAQ0BCdmGQ3KEpQ6o/TkfF1Njge+wVC7vys3mT
0D2sjhRrmoEOkCwA3FjNIsoqZJjpwoCamFlM+YcZYB7ID7HQrI5kpcG4hCIqWzby
MFDEJIXjwCYh3cnpxyfrQgdPbhElO5E/KAmdgD5UTXn12zX+zsBxQYd21q8bsfqa
R7P/WOMs3gQPRhvyHQ1VFzZKM8iFv5VfVuEpNnCFSnSMZfRc32x3LqL+poa6azqb
kDfMvnr9dF7mQHZ8Ny6lMw+SXjXETg9824Po1SUG4uQ7WimJhD+zNbPwmJkyppnK
xwDo5nlXAmMNtbOeENDKO0a+8oJ7G5t5Ez6+3vZe8qCbs+JxMagbCCOGG+/3yPZS
xSzWyvY+inYojKf0jRYmMhFV+5k5+4nmpKY1iZTt+Z9E64kLgn294OGREUeZ22SK
gUGCmJYgGPF3tqHpPyKgMEtR8vNMOKDY3+0sqoxZDQZ4afJw7DAsW+LZAcbGbIv8
PuXHdxoCOZ9+LDIrUcJ9tvEp9vv+aka32LCo1xGzOv1wBmZokLndo6vl9wLoGIGB
T4cYdjYc5+7m1y1yhZalcAiT5df3BXQQMrm7iTHvYQli0wyk088FMtF6oEFgBqMW
7poovo/bNeB/rzwyYCkGJ6VU2D/updORLs0aGPZynh1UWdEM8/YrxcMvs10iN9jd
D0Iz5xMSmOFU+/RMqCzeF4yrZoGCB7B9PoWmnxGDfKXzG1Punk4CHwaFnVkFxhl5
B+bMexITDouUK8PXLOCZwmKpC5akmAwzAA/kLT4tPTEu6a75kbFMd9Dm2ZWsbHvs
QehCOi6tX7rJBnb87vFxyruRbA2DOLxQFji90Q5MzxmrWsUJvVQdj7WmHSY/umGh
TDjRjovNk89hn0Uf6HThuLRdLpppraqr9rx3BbLL3+6L/U82vjQfYnY3R8nuPuhq
Z/yB9bzvzGkH0d9zy0MizD++hGu0LlO+3IlxoOz0QCJzuIwL6FrVHg+ON+/aQD4f
SaehPndRjXU89YM2emOclUP3sUSc59EdoY0/hVa9KAhv7YjKLSUpaRERwynn5QOL
/5M9MGdD6276mjXlBfVV/09ZkajSQxjMjMVxB1yDPnqV/VBJZE2qXXdKVjAhvqPr
KnwA+7/Jxj8zC+M7i7A0VGfyW2YwmvCtd8u31rkMSRVQqN+Dz+nQ0Oy8IfYSfoEs
t7marf5YW++vI7xI+HbsBODJJAwNBUcQIXf/SePp2b7jZ6y2qP80GHPUVwpf3CvO
5G88/2OWYg/cjeycROFBkg5gY0+vgHImYcMHxgYIQok/Ug84P5jWY9YHbIHv5DNH
IV6wJ1/0LXBfDaPw2gkFmU3LKkzK/iw8nWy4EStZOdyh/ULJJOy/NGhuZ1brgyS3
Q6vulv/L7wkgx1wUnRdR1wFsBvUbr2UpH5j5htly4HLRa4hrG0Td9YA12xdWh7/f
+IqkJsc+n/c31XgE64uPZnXLPsxacRXfHU6tbgbkSLRx9KbjLbE9M2OuT/9tnQEO
ydCy8zDM37EZrTEGm8wem0MmW5zANEx6fPgrR9AD/ydNaDG+jErCa/Bc1KrrnNY8
l7rvsFb1/evbYLJGGabCvXdeWzzAfWxmewM8e+USVWUaHyAW4qhFHLl9IYlZ5Vrn
/SyFkyAhXlQQmsnc6Mk1c8MFO8k65Nojd7zMFC0Mhd4XhKVl+oD985IyQWhCTq/e
BlbtZ/EvyIF+JdRmwnA2tkDNJgMDPosVhzzDcBJJ8zjdyoLfUQcAvEO6Ncdp6Sy4
ZnpaoW5t98rQAmFns3qFCHag2O7xZH5H4x5RtDxTlD2C1ZQJFACZXpwkONPZh+wu
b/XQg+OFDSbLzvasQedgdRrJTtITN1Lc9UfWlk73FNkzpIuL/FOva5hlB5dLp3fo
9mjfTPGCkru5uaQvYlDanENSSzI1XiF34rdq1m3KvS2ioUKqL/70dYZN8MjuAHdg
4d+ntxTEV/PSuPVEoeb3+2KZWc/uxAjvkSqKgY+kwLhDOJbdFJVr7c3+bHi2ELxf
nfrC4eYo4lpLYOGjZTvwpBHcL60JLI9s064xmN5ferJ+eOzE4cCHcDpoTUA7SNqu
CXlESraE/MqO2bIn6WzsvTbRYj5ecubB32g+ol1WW/vlrW+ONyzU70WJMgB3ZoOh
amWkpTB/XxHda+jKm6cOe/szxSAS6698seu3nbhPLObaKTOMKA5doS0OBP5LbLrR
miEa/At1CHZ3eaewzR1FdwKTuQZ7GTx2F1P24QbLQ6eRSevkdU0AZ3ydoEJ6Vp+d
RExI0AlmzSJjSuGWjyl+IKWmuLLUZ1eUfDUCVg0ux1Ev1HRqyJNhUzvo7jXf8dLm
qPfU4jzuDxYIpHk4T4m/lpb13eoYtg4jbyxVp3V+pMM86HCAM6NcFiIEo+E/1erY
Ip/irFr1rwOUCjDIHizvpopS4RYK8JtZ1w276W4pXwZbWeEuKMmcnB5IHEIDiQ3i
JA0vZVJkjo8fJkIyMiLFHC1udplqt9+ittP7clPUNWZVan/p0qfldhWGU8cXIkih
rQjTmwigtPhVNPGBkM7RsQ7KCBg6BqjeiCPzfNoXjew5PHbbijwgw3YwkXGa/3By
KaTiqgMfkcBVpaq7GdvEVCIyj3SGfUx0tVR5+vDFTfSQ9qnysS/PVUzxpE5UR4R4
mpPolC+SMhd3vCeBzxyCRyAL/R6gdjJ54Qvw/+qaQEn+1GRjmR04B+ZKwQHlBjkY
A4pR/ByLrrM5FuO4JHRngqY4V32ixMlhwpDeWIpOegHnwwXkTdOZb5pfZ4MAJCJo
HzJj3yYsl7Xx8N5TcX4JyrK1R0/H5PVC0EfQNkHnPfhluvg+9KpNZ8QUJRLXsAQj
rHJwOYVVC7Z1grZVHshnR/JpPlMqh33zXxa0LaKH6WK1hC2FGFgzTmH7momq0XzP
RdiLL2ufPcPfzGvA7U3K86+RLF2a3LJNnN5rPdaSTequGejYouEfcpS59zC8u9vY
3EhqyCFV5d4qyWV79uX2W6+9fd3ludxgp/e8hF5pmyQdaBEJCl/b8dk9uoFFhj1m
cR8uXKo4iUN2Oh9Ur5agLETYCbGATKPd2H7g9fTOso1qVsPealoAA4vAr/xCG2jS
1kkwrXMbeb/TXHQYPquYZHby5wxIyEfy8jJwVKjaVQ5ZPUarURAzm5zH4uZuctph
R80OkxHC7N8ZENgTCzCgnUjQrvGsMwGdqvRCBVYw5bdUw6i5n10jlqTA2ozljjOc
PPLyh+0vhiQru7RkXBQDz4dmo752cM9JCfEhfc66kOyK8RlBt/sqzWt6272xRKWP
IhwibmdFNOzWVhpAIiz38OzjdAYsYG+IzKKnPJS7jkBCJ3hlLRco4+Rl0ZttgFvB
thgXTwBlAVp0qylrFRTWOKHh9cqFBPISqawkpYPqy0DAeojyeCPg6QvZhqHqzNJ7
xFSQ81Aq3VVxRoQlWrc6JS7znzTUTILqPB6EoN2jDDCAdPCEqiDoGS0D+xTugbM+
XsBLRDyLGte9ovPPxz/BkBFNAFT1vuj5zQfrg6WYkZ9qBwj38QOFdHDAKOuFoUpU
DOv6u5cr9S6O3LlMn5qKXujmoQKWuSpo90MOD1Qj06TsLVmOwnzfbQrE0dRe7ps7
gO29sNBnMW4Nlfr9wB2701vCFXJdx9sMk2hvIs50ZR6PyzcUaYDFL/w81+tkHNMG
N6cRSjgpb549ehXQW6Kt6wX5vkAMZt0ySUEH1Z8gBXuGfZmqxxg0eUzbnEa/zlEo
6cXDrr8Z4m2XkrwLIIBteszcL/6krbPxM+CzamY6lTftwHOmBP/JZZ96RtmhZpVl
Z/AHeOe/NZ7GL03GYL/4CSbup0uv68659oxJJPUAkV5WWIAaUB9Vkrt8dv6lrr2a
MI4JltEjRhbcXJeh2dHJrBxpHRVMa5jINMeg/G+scElJAxB+0bLvTDmOZDicGDq8
TIOpsw7/8SpZzeaALj3u7JCA+Gxioja/TIFXOhT8DjFE/qOcR/rMt3W4ogMIA5/6
AsvKuaiooFUllTZLh1EhPq1xM+97SXg3qb5AKXlS7smbmrCrX/DBXJLP3pGsRpcS
1tDKPmESeDBa3G3Ha6lGbQl8QDuHv7Fgx9T33bGGtkq0I795VSlJkd2inwDJkgPu
ChIXWULhhMpzIN2wW88EfFVwDYqTObFBKAiMpPtAMMCSqINnwXfEa8S33bjx+rp3
4PYOLxw6AI2G3LCVSRgXOn+7hipjlh34MJH7D5odAvWWTzqNXb601s16Y2oElf6G
7WNPArBVI97Yitg6O/QcbPB0vWqglGfc57v5xSdyuaRIWHY6NU5cLZPvoNndbizQ
HeWeJEdVpe4i0MpDrACAoCI7xDW5MmeyTTVagKJ49qjO2aY1sX88Jb14e1jzkPBh
37bJ9gPG5VIq/b9AcZu/VQhfnR39/dJt8Vbissa+X8zt4p0Kfbqgkhj1lvcKrdKc
lJjDQeZWRAV/YUdPOusS/0Q5XOYyBsteL9sj0EW/WrIjFHKosr7Xtb4OvoavNFou
oCqU3AGTBwSZTf6HJZKxOyuBj8/p9QI8u9RY5iBl+RHLKnLZuqzuIGyxECzpWFeg
lM1JbxbgxNNRlivEwh3daVgIsZcYZ98xZgbCQJDGKFOt2xPXfT/ynLkQmZ+fZJcY
hBph2h1u4hAfK9sT0OUZxXxSrrf22HMkGiciMisEklC75roXRHEvH8JCohlygBVX
PZtUiMw02kIxAsZCg70t8oiEtHO4yX/TE5sDvx60iOygz9bSzS52rA+5viaeINLv
X5sFXXLJTxZgV2xddFqIKKP/ugZgRE3C0YZdNuufDx1XLvHv3dGpI93iZu/LerI3
IPB2P0c++LTIkmTIoULtHacTPFlCrSFhAoLLEh8gy9VuV9cqmIOvUHL2+lEbs+9x
GDPwKkehDjODQtrAiIbxT1kOIDaazxw2FQd85wWJOqYXNJkiNImSAsAUhlQkLrbj
2O+XeOrgPydM5HMsqbiZe+1jjgNsT6/ZDrqiKOnqNL5FhIDCB41n9mgmawJoImqz
5AuuxCrsQKy01GvbAAvXyqWSJMh0hGRyVK+Jv+UYI2HNRwE9WPCsqVOx7PRk9DA5
tK/JFAn74ebTbAEVNYZNZr0ZoG+hNmvL/hIAPhehFMOqZrJmTtCvk5N489EhiMy3
umi2TQ109Qux0ovJWM1KgSY2MuZnX/Bd5TAPNw8Wx29uNIk7UrhpyKaAtPk/BCfx
C2jRXLXXdK15WNIcV2TlEMzXtdNmP47iHephoDMjJ1ceV5XRCrWho2x8LHlPdyZk
uon6LHCDhT2S670IsBseIqX/zv4irzi+TG1CTD+i0oZ+ijFrw+qCbB7brMp+oKt4
tvw/ktFzw+G0py8NTzDofowYtl8mcQafo8gvqvSZa3Hyw1awvML83NuP4e0i/zVo
Cg1eKaqQwWQrzvblguQA1Ge25hYa1yrx3J3oQI/V3NinjntRiTIJ7PdQKiX/Pgbs
8bAXZ++b11YBqQ3yh1slcUiQwwtPWvhYo9AbQeKuT2kUBBosIlrFmf6huEtkkiZL
oVOhqTEdQTal1dqK2mMoijagVPdmpQ3Sj6h6mdKJ4ixWOTw0iqx97ii5rAwtqoTn
rCFlB0ozNgUFfeBXsnRpjXomPJZMO65fiWVe7QrjGAHI+K8JBI09LWuNbhPk97nS
si3FSCEN3RqOEkDEwkplVF8w4T/RPTncZ+dfxygM9h5qjaFtZkJUF9atS/aaaNJc
uQ6nrHeshEymZzkdppHKSckvVCzXfbsj6ts6/wZgSjaQrQastGfKQSnpxDs2Q7Ci
9dEuz2kJErLab/dDKkJvgYBCa5Z2Z7H1wq5J/3ITeQzJspbGuzXBkpgmrxJJPRSm
Z5IM/xOH2sU5TIc3eWulKdIBT7UdLJ55OTCCOzQ0SPGj/zb/DEWLty3Mu3wII7oC
wvHEMSuSTOv7WZ5G00czqaNA+3B6ttFVpBqMFAzgKkZdvsyHykiepB3A7nh54dRz
1yw5CcNpet2Ft9PksinTTwCm91mvY+hCU0wDHtSSdU79ceFZEGaZz7DLiQPd6gCT
aiSziEPMzxA1L4DYJ8V3VQv0glX+zmj3Kza5z3dOzLqgZnccIhbmhjRugArb+ol9
0fOiD3gHRUG/ElBqEF7UmR8YQ2VYqd6GYrMfnVO5XtspFjrVxglbdhrCW8B0j9Ij
fMPTcscaG0AoZPpniZytliq7uZqsbQrJvuT7gBcQiBNP1MLV3/vmzgyZpWbfv9Cj
/sfTrkYBxJq/aAqNOYewDzOgjYbmZjq4YtpScDWVbW0EpRKCn4VMp1nJ/V1mWBDE
Pp2CQBUSDxtY8KNrct1eO6K2Gg7j2vuNnBxTvdIdN10m1z+1pxHrUbXlnuzzY1l/
ODX89Cwh/mjJs6lmuiEmJdd8SK4BEmarozuC/b4ImpIL+bqS5bl5qjBwR9uUvYfh
PjeYmD9FBe+48QofsIski6HL/Tt3lFrtKjWU9n/cGVGIKs60I5TC21sp/BThwlaQ
uNE2D47H5r09ZDth1yZWvrrObmTnrsg9VyrhB4KiaH2NRHDLQEsuWgzJCExkAI55
a6v97P0q2pe7ifMncqPAIRlKTbmiY7UPsg/K+ZVv6gBjbwkrsQgHRYOSVR8F4Xlg
tzguSKjoFkFLwyYqIsgFyVBQb3vsTrHGD9BdOokybx4hiZ9r8piJ6U0uvv00t1M2
DjdOqZTnE7PLP81TJIVu5Hv3v/2HTflpPJOXizGYxjvGnZrUDii1HG3r1NpyrF8M
CLZhqHmyyM5qOW0sujWXJqefNBkPfuoKIyPeJzuS0FF+jY1CleL/dAwxxs/gRYKf
pqyzroBEgGGFPJhUN2IDb9Gh1JD2Ok8OHXlgPpPJXRkQjsceagjttHtIH4F9q+j2
byt6JSzlDSxbxv5SuTq72bgLR/AzaqfPPCeEdim75oAXfiCL01mv7ZoHMfOtRe1q
gYU/HapYywrchYPc8YOYBv+Ui3VEkWzbMVxvuqacxqPnUbkISa1IlpQmCXMnokLK
MoivNJqtqDUjJkuzwVYxgZpm0HRvQQcVVQXBSFbHXEj/JB7Mt/2sratZKXZZm4g2
Feem2emwToXnILvtclC2vsIQFoPLM2zuY57hvkTDrR2bOXYJ7WMrQTnzPXeAUgqE
K7WFyWpq5oLjRndUg4NCACwgXjSOT8xJ0QAUTIAF4hiNEAIGE45pklSSQQz1ciKx
xMBZ4bs3NJfNIuv13aHGUita5C4sAxAlODHzPblKWoaK/xoJDZe0YoTXR9KDcp3v
4pZLAjpoe5yOw7nvczVGXW1xltMLDaCuegabRXTYIkRr2+iiKkVqTN4nSZS1mRKk
gRT8kETk08j/1m90Rt6g2Sj36heNo0nLv+GUJX1WFGM7FZFhJKqQM6BgaPYAq4FO
WsJy1o4kXssfLPtGkn0iNRdbYZjZW7qhUhxdb04zGgUc3FUI7SbtWJ335pLuy0tc
SXstBjcTFtMO7tTRt8RqeUi2gb8EK3pWU8gFcTaL3/lWY5vzLog75wLU7GkZRuJ4
Ahovg5d8JTmv3Asgwm17R4hsV+aabtMM2KHvogQkhWiaz2NOMeOr61KeckxCsDj1
XZU9hfsHZttXV7tsISch33J1laCFtYpT4tMYIgFNoz4nKk0le4ahPsDLEhr0j3IC
sbCynvs0mzVPQ/3XXSAkw3mPeScnynEGQFyWqUdGBMFjXYqFrWb1OXdvzHkoVVPo
KzQVpsVFrJJD/g/QG6YQw1wy5nUn4e/F1JVA6aLEOn87Qs6JoCClJp+wZ7Htn0A9
hHVHPy6qVkLu0h/g7iHD7uE5f1dCekD07kIu+J/XH4BT4n0FMEP4V04xFK7YPwLz
vVDAt6ypopF1KrHL5/uMhL3kOmYoN8MYBQwiSXvMJq+b95wtS2kG9WbOBh6YrBHn
c4EEvaY/FpXvJIybqMRKEH+k8pxZKsO9Khps4sBvGi+TzoE9eiIzLEamfHd/cVMX
Vc2Z8ncGmavatfKpwUkU4KRzQuwRU4ip4cb1I88kAIubXevqLGUpFWG7IdtKFenF
VL0st4Nf7OXJZ/qKb4/7WWMpRsexQ4t8djzG6NDpByFMbEL2ZMr+qpBNrG8l8ow/
/N+DQUILF8VwuvNaEwX9DoXej55t5Ugx0xFRUWLZ0zh9+loypoIHtEsjMkCZlgsd
K8it88mI1WxcCKmL8RlKvqe3nrJu/2yHY0VuiQg/T3EKI/m3ak90owfJUN0kvKh7
dKcMhHTlqepfInVzSjlt8wsEkRpcROxMbx08yU4Zwgx6ADMYAqYNWELoBw8ZGGcn
mCx8VOPZN4PvarMy/4IwTtD4G8jSsnJa9d7zkuAGVtLF6Wi02DhTIuciF5I8BRvS
Sl7OB4AafHRu6UJXMrXVIZVKXVSjsObofV9PMqmJHY5fsddAesFihb+SUBEqbfNq
MRWFPWGKhcrrNMV+ZMN9eNJM8q80s8ZI81kB89BWNG10B6yufWW1mQ/Mpjvb884s
Z84nJ04QJauhZgh/0hOcHABJvnSmzEY5HmhjZF7Ki5PcyXDRV1Idzt2VxssX3XmC
qef8+pYcybSyzsLLpxnsx6AVJqSEb1tsqkX/PAuaFfBLP8KWvfOwYeQkQu0lGLMZ
omqRJzTloagruEt1+g4BL/W1rAdWwZi/CZqeV6s9jFjCjzlSQ4U0F1Hn6Wz6SFqT
4b85YLUF72LY3qUWxeFTBKgUM7JaoFESv5n+d5NdYuoFNutJLRHZyXQeoI3zKohb
0Dk4t+ppJ+wETv+hgNwdTMsNWK++DUndAw0w0/XKP0XoBSLysUi1XO8tqJ5rSy7H
KBtTrE3+LZYKO1Unnq7pYj+r5tah6XM59OjKUcoIuX3brQlhgbrcmWmPZXBZLPFk
65XK1UghlM7/4O0tt8aNM7AdsY322eg7FX5PbJZTzxXEbbrfcpn+upDqQnJHSSBy
WjlI7GDRe/QndmW6SLZJIwZl9WKKqRK53v0IIEy1Jey8KUYjPNJACBaHOlfVstES
1zi6pQRaBRmKM2cNKF63u6hZRPAlBAZ/coCUNLw6RbWHlGFfwVU83NhOm102UjZK
EkI4gqnpphT1rkH+iKFdUMTqWCZByQtu6wzucF95pr33y7mH8ig9B4KTdpeDCWMC
ZbtcK03OYTtECb23fkYONXbZA4dxcrt060v5SV/up5btbtFvCQUlzrBvif5MO4Y7
PulaLDxP8iACQMsmxdKZfXPRNrdFUmcbk+hhqF9BaSnpxsw3NZlciVTixh9WqAv2
g3RwB46wFvDNZqOYSVmppCWwrIvfA/9Wpdubkm67K3jUE3efRrxlMjcxFrwxfJji
+1bocGvJejDcZj7hQxAojsepmL+/U3V8Hsxcl4Axlrz+dYhu83Q6+frET8ExxNnn
pZxR4dJc8EyXE0mQ6/Ly0ouk59cMd/oIldGlkz574JacD1z0YpiBvW0oEgOdHpho
Z5sUYCq7ZraePSHaeL/jRos/nAm6u7JLXpdbWpUx4hmYp7ifDrIDV97ad67JZCS0
6jfpIwuS5THbUlptwvpQ3WuEhe8PwpxS5iuV0Q6offK4jO2cWQyShKWJUH8Dd33u
vM2X4H3ccJBTvfhUmIi/DXCsF2FHrFNiQlTq52Ih9KtRT9LfRFh2Ht6pwlWNWrEZ
u4Es1UMS0vjX7vUkIzjmrVybMv4cdaP87avk6Qk9mA6y9vK8MjZYjPcUko02XYZS
rKcRAo7FsmqngSltowjnk7WT6oxDlmLid/1riJstuGotIJQkyG+n+fde9xU2NVbt
C00A3CAsgD9pG2UjpJAgMiaiXI2wcCWApeoOtb31RV9Zpw5WOwjSc2FW6YFIC2ap
Q0CGhVNZLAtNzbUfvHFo2P/xANGhTBPuYumD67/UeOr+zhjLW0Sm2mlQch0d3KT+
lf4y8/y9z4ROVhqS9vM4DKTcQ+ifWl2f1gD/vUoFMRteETHEFWCyRK3Bjv1yO+av
5Xs7GpqF7emJsEsoxz4DBo4VhonjNubLpgPisw+imozCV5rYG8yFSRMM2hWcZiYv
vV+1AKC3OT8Ppc1eYE3D1uOCqE514Dy+tM8PqLFCUJcfaqdoJ5u3LxgAwXfKIJg+
xd4Alpmh7vUkwfi2NYCxhwqcrVOdNuUI6Pojh2fC85IR+Mfxjb+ZCJxtzfq9xOyw
ZgMAFwk75+rzGnkcPXDolLA5PiF7I3uaOzavqYNeMECynohOo2injOBLnpsRy1ZD
W5fr8PBuVCV+7dBen3mxr5ClmNlGkMkr5+vniScM+avFerAlpoiCETh4W+hXlDUi
AqfcctBBtZBSTuaHULLBqrehkwE3d+MGUid/QWAr6YseQz1etSX9lWV9jcDNP39k
CDY/Pyug3ijHGgEtKw9vWvkX+GQ/yuVrgwTp//7axs9rkPDG3DAPIqxNC1I2YNuU
3h/hmERDcOGr59TcUql1q0RaGLRCs1NcMgGebmJ+0pToLCoVvQ0a6icSv8uL6bE7
EhnaLBKa+mEE8Xp6mSXGDNyzHMg1mNJ4Cdm2KkaaTxQFY6m6HUoh9oOAbL757eaR
w4gAneHxWsFHVIvhnd5n5rvNRgIovXPKEkzAgFBC6SHixXm9m7s/2KgcCzBr7ZPo
2BsBwYIzJNhDJUGSMYoOp4eCm0gB85w+HzFqrT1mgi3R1C4ZcK5lwhGTfl+hHCGA
drAAmNv9+FzyxgH2mZCMFkwug7rs1u0SuznbbrA3nLNROOfJJMYzY+nvDQPVzYJq
JLvvJqxoyQdeR+l+xgR9/MKuZrFP+X6FM03OFPuw65jZhWJQwkKJW/PxrDgWzqQ2
Aoj600kAsvOtI2hvWvVH0aatY3BaAyuQ/5cIVRwdbB/Nbjqauumk9Raazwr8TBVB
Mo6JEnB5wn5EWKPz4H/n71WZhA8H8oIcyqLhMOqJVg3cHlw1Rpn3HQHtxEvm+gh+
wX/AQy/AQrL2E6piYh5RBQq1zfaluzHe/pvedqQ42iZoG2gpfmhpmj7XsL5IOTIS
2vT9Q9MGnV1DGc0tw95gjlp6AKk3gQ4Zq9q3hfKZrKYm7iZGoDnHyc8K4G/RQpX3
Mt65Y/wKIGtWtEFzwKZPd7rOUFf/QgQ73fs0mwV6zjfBWb+IsaJyG9eTCGBUr9dV
QD1XxR8JCXWdOM9KGohaU6aeHM4tzXL96ivwr+iiCX/Lv+Uk98OanAN5Uy63B9/E
RS1vZ+j6dxTUUYW1zRqlQr2xsPTelIri7Et0YptX+ZHoqv0Et0Y6D8Jl36iHmHkT
IvEBy5OlHQ602Q0L/ZAai8UwrgBbgB5e1sHVpV2rYpT2HSBE4ifNL7TjqvNOKVEh
E3a7Xr5NBszadP+u25khSbTq1R6+qisR22e2nc3/yrjie2yoDp2mPxsMjFdo2AMm
S0dYK5+zLqlGqeCwlkmDo81TQT1mugiPmUbR+nTjr2MuniLmeun3uw9XpCK0MR2h
OkCW2EZVPr3y7dcuNAfcbKIRFXvx7vxsx0AeakesiMZCmjAiQYdVwmjqB8fMzAkW
m56GkxC0uHVdC3BkR4hOA0CP+KphMbKqdvT4hh+m/7O3qjvZ/rAKK46UehHCaQt/
QPUb9kt7gRXfN2VVnl3HCKCKTVbLcUdNEwNf3z6EVlI2uZovDDlLk0cW53Ee12V+
MzElQ+ASz1ytreOiJRtSSXdW11xCIeaJgymobbkq20IwGTV0v8GxTHhQJtNjJjYM
hIKbM0DmXPBl//ehXKtyR4l9u20wrFjjPCjhFmIi4TggGb2OGkKtf7A0AyqLdrZS
DIXPhpoqvR8qsUqyAldKdOqlPO4W/uyOxIQap20u6FAdIhNFmBYD+ULXe0x7jsku
Nf3ZUQ02vRThGwA/Fcdr1aVglNvLYdHJ+XWnsrXiScD0xyS2UOCAHdCDgaYsoTlk
P0g2pPgnNMxqelbKzRtHxw3BRPDClcz5yBfFTaXeHPcyENIzHyPqIsrh2hjwJBOW
lb9HvCJMIUc/pSepsvbnVghztGlGSnY6yaUfqyJwhw8fP1iE+atJXFiIvikZ2EV3
o9KEQxZ6Ipq7WcXRBvTjyY7pq/pCbrA9T+PPyHTPrOUwP7rgd1cdt+wLq2Fr6VAd
HltjxtBZ6Z7TgLFdtbuFG84qAaqtvmZndCaO7HF088SiHpH5mTGevLeZC36fN75y
6gfWQRcD4HCkr0x8FpwUugQF2UYrZoQmAxaEswqnpZLAU38/rWzaVGXIhXvixWVn
mpawo/4fRSRnd7ycebTxbPgPGEb3C6De7bfRPmNwFXRt4vMEtwl/vXQ0OfWwNW5j
JJg1ZY9aX3Q+tMIu2B+Lyk3PjC9NC3QMfA7T6PQIGO4YdNHG8XyKZ7XHaXgx+ho2
iwXHS94/aEpdOo4TTLSlyVnFsRCtWQd1mw9nbW+cPQ/fd16NBV2jF4K3wpo0LujU
sFeKXEITE4PIoZ7hWjaG87OQf5MhmRUTfQCiF561aM59zWFHrcwEPU8L/8pZlb/T
aeBrL7Kuv+EhP/CIAGqculQTwXO/2EzoZYNYUYpTq2uor777x6bPIaspX6arPwlz
sQZQnZzFIWYsDfK6IEri67zWsitg5evJuDW266TyY6ntNc+KW/4Q9L9L4PNGsxrW
3KlsTmhyhX0zFn5zfi+m7ulA5pXLMlkg/gK4k6reIY5ZrbDD6tbCNbV8k3cMOGSp
shFAGSOlx7ezOQfVIY8buXIXy+p4QE41aU1M9MXEyyvFDo1+WsL1L88RDo85vEJm
CVF5Yk1U8MRRrdLd8+mSeFeMv/9+SYG2jf99Z63QKE2KCSBCbY36g0K0kEkuvEGp
HTBf2MVqffP4JoMKMksx076Tdo4rTIboetnwBXbLSs8ag1uzqVpBEYsv7v4DKil2
D4gsEbC/x1hxIlI6mu+On9eqGaM/2tEjGvZU6vrgoRHUy367dEoOMI0j6KRlHSEE
/MSHKyqWwP8f3zUXEjAHamCaCjqhBDQUPogiXXdB/wjZIGStLselFfnz1m6/HP41
b5xNo/2SxTUMsKTSw5ojA3QJJaAXd7+OOI/awP7OjwLoENCghjILoy8SqwgRBbpW
+Q5p23loBIGOkhQ26hojMlvxcvG3VvEwPXrgQp8LurcNdQCTkz5FEuYSNHToJu07
B3pjhbiXQR8+xwQkDS3PywJ7Qtdt1Q+8WnsHTXXqyDSwmUPj8A+UUM2SHR9fcyI1
pM+oQMEB9JI8tZ308evdPu2/5r0tP34BnORUSon1jcv8N4w5T1jzQF10GI3DP481
xfRz6uu74NxAOchYZZBsqwS19ud8LcaXjkuVf/PAhHH0zPYGtwPZ3z4nGMpUST5S
nwhoUDsQFHXNWaN92ukuExTx78XbAkCqTIvsLHlFmmsNKvxgjfZfTOC0UraXAZXn
XukflUL35p/ZQL5WEvE7y47t4hsiK11/wn9rfIHvHJoixrfKcn+68viZx7YW45fv
hjQgQ/D/CB7F7fVnP8dLYUCaCM430cE2Q7OVJOoknblpP3EBq938UENOcgOtKJxN
3//VjuqgV2NFeudyjZiZY3Ldjxm/ZshRIiKMzE9PlvNUH4Yvk9nmU8v81r2MOSDR
w5hcP086eWEmONJ3Hov+qTH/KzJB5l5WJKxXor+DhdK15pRcQ2VdhscYfqGXMIox
JBNKQL95ndPALPeE336rjPrntazKkPKihT+g3leJ4knBE3NvRiaw4ggFKWkW6Alz
yel3O4+UamqCuEFcYBbP2B1nDynKXc0GvErBpjohNJpVdFoRdb7wG4L/EKiTsx7E
Mq308E3G8HgqlNMj7sh3+MqTO3qYYoxAz3QV1ICW8q5LrUjSbSg5gP+bWNUnptBa
Dajiv7rU1GX6BEnWi8OFDoKMC22dEzM+6AMZOpc/G5RPsXSM5BMk1cBsJpoI1qc/
czV1ZIJFu4kkbWXRNjOxbvaA4L0zJMBuRwwMlpS7MsVd3RMpervGgKGgh4OaDDda
R9ILF8iCqF1hII29I8iRXuEK40pm5kOor645Z+wDpT3tyUBz0JVaBHkUKMmqyWXG
qCPzK+csB0fPNvvDJy/Yx5/HH+dgJi9F0XEAIkCXQy3qQuPjcvRewEZgxF4j0in/
F3iUzh9xaLt5ELMBE0lxM2lMVb7b7vIlQRHpqIoHqdJDSCI2l09ta0iLsZfz0xOa
hUhEMdsoyibPoaON1dJWpP3LWJj7KzjtUgWjUdVbhN+7xoBF82ykEDWeAnwkqwHD
EvzcDspRrUPKJisjqiRKyIWVoShIlGkxAmVyAGVwxM5fgh6i/Igk9peNDgcRx+HQ
67Ni+JykrvYskaHl0fEro40jEAF8H6UBB7x/Z40W9/6V+qIj1gjVD+LyrGDwkiTD
P08yzG1HeWCITZr7TCDlEXhkL/Eej+dfh+zrQrS9xf7c5+LWn+RcOoJN43RXXTNR
X+EXPT3UasBGMLwaK7MhIm84lq4Op96Xl2Dn4L6blbzNPwm5vr8olIRZqhhX/lAy
/1jEiK5a5PpaxsECBRe6ecg6bUZclS7PqPKfBW9G0UtE1sHRaptxW/sNIPUMKBQq
XThioxv9x5VvGRv8greuJ1mAODcrSAhwAJAHE29mFWbGtiUouwB/qtA+BX9wUpwV
TW4kzGLNLlZxfvc/B02RwRftzh5iapW/hXDGChajWiwZoV20SNrmk2uZ5cqIZxEe
fkTvA7Eszf+oU5hVZ2SGNvysnerm9GkPpG5x3R6KbhDbxrUQY0DxpJOX3RE7SCpX
fHhtliWUS7nRksQQmES7EgcpJ5ld/X1VIx9gIMjR6Fk+4NLyLwpkIjYamzQIOTez
ABGG5p/zHJE0/nMiOv7s/d7TOoHyI1jmiIVZY/Z0x1DC2F8//IYsHm28SK544Txe
TDWssXdUSWGmXdnketzyWWZfChGOulbiIlMBOKu+Ji4SJh8QT3chZx8vpo6ooQHk
VlvdjaBhJx2M7c7kDUS7e+LnaWZ6TrcjBLC9XVxlNX/aAAQHxDl39Ow93XsZrVyw
pG7wC7h2rovpskp4mreExgeUZrl+TquyEGSk8pITo12VzeuN9MmU/jZCif+IY1DG
moeQ8QsmhjIPAcyYS+7Ynb542PA5MYC+3zaL+p+T2+hVwIGpSV9RJ2e1oMmTHNcM
/CKbu+rRQ3Tsl6We5O0CwSaNaiwENfydCDhf1LMB9uth0bfou6tV0+CB8oS40sN9
MBKNh2dfMKCUPQjAoF004W0jZxalHcpj5NvsIhFStN9djHabcQUgM/v2HgLn+TUK
8u4Q6Va7pCj6uz9hMkk9z//ZEK5SrnLtxa9knpfT/nGV2NfzR9G0PQtLL5gnL1wS
yMm1V4PDHOyrUnnHb+Zt8U0GdkquKTeeEGyDw62MyVCP+YR1pgN4Z77+CFQVf+an
aEfrXdxuVlXnt5/YjiIryAPUz1Fd1f3q/J7QRTbo65UtXfV7k/L68cd2DpyC1y9/
e/QAe2LcusHTB037KvzqwTxoj5eIGTYtGnHjDfzXo+M3dfXXBVe2IGzD7mda8iJ8
dd3mVfU1el9TkV+dD12cnmhQb3lT9fBpneYqWv6gcrJdDarfn26DeD24QTotU1F8
GF+blQPZvnLMpYyeK1yIHKeEhxChX71TjM8djhbau/OFosa2XN/QZ+AR4tCy/ZE4
Xwk5eXW7Z/Ev2Hgfg0zaXp+kI4Q9xlQPQ9MvE109mDh/zew6C+G5Y3t4UKpb2WdC
sQpSPmPN42h86tdy6fIvs5Q91yGlymziNfXLcljYJB+SgacuJldtbUdvy9DtxTRF
LgSOxZtGj2TojBQU4wazjhj0Qlub/CTzdZU5HdTq05SR3128xPS5QIoM0ZUVEceE
Ul42cHA/1itoJJJXdOMYZuLUUH/hqMKJjJRLv6IO9/GLrExpB+quOIJloqzYavtK
CkGSYAjKQ4TwnKUNUQgrtvz7Gdw/nZIpdZpZ/b77mZUEm/fma51M+QNnLzJ03wOj
zf2DNkv0dW3fiXmAD8RMFjwBbzWZjbW6/IZ7nXSAHXHuY4wMOQ3UiK3RlAPkChP7
P9uda7v+e7qow5Lwac5LSP2Jucq00O8obWdwjuOGjYsLFZA3AUKz1QUBKvYKIsoW
r4XQQHWuSoArWbGhtGweOvdjPxNeYFkL225Q6WmQKsH+W2JJNLHMj0SPeJUiWl/N
9q3dXAQ8pp1CpAachnkE+ZjC6cXXWQLYbM3krFzvQshhp4DnI21NfPhX0h3xp3N6
O9inXCr4aBbsztaAFQ5EWFjuv0FnZvvyiuaMWUqlO2wzXOV3OpbNULoZeSSvh5kv
3J/lYHfZ5HOfj9zqJ+0npxqzALYP9wAyHZNblxD8iVV65uuRce8fxfpGkaHwGMnu
n5aXGNT3i4bIQWYlTQFUDYUGEghAq2pw5v32NzhnWsU3VwF8k77rA16ZyeYWQ4X0
Rd6d+/ylb1XwQIG4za4/sHhGrUJdFwp7C9lb7wdVZr5tQDVqORy13H3VGKXCOqLp
1A6DexbHCisHe7FI4S0irRxqRqkOVRcTBxkg88Efmk2hxkigsAJChfMELeQA/xq9
f43A2AvqVXFU07xEKARApZnQC7Ki4F6jXkXKlAWndlfVP54TL4dC4iOW3neCYCNi
wrfyon+wPVWyO6UeuQ6VUguri3i+rzE8MmK2FTzzdhBGoZYEqSVPiCCjxwOKyEAi
iLUg3obZm3OisMHp6ZW47fvOVe5RxH/eLWa+tTxQOUH5GXFFWlgTttKxZRn3H9/P
NMMWV++i382pbj2DIoVpidMe1sgh839XPG+rtOxosrIqEyuvrL7icHG3WVghv/DX
FHH24E+9hy+fp6IBocUzw8uz7wwH6rXmRoaHIKdrXPrsmFjnB+qZeoblraV5A4Pw
eAveo3iR/ySIrOVl3b0NQt5/ri9Qm5F8kz2WjMrdNTR3550bYjNcQ6bW7/Jaqt0d
bRO78n+df3xwRD6LVz6uQ2yG1KE5azoFIYTb9fZpmzSvFOue+1qtyFLPPJ549n0g
KTVPzvroCJ0Ff4VQjmKASctALRndZC1weQPAMu1sJf7/f/ARy0zT91bGltU5v44S
LC5yXsPgPCZJTjHuCRmCTQxq8fFElozWfNgLMj/Qw2KwVpRgidT7YuiE0+L7C+Ld
zfYjadxWyLKkTAdpa0yEpy8aNTy+/rQ1wEPp1tQ6IwIKoZ73r18N4RjUPNC+92DP
24OieYDun5Mv34w1yAx0ApZnZxHITMLjYlPphv78I3dbEkR6BAkor+jNseS0JSs8
JvChFOhEpmtFOkbKLGtriZIEhpQCNHFISYjW7TKkFHBe7pM2sysstvvPjJDWyL0L
r2hE8hsEMgCfEmX0cmdJRCb6XjUxxzj0aGx6ez0J20txHap1ymPFkc7kIQwwvy8p
UZuNljcNx4mH2fSkdlZcb7akI7ZxdyLBC339mksyU0kcKlRhfWgnznpuZQSFyf/+
HHvGkanRxhyriQv9cQMx/h5b+rtnsQvlVnf3Jmyr0QP4hOZbtqwIOgUNPXklUF/2
5AVELQPCUcXPp7k6c5viKn9zKFXvxkWmlIrBMF3XKk4bMZKDE6cxXytXPuONB3Xj
+LNbXuwzVoJp9SBNH2hAxU/F4zar9v+nHikQeiwPf17H9TzyyGnrl/0WqE/z34vD
lVwSpIUQ2wxe8+mYrSbtnRD7bmNUXanvxfG8viDwDGnmqMDA8Sj44HvGJkF+KS/0
rzXLhQoLtMeIcjHfET+zUd+woHgJVcxWuqzcLMYQoi7BQcP6pVLdPC4T6L+m6KO3
74JECnnFFaCawXBNO3d5jd5rPJb8RblvJ5ZRjN1c9mqzRizAjwG6fW8i9hnrfBTt
q6mb11idiubYBvF0rqwQo8tRjcI+JrzOcN6bv7vNTnRwdnSzETaQwWDy1e4LLlIh
iUIIEtlIOwIZ8N9rO6+AOajJ9GqXVu2pBPSGGkBC7PH6StGV1M1HL0MlIlS4TXZH
9zB633DWO/or9BHPo2hD63QJib5wdb3jnknMszv/jNJSWAegGP8J3oWM0r3FtGV7
gJSMgRSWGMyEFPJYrYapblpr2DSVJLv23TiJkJVo48g5uywW7g+LVzAsAs6dYikg
/dFuXbHw5diyBf6w2941hDlD27gRWddyba1WAn2dxOfKF7xat9IHbCmiSqwDQbnB
FLSjiJUUlPWkmU1ajUPKSntykpgR9dWSzxtjaUi7wGGSHoDutPmowH8TezxgHBKx
wNaj+u35rwLw+IIjn/YPeKSx2ZQ8ltUIjuc0f1bIT0PJyJbz3lr03xuxv74irVCy
GJ9HqIoWgoO3DlzIkTdKjsbaln8xjeqyfQ/GACeF9N4xEi6Fi02yUMIb5F9bh3qZ
mxLP+801L3uvjVwOHN/CpdANNzgwiCuFYVm+LgqOhZeWzbu6X6Y5pzkSpqi+6X7C
TeoeJEocnv4eTdtrNaDstEKtpOE0Egghu9flnTUiiLTT2d8Hnx9Mgo+3YmM8LERx
3zOTgdjdbUcGn+DuEVkCg6IM2g7cLoNCaF/0Uht3DBOqyy0PYHs8sPhekoCxGCaE
9sbret7YQE7UwSbAwvEM5hDFa8iOAK+eW+iFnM+qspNzdX+i38GHs19aSnsRDSyf
7WuyE1cHpfgAbAaebSLIdSyam6cjsiHjt/ThneLm4tSxoYrc0kA0ZrLA6VQaqB3i
+o9wOTzuatLT7YaL9wfykppVMOTf7hjgo2PkkjrkmmDP29yaS3w2drufE3jA+Sl6
9gwBsQAMaLumdqk1V5aanuDWGqBVg8oemniuW/RzQrC21lGdify4QE89v1JJHh7w
DUg2P+tXYqnEXe0zFvJ/mSgkyw8yWUixTvlnXSxQt2z5+6aq9qSHq3ykbaJ8Doaq
STZ+TcZX5yx64UaWU2/a5LtQuKML8xb+HXMwckflwhXc++pq+d8A6twV4DugeFov
JWB0bUeRdqJ84AOnkxyRiSuwCQiKi75i9FP9oDyCVargy5VcDkD+69koPmZGUVYH
Uizgnuo/FNxlCQsemHRIKkLUGbYv1xcbq4KAfdn70eFlzlsM4xtufx0ci31tKR2M
UPRCRySZbPZk6ssS6+rLISU07RTVDL+R7RaZaucPZQRKSswXQLAValucL5eOXWzs
rV31T8RvfjollTm9TdzrFAOAOgGDjU8+ABnnvNt92z7STuO8YO803t03IO4hw8Ae
HW28T2XvUpKLngWHbdETyxzAoyS1P9guz3x8IIH606bl0xiwJLKc77OBKFOd5g/1
EguuNtJ5z5w/obYDFEhCxMQE7YUtRPadezvQCqTATOQBNPJVZ2CnenChQV6/j1S6
+X4zpenvywmBuM8Qeem4phONQLGsNnpZmdjwOnJdZektPjpctIblE1IDGRWHUnIK
bpaMwjC85NyRrpKcbaPpeUxmK8p3D4LyHsVzR35IyauA2thw39xguGW1hWowSsWo
RPOkCnK+Uaf4Gx8oQWM9AS4BUfcg22+VQ9KLs5W3C3WXo5Y1lGG5dGRR7OiPnUL5
nXf7JQITV2nfTnuLVGPVGLxcL9ygNYLAoIbadVCKiIBo8+Tn9UIRphnOocv8XVCt
sflC9B7uEZl2ZZqxNzZ1sXC7++biasYkJmbdPVeLV9lZhb2shXIfsyPfGLfjCPaJ
4oq9lczp0Ccch2AURF+2grsUW0KTTQ6MTlYce2PD0L3ikNw32Qs3urGSo2qexBws
31goyleJCvl5JC9e5AR5uPu3hIIfdYml4llXf4t+ct+bWzao2OXlaLAYOD3wl2tJ
Zxc3btCjjN5iul8nIyzqSkCezJbUCtd1is56DTN8LKdCGFCFkmbZ723cpJ9J9/J+
1s+3PiMg07tIYI2CSy1501g8zM9DUz0cqC0298qfPsmdkg9xqNc68xH1YZSVFwm0
vL/qMJFsiqdtTcJV0sUaMQU2cnNxh2gc0TxP6Sla/rzsQWIkOJ8aGGo1ED5isDuB
gYz7+s5zul9+jMSfpJEHEI0N0cX+89cS/5xihiT6pWQnLax5lL/zeKo+Sl/BJLtz
A/4aNALPptdCw2qUeIAyx5HI40goyMaBueWE9wLyqfAiWjwktK1EfP7pJAKvBojp
0DMNfZG6+JBOljSIt0XjqRrI/+mbj4Q8xoD8bBptPB/BnF36TJJpzvAaokQQyWR1
wHOhfKejZAUR5XE+whkjBEQk13yLJeeDcS9QTZS8hY08HYOUD4p83/2srO78zDgz
ibregfwPoY/ovhnD/rVwyGAHgd6qfiowBiyEbY7iLhn2aMfSq7kNYtuzE0hIf1E/
OkuamfgJrPiBcacjF7XbJEmeGdtGgEjGK/2Npf3dtrzJwPm7SQhEHQL2u17ZKMZt
I7FHu2dYqzmP4YxoITzxvKQ1a5GLG3u8kjJ4OnwoxnctwmLiVkdyQtHd7KXP0Sch
SC4oFF6lhqZLr5cGKeiEbS1G8Jaa1n0TDEbTB2s0Jifmx20RJRBruWOEfjM/aeHM
BCoNk5VQDelJzH7x12IpRvXxRIHj45goxmTItXFvSym8XaCMMpVY+sJXwspDMeYa
62te5SlhCWuB3fEcCaBxJ59/b3vfyxvuNkLFGmx+0lrvWUhEYtlXSDjexh7vuvd+
4bLH+eDwpUYhHxlbs0LuFiNo3OvjXF3m6fJ1EREkssj36q8b95ah9UW9hc3DokbX
MbO0UwSCWgLoMb72o8TXXyF796w3FvmnQMD4tnvCKDDeLjmoUFNNUflwbLYHfUcv
fXs0WqucJX84/LuTOSEvwqTxc5AjOEx1pP39HemHfd4h36rvBiUQ8fXoFJnFvsKl
e4s2J9+egEfBnKvq4zryzbeSN4RpTGeBO0KUT8CakM2UfPujHxlU5ZxJPNn4VKHN
wmzbFOfhjFAD6Ch0aZDCfpKwm4CoCdfj2XCe7okk3b1WcY091rLMaS16j9leI131
Ahf7HWhGptgAWDB1mvZLvq/O/46IibSPk4P6WQ211BVfkGNNHxZRYPEVjlmi66mK
5PF8eBbrRMhtgPmsiv3YZrnqXyQPXeqNBjmvwRwlspEEvFOyX57g1dpbjN4xtMxU
g6YAC/A/tlk0YMFkpsB1N9Q2oD793ZPCrYxBxGzq7EDLQUcj6UNinWKoK11MG40o
CHSaUOX7RDpiGoGgDOHVMmiVbDDatu+nYWktLg5SHQfUWuYeohXqn3otwMnL0q9E
MoSjd6AQGSGzcmP/hd05QdkwCoqVI6eS5Nbu4Z86L7amqGY/qvSrpqsXbG/If+63
DA1Px6RIAvVuqQmEUzYLZAG5U0Pojc0+mMTN9QQUOfVl3soeE9Oy1vFdXGSmXkrg
JyE+Vi+fO30pZcrAXXdoEZLF45bXGXi8xlYOWj1CKtcfDWFokPDfmLvSKUJBdEpI
0eBmqVTsvO38+65jdFLxwQo5PqHvMARCQWKMPQdmeQCFOPgSIJoLQoCtQzKb2SIU
22hMY21SKp+A32I1QiD2d6yEv3mEk71Qzb2ULSyZED+WcyrzIbUVrd3ilBG04SD3
7PHcWXdSeIAL0qMPDweDjdWZZWahFFa9KGjcQP1KR0AdQRK9nxC/osEQhdmpUzJP
ek3mn4+RdnJ6A1clCqdVqbl3NMIded5yfSfR8qzaoZEOpkZRnZtpNW7nHADY9b/2
G4ywfmKggRHD5O1F/O0Z0bXaByPiMSEryqPVHb0KqQ6RZhbwRAFL+jsWEwfcbT6u
MFYVaPei/3fN7Hv2BH4hC7ndGO01cMMbKGAxmK2n4SAMdG0Ssuq6JKOxO6Bq2tSD
CmvLiq/SVxPUwm4xfLPSOxJIabAN8QF1yKJ44040l3QoSiOaACSr+U+5BaMnydOj
/w24ya5keLDAr1+Ku3Ay7otC1x6irLWdio3oCDB1JZB2MDf088Lt5iXjXldeGo9S
lTl6fMxNejk3Ew9//z0hxfHEvv17ERgG8JyQN2B8UoEw2O0rnVxOB9lS/aYe49YB
cpCUgiAJeTkrX6LSMryzkTz3LJr6+i32rCIiM/tmBEZRnhEcKk4c60HpDgCryGsP
loM2VvU9uG9dYgvVLsU8QDy4IHkFipiXO3SZNoLWHksTfRT/pcFVifcG0Lr0CaN0
c6Z5Yt1rnqSSMLf+kqMUK3kkOA6Z+CyPArth/5SnfLXLbcGFhmmpS3nYR4/g+UAS
QnOtPjZ6YBOVyWxL2N/Vf20V4dSDZGSch4Q8Xr+iGVFX6uBwIAPSCePES1RPEKH9
3QyqF76YGQdV1mx6TSRyK/XSmrdTz7xmIdX5HdaX/Pk25I8pt8ZuEuV5su+YVkqu
FBBpDbqnimSLP3dVC1himmlA/aPO6CSOqCEVGryWunRHmmwLRlw73b/CDX7h5X75
tKTr5M1pxvASTcst9BnOcfdgFKsN6ThNfus08GZyToqEGa7Z53uysRrEK+dvK4kO
7jWzlEvYUC0e7wKi0GQv2j2p+0XEVgwy475BSOE2C45FKf9yPN2DDfBqeK0WTiGK
X/UOXUEaDLxGhNWmgaboDFAu0p8nkAHjOsjEN1imOcligE+v3QZzoSXaxs0UgQyn
L1EkFQQ6IdegV3w9ceOoXsCUaT5H9ukoAnpgj1E7eOwVSyF7XZ4Hn4qdsQNzwqfL
FcIUIlODW4QzL3SFKOvCsSH8uTv1C2cq0FPw9w+iG16CBtgmf+fQJl4EaRR7BKk+
q4E8tZawH4GMfYKHcxSBi2HzxZsdytxLx8bO5HytlgdyvTESmReaj+Nr9JoUstS/
aPM8r9rw+C53RUB0szD72NotgKqm8v/GKCBZPXJ8aF9uSlaM8zysYuv4vNvSxX/H
cL469cnQzhHP2LYc36WbkPWPpXH8afaU15WywbVIRftp2FC53KVdGWAbPAOEWoGX
CO+AUcdYUsyRE+4WNrrlOlIRK6FgDmfMSX62Wyvn4c+UZWfYCWnxBsTIAIMLV5mJ
x4y6dN5/jNjzItTkfnZgMwewtb3OT+T7gg+vk1WCMiWgVF+u0IM5Kr/PmuGmhPw7
9HEbRXWzZxLEOEIyBtvQgp87Mpy+iCRuXHA1J/17wHhTe05Bbh1YiC+/kARHE9d0
D56OgJkNhJouY0bGs3+Kn96TzrVUKgAaWAwSfG61c0o1l4BY3BFlTYUVxeoOKWOr
T/RSjrmrwfupXaRW3Lb/yIuWBc6ew1CvZvO2p1ZQx3JMCkQGPZFuKDcT8cm3WrwG
W03q4bJDsFm/JrrhSYJfx5hAZlUh0DRbdqTh/qPP7KPh1gg9SNsGrYIevoVb/GsV
6zG+/h4eS6Rix/l+2AVVvH8JeelrNSuYUlmc+tEsggpp3fKoTkz0P4tk6wj9xBQa
53JzuI4pBw3x2RmLd/EoXpKXQdozY1dRd/rUP9UQKIgucWnhWIT6PnjXbgEkRBAm
5zEDMEqgdxKSZ4YR4MucuxqV7G1NU1uew4SHfIO9vF1QCn+dYKanj9zxgb+k+7/X
ctLiCGA+yVOXx5vbkIOlGLEidhsFDl5wbQVF8U5pNK56V5bIb5NnzCtMWS0m+rA1
/Bque+2BCREtwvLsSUWn17FJ0yG0aTy7ng1NlBVZ2w2l1ZHy2VKR2SJLVSnyp0Od
FHdyXwfNLpD6Llc/kdbG3RjxyOMPvhrAXT44LU7vXTZn/GJCcAXay/A9okLmLYwJ
MJiglZYK2/fWTxPoHbB5ED7QInqHl8PU1MO8xFrjexvt04PphN5+L6Ehp1Rfr59d
KxIysd5aUSFtZ18hn4IkUlFqIDHPXLNfBlN8OQfM0W3ZTj8RlhzvQz0kKf5V3ogc
IGhPFT2uCkNeD8qwCFUJNddj3U6mZOUtJJ4byNlKM84CcqVqUzVTraMNqh+4yg6J
KoSoCtBFtt8c1/5sEWmqrUlRU0pJnaOTEyTqoR4rQPEULimLCVqWW7lRWk9lyhDt
sWszrKL5ZY5QkfJCy2RYshtxCHsmXm3zUABuuL/Nb/6gI8oAUqAX0ADj7SRbDySN
ZaFXGH1aJklkcmH5VWr6iOFfO1lSGrvYGsKaF9YPL4fcriIACZI4PieUxx8wJOIS
xs+KVBSlt4AHxjY4S+3CWir02LX5GmnZRf3e+JagPjmw66bABTEaw/OmijXZ5QPx
ioB6hpxlUQlCU0M2jacb307I6ZqHD/wJz2N9ebmDBlWMiwvFj/YGutuVun52Td6C
9zaoIB7SD5Bjp8Qyn5l04TyMeXiwNcKFTz3HsgsFJTywtcVkxh0bK0GGxFnIBiZQ
kKbZ52l7xuWPBI9cVdxmOJl5/OWex62TNVVibBJGC229E6xhj5aFGqbAFZir1iKi
RPOGiL6nq3WpAgtiCgZnFtjZiUnfZhD84Dp9ogBGQpWwmTjlLBvpPWYdBqE6Mj9J
EcBS51p8iX0rA2J3Muzva8or8Ow56RWDhVqRkXcOp+eYH+UGxXIz0ra7JQlrsZiA
lr7f5OwA65L1Mjygl0MjrjZQolrdj/0/FH2IpqvaWXWBzBCvOr72VO143+Xql+rZ
YLIMR0ixKljWEd4NEaHulSm2Rzc2LienMDwu6Pu8FAf2p4YVgxVCFRaTV2Z6QdoI
KUkApZsmxzlcxPDdWNQQe9eD9QM/pSpZFtkfc1zMtby1gBHP9wVmIfTXCcikWnsN
TMiHoWIMWb8Z4fSt/+2UKOUV7HK3PWVM8VKMSohoZuTVSgF2Lryi7JFXesC23ZwU
y4qDy1581dKo9gb0I5wSI0qv9mGpe+a6OunTPUQNRmWnxfjXIcSeXhhmAs1fEPMq
wKW+Q+b7gHfDCznBoKJu0+c/tkEdd5L/j4Usi3LQYUeZZJ2uTyWlFBQA3Zi4dF2f
J/Jwp2e55CKTXzXhldbY147jMc9dvTZwTssUzDzZ5oYaRdEqWv0ECjx9WQ6Gql1N
3kbrYjABT7kVf+c//EVCrGNfXtOGBll5eCcjH7VrbDIu8KEflGcET73wLq8DDqHU
lgyGejyZPav4NjwTen2SnvNbosTlXHfqWDWQ/R/3YPY+eXBKyC7XFGGSaALRLyN1
AY4Q7/giiUMZnIuiUQIUNHK8iZRjebiYURW1SaKpy6yh9QYi6jU09iVZLKvdgXBq
xHVR+34e9mq8HLoOoBFHbxwV5OfNl/HoYpIBU6w1IjYi72Y1MSuOU3EXjyFUsqBH
o6iFlvhFWtpvO1LvP2TErVXImCb1uT8dInyDolH2U9jHCWqZiw6LOrPTIailL1vq
+z530Lmibpgl551CmaYE5qXDpqEjqZJwBIV5ibbxB8d2bPuYbiooAmcu3ojjqdSf
w0NasBynjrQZchOmI3QxSrLX2Jfq/IyGXwCm/Fshb2SvN27RaxXnaft1K1wpgurz
vQR3HpxfVjEP81qikWvZWdd+1vVTSyfGr0R+I0RZzbIAdM5Y8fzAn8LvFCFfbna4
fjM1Le3C4YL6ETeaDcdJX9uyqMQg1QU01c7zoaiWXyyzuWWwYtR3uouL2CM5qznd
whwCd2ivpmVxJm3ZRrLIk/Sm5NnUueiSU7NGENvnJ0pmN3aKWX0vUNzrUmPOMWmN
Gw95OBMPYZDJdYurzktpLnUkrGtSMC9bofQnubP6QJKTvawjebzYeclXoj7/9KB9
8EuG8MKfGPJvXgwDU0cqHkBS5FM2HiqitwSVyQvBmAiY0ug+eEOkuBwxvc5Xf5uO
kjXCn1XlLY+AZA+0zHA0ABexR0PzRBGDvVDoxHEXSkzW7nSx/+RgKbqlcrr9Zr3u
m7jehXJnuW2PBlYnsV2Md5j271yP5YN4E4TNKFxrm1uzA/oyzzOpj76n5iCTBGXC
K8sFc0x/X5ABQ4pEyAOB6jnKZhM29ddhqIZMvQTvyUdcJZb8+62iFVN4+pmw8wnL
s0QI3mVd6c92GZvnFdfIYwwIvWnCqWM2zOBaI4ORiwW9laCqRuAo9r6c9guMJrGn
tpbBsKssBnERlUhacxwKoHKksl++CaPV74WOkmcJOEH5OiRmVAWeeJ28+hFNJ+M/
PSRVQeEqhKDRlEQUl6aYuYHLhHAd+YhZFiUjtsMeGaPuKuItJc9yVuuwxiR3mbO9
4XfF9Yq37mfbMZtWZ9OxogEY/7RAhjLLHmTeLmlCx24E24gvC5xueJLYHLrV91c6
FEmTXSFkEEGkW4W2w7DPY21FIB00f+OqcCltAbPGFdEqShx7y3a8RjNUp8RtNZUy
+bN3My18JZkqADghCzIWdqPZtOjbyGlMwXJoWReczWfwW86Brl8Yexopppa59vN7
V2MQlug2oqd1eYdDA0j93FgCi4A1uulvfYK+6ohX0e1+sMS2BzlIuiixpfwZSNFw
8KQcUZqe+0CgP47OkmFJHihhBM3Xmm/EN6dn4O2WEzygBFmL9+wLqWBfYBv9iiSa
g0sUFWZUlzDMXC2FcPB/iVphR1Mk3O97hrHYAsLiAJmJVBxtfh97kEaWenEog3GE
PIrakDobYMF6OXvNYF5L1vSzSWpR0OG4fku1REfjrHiKHLB7z1rn+pI0n7KC1i7Y
euv3q//BiRMMhk6eXoIsMWZjLXLD2gmqERS2+X1B+ng2sQassasDagbbvVg5hgOJ
J4PA/nGCIA5Z2MZRx9HKFbroeL7PzhFcllzvLNAqP7LCkphue2GCK2+tTnT4kWSf
y6VMroc/KNHd5DIJ2uRJxZwZHFEquy7+pzkPzbuLoj3tLPSwPphslh24ddVnpiOd
dCyjtzVmJ+II5oOpwJgUE9MrRZ2qR/hrC8/mP8tImF3B5LNf5HlLW/Tc/FVeJA2z
hjSl4SSfPaf4DDHQL9LkzRSmDVBsDvErvuuOdvzCICAmb254kCJHJBdX2bXU98UA
6v/F023WYvJfYk+UsGQL4nbwkk9M2MvOdL7AaNr1h7JKiJDwkTn0JdWC41H5+0sV
5snkP7USFc9sbDrPWmdhJRCQiIQsg3EvcR0HdHw9A+HXdrI+wYZ8DGjaCJrOGNfq
5Ak8bd7ZpUS2CWQSdpE9aNxZ8gXu7i3b/kwn60NAxNV8zE33AlPGJezXGDF1gaiq
/jH7yaBqcJcvcGVTXL082HPLviCb9sNDatchKai63LSKEyqXEFQkdb4N9HD0OoVc
iMIu/tLJOdOviyu2CCA06mpmtJJRXsMljP6l/PPZHjpX61o8oQF/RG+H6TGdEXZu
7BIl+cZ/7Ghrh1GmklCzn1X5Mbz1pjdwt0K3tTGAuGfYgLPJEKcgLVZrUpPKDhsa
Vp2iCTjmb42Mk3ZraddbcJfxGKYbf9/b3LJuDP8sdeBLNFYvLQa1N8GUvwg5D1LZ
D0MXiEMvDF99MJbqcERfLuNtcptdez58r+BW0LREnEZbReSZVGdSjKc11wi3ILAz
N5d02JC4JkExgiFHxFImiyq/7mG/7zeXfPHSs/vS/ulMQgr4BELLBVq5DoqaE7Q8
Iqr/9aOrUtoBZs26BRxNlRceKhzNxo39c0XELGrTpZQcTQwIPY5sy8SwK5YvWLFf
Kya6SL5kIRXAlMW6Ikcsbdfe9OdgWGloY2+tk5dXN/ogJG9iDsN5DE3/tGnWW//E
rhURBIGA96gBohF2aa6tMSlF0mi7F7RceS+wbrPN3S5OAV66iDa4PnUvMPYRM3vR
dzBIT8WfR4HgJO/WFuN8Eg8HZM341x0D1aB1SgSVqNWgVFiW4RReNxufjSIpxkI3
BYcleeOr4SPpLwkEkNhkcSqbza6Q/wH8x2Xs5up4Iw0rlZuhe7KqRlKMXUngB5iG
B0+XsLqlaTllq1CZuLSSK5u2icbDFhvoKO3PkI1V9M79oEHnmjRqP8++++JsvmC8
+FcP5NqWxEQrKF4nidjiWmaNQkSX/Dhebw/fRY7W/+QA1QLQSfRW/YUjWka8TnEB
L3vAxQjweOBnKSxxvobIxAg635+eSEAPk8SS1IE0LB3YaoND1BTBOGF8nH5TICPY
oqN5xYAwkKZPxz0yESoPRowmnMzTxwxKSLWYljmztM3t7x5Kup2Vwprmy+abOvZn
SNp5Adp6M5RaqLVL4w9OAvhR3kU8UtPFPQAvt/8fcHj9wB1B+TRmLpbCM2ezhi9G
XDHHJKdMwUV16Rp0CsWmy5zNK8vBQw3miDUgPm/BoFTqxmF9s0wERmuBY2qUd1y7
+AzDohweTw8NdRvuV5dV9XuZFWi+dzEk5zUhVpaFommhjjBGU3XB+htUmGG2ncMG
BiyzR5jnu50h3/6ETQ3kdAo2kYhjyqq+VEVCcwwVDjLjb8CsOa99lBTw7Nr6MpMW
9EM3AZWH3DyBBjnqw+WKRIzKNigM+eFOw7KAcT22EoitRAvcPWf1jD6rQeLsTUq8
aXPnQ1RzMgLx45eBmjDhRewh00w6o731dYIYq85aEHgi93vvh8eL6XErz2ESinYf
Nvmbo2POvO/kBHfW5Xozpd1udBiakOXHSVy/MKp741oGLC7SGivOT+N0mloQKTvC
JdbLAJq2JXTPb2CtIUm9pKJv++tB4agffUXs6QqfhWaSmjRIwkOh8gdHBYVbnKgJ
txCAepPexM3mSmiQRyh/RLuGjLGGtD51ravE8wvcnr9GqpWpiU1V+NzkfAJENWnn
w7COseyqT0/R69MGZRKtWxv9x6VuGFQDkhT+Y9HZ/EBYd87X0SUtgoHDuOKFhWOB
sDskB9DY2x1oHKXrJq4mOIpE3DQBDU1sH6Vl8nbucPkoICJG2aRaMoQykDidMJOF
iM1JZuvG+nI4Qq8qw7D/Ta9tXMdzfWHfQYXYJo9beXvpQ2JTCAB86h+eA43NegWc
BGAIgljJ8I5hkDxEiIuv9G0G79chK9wb+ZtvbHd41Cvpj2YlW9Y74Zpomx6xI1oG
9dUchiLTTMgrwv+5M2GzuUCZWLofvxCQatl4EWHR8IWgka00CZpUJS9m2pqgG7Os
oYXehEmSk+p3QK2nM3ORdtuyxSydjMgUeQu8l4073P0wFbVMDBcdZ00CwBK+cBpN
EBi3XRv1H5QkLU3mmiasX4vsmkQ9CHS7oBj3xowIOK5TKvkWILv2+EW3BO2jUW6V
Wnp4jK78PtxNxng0rDbWrxMG63go5mWzd8FlKGKu9z/YkGvU64wAZ9uL2BNdegwZ
CgY1OPXUXWyro+AtQLD+bgAIChKd1+dyft+eWAVhWyxwFvUXY22gun8WpZHuhnWo
Ij3Uvm6NYhkW9p6CxmBPHgnB2JHvXXN+BX3dFQtY/qD/Okisj8hdV5OCfCtokSNu
K3HHCaOj3WD9N5EHBEDcPdqYXJAnV2WRehAbYHoCWJpQOJjD+/UAZ0gYd5MUtnz8
LA3A8kd1JWuDbLqYl9TUZ3oqiDZRXuXrP+zZGHeDZl2DLO/Nz4lmdV5b5wVsFYvV
msNuf7IxPyvDCUnxGB13a1vcw1hLR+/SpxSgdpJYew/SRbyLTEd8i1RjZ2cZIcjS
xOY2zGwPNcHw7UgFdx5ogDKY7LyAXVLXUdzTB5Lta1LI7LkcinpSt+22z/XbM0ye
M5TBOQ/QIRYNT5IP0HepaL4Qj3aJ3nfRD9Z91F93tOlSE7o21OAHEPdSEH+XIbjr
dWHeGID9oBMGZDxACZBCzBjRxWcxSjacHmpP0z33Vl62IRk0mEOus1r6dtU3sf0J
ybIIg0+mpIEiPw8PNyMmwYSbbZe0+gcqGAlXqGO1Mch/jtKiSu3zCt8/TCCWF8Fy
MTmFU2t8pvtEmtUKh9v2UqmhyaQjTmo4F8PNd7QRE5XD81nHbCVQJAU1bpu9CTZQ
beGZ4wSSK/b3enKXmpRZtWeP6JY5Pj26Yabu4j4sYba6kdIW8sU1A7UTGYaBZx8+
0Hl6oxV1sEu1u3UibcKASSd0FJ68BmbXXpZobYmIPhMInLO5rYuwcQGi9bMN5H9P
Y5JG9OoRr4mx4/BBd/dHvBkfz0LbcG2pdsBJaan/NLV3tvB/UByoPSuwSt0eiPWg
BZsRXSzBoyZnEYtNz0ie5nL0O6FSN00FQ9HLawbZybaybrNYgJFs58nWAg+afNiG
JP1dNeecHiMlLbkGFNCfjW/hOJztsq+naIX+tr6wNuE6Hr8BjQzm5ZeUv8zbSBYG
KE9nGvBIDxbz88s5o9HKhvHs1/gfzQxFOytO8WYlad2d/Qlin9c0W7xDg3yEez6O
kLI4JJ457X31fR4MPHdtxjO+9GXehQKAra7MvwH7kxhj9BW6w+3i4pWBVeD77bFa
lCE8WMPp/Hr0J4o1d0p6+IKlrpYpeO05F2myonUGXjZk2YUizw6RsV9pmycap9JX
UNJa7CHVaIWR3FkzHKslNVHSonLgUgtdclu1nGksh5YTplvIk+lgp5/19pK19qKK
GY17hnQZYfypv0Yrs8tudIAlw++00Wu8+7BkeEqSzpHBzNz61LJKTGSGD1l/bKN2
CpG5M8Zww/FW3sKKNVOsw+bPsOrO2LmpIYcbhpjLToejEm1pxAAHmCXiZHsLBDHU
DDYD/lnr/rm8PQTeoI2muWIBO3IFSkrp9LaXAATisEUm+uDFz5aVdmWE1GSvUeM5
JKLe1ibqjCwifGh3zUVkMIRpAgDLdKr63z/b8QynwezgHI/wxcEKOXn/y/c7ceqR
Sr5rbto16EcLmpQTmIo4I5surNG1IhmXDZ7ACalvmWx3YpPP5pqzN7ydNyTV3K0n
iAkGLpm1x7Apv8DquuvPXxyylbVb6H5/WnlWYj+U5CsTC3jdONBIA3GDubaRK5iw
i9NyTY8CqEhinn9YcsKSKPXHpbxGEQDZT61lRsTBmR6u74RVuJXWFT4Widea4W0e
2ThbcAf0q2FzLljqw2t28xRTrUCR/8PIy7VYp8EDzOgZ1PL9ziQmhXKyjmPbK+xK
LPiVnCGmB3LtzpkZDgncjJMoz4KKmCJ4L14Y07hNQ3wtuYUSkxCuaiYzLiZJ22HA
j7sESqevjyF+ffg2XInu0u+sjrIsLURyIfSFFaYgpwmaFj3pASMdnm0plLxA9+Tf
mMbF9T1gybrCbPQVUGod2xZ6QcJerLv6BLXzZYySe9VP+AZjdEDz3cPXWn4BiMjW
oV4XNGYFqOpM0FmIXAxGCSPA6r2LydMuAV1kLMbVfpeWlk/SBSE2T40T5jq0Mbml
nedrsKgtu/eG/KPWugbbevEdOpI3b5OvbyAnxKgcbBO73B2iEcgSU4c/KleCdxY/
KdTDV1kPaU+K+jElT8Sjs2PI57QILFz1XVJmTjgnfpG14YWMK8ZZdOckQDdK64wB
wTDm8DcZgxuOAMffm920HoOQ2IgWbuDsD3QH8WSOijQNF9e2SibjI91gnUOh4SOV
Mg3u/0kCnJJj+AbQFSyZ3ULvOmZ8huAeB9BKgsXUxCcrzVxc6j/pOJfbHN0+0yB4
LmkVMM8jzgcp7Hv6hqA9acfzmK88FNoI0jPh/pOQyZE4Cm8WWL8XCaAXFHErCeKv
banDGcB+FrPEvXRJuKYWhtycvXbKjtNWXTbIUlSq6pKo3rsMUU13/coge1JOQTlI
c5nQkw+r3raLnIag5S0uDvEKMgwNGbVRnDh8QCMCer1bU8rau75cs+QHwywb1Ggz
6jJr6nsR/H03efrAH6O348S0rDjYnbns8Kgxr/4Oym8NXKaUp8LJ9IX99UYkXrZ5
/L1FsDE2LYmscXOWb0GtSHsWCbDWNB5aD0ONpwga6SNoLbDKX7Bodx6nPvJF4Mnk
ghW68jjVglUB00sbhATui1icRbpP0vpQhQphB0TDlnGBr23We3hsmjPBClqIJIOG
JQrTOyJaQLUMMj5eHlBZbRTgR/auvZZcSBfwO3X9mA/TMpGrqJHYEQTVLsqZiXK2
JyRxN/FeK2eEjKThmIrVmbLTrqkpPddU7Vd4paSFRidsIsxotWlnvCKtICLzHlOm
8YDgV9bd5VMKyMD3ZXBB1wbVpKscutLh6ue/r6wxMBfHuqHKwe0HQ3EjhtOG0GBY
jjMoRwI6e+Xa3TQXap0KY6sMHp57/+/BG150QtyxiTIMakqR2xyocBcK9EWYLjri
KzG1xBlHIhGvRNTWa7uu+9DZJN6mp3GLvMIbUxvbXvJcdubD2Wd3JpZkammC6ZM2
DRyAGjcyNn73plj4HVHEkS6fUzn3Gx0j3sgOPGtqWZMZ9IsCaauxBsmQely+tI+/
NzQ3Ja51g/3d3mQ6/MLqYdS/qQbPzN9d81gaqoWoyoCwQ7TDvVQOxNaD2r9y7ENe
PRuGs6HT1zUy99IIcNZx012Or8wQ2IrJR30OztWbUlMnKB1Iru13s6FzHo+tACYA
c+hm0y/BpJxB8s8dqb3Y2zBep1kR72n7nsFw7OTG2bcrG6DYR1E7zhhE6Agoy5Bb
0rRc8VtNfa7GaoSrTKFVq4sKUUQjj1jqW4W73iIIxmZLq7oTAZUXjblIx7xVL0SA
K3Gz6M5pNW9OQoOanPHG6yGmdc1Yn4ryHRkmAxL8ddkTg31YeBof7kDiPhWAHO+k
qu2Y8xs63Qp7dGS3sKvLhErhXovHOsONfuWA9HqdeaQQPbHO1+cItAcmfk605CyA
RyQsc30FrKXqUDKxHpuar4ka8RwXtWaWebrfATFJ0h25SWekqZhu8nEV5QNvDD1j
8f185pXgWsppg6onaZKgvOzmiZFDSA8qNloW+KAGrLJSRGYeleKBNrhf+/jgmDry
M/27oIRFFOOMXbGM2Q30DSkbxQ/wCTaUP5mGGiGQZUoitshGwn5UA6RwuUior5kz
6hr41yRqNuhQQX1Ijp9Rmm4ogFzNKiiVKBX0kmLyvRX8ELcPnp0RaaGkwrL629sm
UWz09yxkxPquV6pIlzzoPJ0IizuF6BNBbk0mZEYFiFcDyDV19aLzShva4orkCg9H
nHNOC2rPRaMicGC/tZILLD+bLDqruwzv5+30lgcpEDM+s6JO7DgPQXNTWyghVH1T
3KXC6hBRwsLCbOORi6Jitc/i2FnkLPLKvfY+I54hLNWibOT7hVwiLf6nwYavGE4+
92XSm1MT7uv2Fg5S6xDWVU1E8jOVyQhI05CibbrB+e1epJ7N3zwYeIb27Afn/Iuq
95Kub1FamKanTEHLwiKIaegjGrh/oRNHajlsi8F7+qy1MY2rPBM7UKWpLuemDRlH
JeqdoJDFHIXsU6F6A8WKZu1FpyDqiSxjTqa+qVTKslL/7ySATGYJg565MJ58IwLN
2lGZDBfaj2YlDOasA8jrOBHjHOUh7lhFWTxz5GERGsyLE2QJbpmccFHocCXR8jV5
F/FFpO3q/jKIoThwKD6gKV/Of1mZd7YZmDjMmJQBfs+e4OiVwEdxvUpfP27JgFhZ
1XbVf4cfGYlznn5QAatXZm0GV+eQ3X9RRI0PJ0kqlT0Z1fQDdVSPlgk7IxKgWgyX
x5mFDUboJbA0k428LV1m4xq5uBDOgHkoLLIY/5mPZ4U2FGr0SrVQxNJkEGY/uwP6
YE9E3qGOAsR77trl5qsBDyW+VndeAQhIsf6/pxhWH7ukkLACypKXV3FRoHkbvmjR
ycFI8lE1PqZjGLqy1kmbVmaKhQ6hiQNakqqWLR1m12ycVN/Y/Q/YAq61bBAntLxT
zY6Kp7YdFKVfDJLjinkQw145E7Ydu85HK8zqBi92bbVLpr0p1HeDrA/iSUYt3tJn
/Gm0Vd2K8IVxsWvGhCo7/j74lzBKl8/l0iS/6NVIlNHAe7Ymb4Q0rTfgoUBxG62E
8ykJ6Mx6Zmn0Gz916SAnVn2eTTMAbeVhuT4Uwd4srsH/MMeA4wwOXYvDy5K618DR
a8V7DLmAZXXInEJ8G4gqMrClM0XDOuGelv+Jjr5wTfQUJoXAVPDMzTbGzffrgIga
I2ooc8ukZIfwySOpdIvCVI4BdRVMnbF9HQkOI9h41LVTCJvLHgWNpzq+jQL/6lha
1H3MCsPfPcorFcFZKRRav1DdD37SFyMBUwRAF1tx+H5R6CJqpGZvoXPO+giPod/V
guel6LJWk4OYp+y2MXWHuOa+iqk3eisRbGJBszKn+K5XipoQL5uwpzEj36nV+hsn
n4h01FFsghtDq/oQiWeQ1PG/Oq2A5kwGAhJmfCzNL9hzfKi+XOelCg7Rl1oPxzNq
NqivsKNgX7BOgvFGfwSY1y0XCAiYGXfp7gxeebpC9/3IlgdND82EysNro1xRP3el
VzuRQG1cWkjz363/JQ3XN1D0vo+SP5IEq88+TrwOjXCLmkj0wY6g23zqwz7/W36J
aF3WTQ9nWWHGYB5wLoUBdFmasRQ8GrsiBlb2wuHffY0fVsg68rEo2PUBUkuohOiJ
geclXOxRLspj/iz+HgjlvdzvF2LoPWQO08BsP8MQmCKj8bFcTXq/2YLuO2V52iBu
mHDY4LAahnC9mkQhg0h60BkUu/hZRASCOxMXI9vlC2g/DQr1mCcOBbAqlBHfw1Z/
KUH+nypSykgpHXj7fijDonZ6ZsimouxANIXXPec4AHuwiJQLoTf1CorC8CRkdXHI
8Gn0OgLalQICxehM8QLO/rga8wa+7jtKiw3ZJUaaiKOHUeF08Z2+UrnrUcw5iYui
WWqK9ik5oE4fqOxgHy+K+g1AGJwZ62/dF2lXAKAGIg/EnU2ESbPrpqM4kI4eHMox
U7LKiJ1Jsx2g0EJVxBnoMmLd5eOOaoTLJg/JNLLNKUuZn3ZcVZXDlJCbprC8+EME
qMPAjnkshng0ZjsDK/PzrSNpcUguH2DVmYTj3Awf2r41MKGYZSuvhNSdCPpGSlxP
i75fCFYikw5PTx+87nxqwoJruPSsqULVcIwgxrf6Q7E6oDiiNu1SIHgPv7SP819c
4eu9+vMTjyYsJtib1tvbGYjFjQWeKMoE4Um8z9QdwZrqs+UUBbdIMCbvo3ZT/9Vp
mRn8aCDHToHRie6ykEnn/8RvwYrpkOeFh/2XLC2+vKOB4CQ6LgmTeO50ckTUJg8S
QpH7Tbec4MWWhpBtXErlVbUBIS3PUhZgWvSYJV7PPtGSZege1Djzqz9TuO0BWw4O
bqr/Vk6dnr9KUBYvefjaToSCLM3n6iRURrbF3i9pXzB1TM2yUlfuPrjsI2+lqRuJ
x4rtBNl15p3suM/29AohMbqTNvRXqKdT7EaVocYCfMuS1TAK9utOFBuAf6w5Gm7A
+PMn0/Z3KLLpyta6qfkSzzgV3wMvLcY7YbP/+nWXjq/AT0pDvDli/w/Y4UK3bA+Q
PPnOKPXw6Tv3LNP4JAGZ0G/h+AXTr7/JIHJSWCLj1OfUtA09fzPvUsSRLaxZb1wx
ePXpvn/MxJQOwmw/J03vNylNJdB0y82m4EsDIdjsYzWkDIiStM/yv8wl8CYPF7Fx
oBI3DjFb8W7TAHg4vXV5MOndbDe2yihDJJ6v2J8EFAWoXT4fjIe04OeuXe+eNQ99
O5GpK4lSNv395E/xHQSnVFcuFA6g3K1PtiGHCE6A6b0HB5neFtW5d+KFZh4ViB68
HWNLAHH4ucNQEg7K7WYNA7UI+eHNIr3LAAy/+aJZj8y7Kq6KZJqvDvj3eWRya2mq
QkXmSJ8Q1g9TDPhc0i9QotauV8A0d4ZNz5/T6FpeR8cg2TUrFYkPLriD5zh4Yhdq
zoJCI3KXspl8U+9isbeQEKZlQR1QBqvIYqs0uzrPCU9pL2gAgginQ3JKkNfo+nMW
sLWLNopxl5AhxqY87CmvKJUXf0Vvwk3AdXHByQcvdrKvxbUDUYLEcMcIODqw5agS
JP8zExpiNkK5qlOXz59wRFgUV0EyaN17aB5FYxjFtlHBhDKZQxGMjwhr0HIYh03v
9Md2ayKkWkGgb8iP0XxXSvknnS1ZPX0W/hfacOQd9/4SmrFJokzS4V3Crx/O/TPz
2DfuQKLKWrFUmZxjWUJLOXlV9CZa8mCepDtP/Xd/tH1olzzACsAGPF6IxxL3WrI/
wKnEd+aRrTKQXwYlv47lrA2Ztb20JX0Hx0NpC7Dgdm6qpNzXA7VInrtDwaPvmDIj
t0PhSDZ1jz7XD4UtOwa809gYz9VyD1OJmjBBefYdosxvINbFbyJPfaiLhr9PohVu
NfxWnqXerCqpWgQtHmUHIyix/JVQu2wBXy9TZ3ZGiu7CHwjGfAT6vQO2IjcKRB5I
8PKHG3OjfY6Qfh1kJ3j/BrpofjReZZLBm+x+6hBLuOkVgDgwDUeKJSvyIuJp1WW+
zjiZAdk2291wdOhDRQkzsEb/wYUWnHrV0PIHdQ8gzUinIqcPDpBb58m0M4vUMEGm
sPgfaKyGu0Qu/cIVcvPS/c2gHu0q0BKN7IqBT6NfhNIUDW21LLj/ZV4s4VRGmqct
9Yu9xVRzWfCMCZkmKbqoluJNWmtfim8KD8mdo/zcTwd4twQ2jefwGxcebJ7Ir08K
g9C3gynlYYKDu7IPKDTd8/qR9EeKvomPUJYvbRExwfx/m6avwE/vEvqpuJsbV6CC
K3m3P+77+1IYUmPQ//1DofgfSqfR4xjGu/bc6BO9Eekq3FnRsEeQAkw2suKMAyxB
swCclVjEmIV8UOI+VuOMvBE2/NKZJ/9hqBFQ2StasixJwB8ppPWjCai4umzm2+c2
H8yGhHGBkFUWbmlf5mw8I4hpzCRP+YE7MRZkyrTLwlC1epTWMU1vCHeT4fyOZOrZ
kDNLn+n0qWF6vXmUEnE7/vJ9ZpOwx0irFTnR/17w3KduSZQJapx3+jPU6Vzz1Hq1
YOOG6sTWgGIqwSeJXvJ6G07OeLKdS9n/p8nLv5sRSARLlK57YhxdO2Z0b5ukWk2T
6csLHzSiBt6dQuYgPsnuoFuzugMkUk9S22rS6VT4gPehUPsbNz4luvYnndDQVp5R
l53SNcwlDUqu8qzl2ywObA5bes8nsyOR6sgQjVICGm0PAAGg+IRlGA1oE+x3OoFV
Idhgpyy8/rx3D4gomwpflkJgpaNQeHEg5fiv7siSitSEXpnBJOaCRzXxNengCkvz
cVkA+eQUGKijH62ocXRG8lEh3O6b1CDboAT5eghzRFo/Qh+d5pRSSvIAvik7a32D
rio1wBCOSVmbt1Srk3+yuRG6rnH0ihQWnoNexg23TZRRjruu3g0GwDtKaqCYDd3a
kX5GtLrBYQdPsCw8lj4boY1PthVloxu/ml+9Flw1VHJ54TRY6HjjFrWq3ngcRqIt
9jfChKHQjoGcJ5VOrQq4OvU8/d0I+T2t8DtKTQlcKplg6BQat3hYfhH6gpUnT3qb
fWeNeJgnPryPv521f4FHEPaYvEze1KEG7FkvlqROi5nsapZHDx6mfJ8XgmRuseDT
k8YMd6FqnbZg86e71tmm2xK8kpkYUMLVMEtdgjdzHVpaKe644sqo7JL7PN+7St6R
cNkeZ2+4hqGI1Ozc+naEeJD4aCrnG+6IuUB496HhOaPbUREW4lek6JMM7sOHUHfQ
h7IVkcF1dCxVBQ10uzJes6UlqfarIkjOPYSEMrzAKAKMVlVI8QeT8l3Vq0yOjvbh
jhgUK+aK/gvP6YoyfnfOaWu4MteOvKZYS+aQfBYj2WUwrh9d/jUbEtS7vxvEOocf
379b9r6a02HRhLDeCS+t8L8PYmW5uNy6LwEpWZC6pjqUPP56dulk0X531BGr/L0l
kBmzRnNocpKxmzsAfl74jG2om5Ko+ojlDrWtbrBb0A/xHeNvqCgrnZoY+smKFjYY
55//bMQJOFsBjw9Lb5ujrmv5nnMh+JFJZe467Qj5uX+3ob4Yz4SryM7/CFZsxjmn
Lx/DuANf6ejMy3uNMV0jYnB00rDtRFF9Dc/p83cXqlvsxdyWcwwLg4Gqg8Dw1hKk
l2BtZ50LnXSZlYOU89PNfQqhZEJNzEeIrgxlRiP8gzM13NSM3hHNHTJ7FBpPBFw5
EJSRXgf634/2ib37GB4uSTwP6nHkeJ3Yn07OODHnCelkmvqHZJBxIFy0uGFb02zP
LdSYtTT1LCniUhfJqM4GsR+X5nulqefjFzT0LH2ISrIl5fR1IjMYZgEJyaTiqKpH
wdeCKjo8QoDXANyMCSS0IOQHW7+r9EDR30pcwsEPq+77cmsZ9fZO1fCql1s9hJgJ
QlRNi73JW1Td7px0VfumyTHYrkeIHV300C7uO3M6WwNMuUCiywKw4XMn7EswYclp
rxBsbg8uh3I9JGNoInLSMsXeSuMPyYnaTO8YWv4MpFdJ60BeeOU9hyuaV6IrzvLu
0pLxGV0jDFEXHx9RwIIujv1uR/mG2j4XwzMWXHXd4im+tTFJAlxjpYeh95mh9MUF
JLusOamCy3/Vnj4KvyVkUdlzvmHYt+5hnZnvpDV8dRFk13UeE7IZKfZ/wSacAkYW
8U+u6M4T9R/TX0kbYxCItaqm4YZ44ONSHaWKvP16y1TBBU2/O0IjcC2JvlXLQs+a
sm5Cto1BHVtXhvOCoo0l9bWoque9RJVIVA8kecQ6vHeWqox8iV0TUEXyhK5wmjyu
pgME8rs4E86S3x5aUC19+KcP9KvPwYHTzobV82ewV4oTe9Nq10pEGV0LLthlokho
lW+z/oTuzmWA4p0piv6HcwaFytn5uJaCSvW9syUAHlfUMbHPFnWphpEgWx1VdVDy
olBCLeQd+ylfFTj4CgdHvxDythcmO3+CH+yN4V4xEH1li6iWhWgQbtrAt6HJzDab
zJ4LbPvUWp2NO+0GHtmemIXrpHqgJoHOAnjO+M7/y2WoAG+jMAI/b2x45cooiA6H
zWrphtul3qdqsYkWXN51/ij3aaoUgm9JnVWjL1390F4Gwe2gvLaqbyRCY7fFzhuO
ZpD+kasnLYWWUKx5Fk00PtWQgVK+mgNr4euYhfuhYFX1ei8mb9d0d3NGLdOphomc
n1wdlN0n2JQ77hr6EI9fWEzHLiYHT21NVwEdpe3+V5Hv7a6BabH1UKNeeoCYqD5Y
lCBzTLtMQIS9lMhu7ykRVNgHjGMUyUtZ0wNptMRdUD5bYgQlW76CRlUNzkzauha7
fdA1XucrKGMuwtt6uPxwr7gJkEVGBYJhP+mBoiLlWd6WA5ik27eN/6b50Ic6pHz7
scPmbtfgj/7PZ8Xx2BVI8U+E2ES1ukkdSWYM0V4P/bjLV/vJx2TeeJTL/zCSh7Ie
7ZhsEGZ0+dxEFcvOLd2uAiyIu6ax3WySdVlyJ7VZiv5VtcWA0nkiYbLwzn/kmvVD
UCn7Iic/2I4NqpXlCoMY9OxL0AIe5WCfIXa5T2GyT+umWGeoWrebHS1DDwW8QBQ5
wM0yP1j+bPyv5BM428SEzRoCuOOgUSuJvCLY1YEP6kFNWJJOb5P9aB5L/9gFPpUX
PKTJQI9VTfKQZY4U4zjNDN8pN7DDSDl9VYiLLUle+5/uzxSETgd1TnBExRFCRAO5
SA2MGtpErfwSZnkakq6Guq72DHrrqnAspT/CfZn2sIgyKz1Tfcbf+JhvO7KZd7wh
dIJI//EmTP7fRm6yfGwqoool/IdfhkzJOmIAw3qleAihFpRSVMev4ugphadWvfNp
i61WvDGIGoPWA2OxmhfEUBvnO9uuxlzyeVwCMz03v6fEjMtFgFNEvcge+BKgdX5T
ktepalkqwDVXGmF2FBlXFSMcrS+N7G2okaRJrXj373elBvCbAiu1ZYtxFm8kHqNi
ttHajVT7U0l11jUQyMI58ydtrqvq0rhXNhKwhbOhCYvJf/zutxsO2LHRaZsvGWHJ
Bk1Xaqon4UHth6impaiCAdwbdu4nez+olQP8tEnFq+mvNOobysew5U/ypcXBS2lp
9MoeceCLiu4G9tCPvrmbokJ2OtZ0HG3H+FTAwsZyYpqhjrYcJor3B2RMAcyzmFqr
MqLKXY03T6IPxDLOZ8bnMrJf7ujEZUnplS+pWXuWGA/qJVDoDf9zlSiatZFizLou
fYWKVIZD3/M7neIgvgvcSqNtJQJeTi74ESQkS/Jjh3xN1hVDCOzT1fAY5Jp+qsSH
EEc1Dz/qW7MvflYEJm/OwlTdVCeRMgaMpzQB2wKhWn+GCG2uC1V9xh5MYBKBvLtv
szb5rm7xFb4LvJuWTKtvw51ocjyUJJIfMaRgarBn5v6ralDUtG1tQlRP7Gto0yqS
i3yZvquJz82FRCwsLwP34zYeEYCYJZaD8tDnf7f/rDoowDPx/sbmJqFQn3i9BPbO
vVOCx7JATOpoveDQqmCOX6g6RneIVBddLWbGxobxslJpRYKJK3vrw/4kEYEL0vow
H4bo/seMjSFbv2TIvxntO5zdLSDI+HspBO0QQlRKOVtVaYrLJdQ9cL2fZ2LX82bB
jOZn4G151TRFfNbdEnNBpnGXrMIHXdIOzZzqVwlqvKDZhSgWZ/BGY67zvf1C8i/2
bGZsgYOTMULQ5HGjB19ZbV+3FkoCEckNPqDFg+z4qrkJtRWuhlHJsPbFzVtvoI+3
ZtZEXnRMMVS+vvsv9xvvnPKapfmIRFrNRgliEMpjX3tMdoJJpIN1p2yNiiAazm8o
SBjJ5R/sCDX8h0Ze3Lx+elA79lMKzy8Thrwm0ZBQHuu9oXRvbOMPyG317Pkp4mky
OaHBVEnLVKc80Yel7j+TN3ifU1+WnivZfQjZVE2rsbMRZQLwMMb1mrb1R5CYCrpQ
KlQqNx3Ni4T4GYDcG3Jz9jVP7uyeVuQwd7hAeAdl99waOVqDQP4W6vGzXMttP5gt
Mpwi+vYPbhbeJVE5FJuCThMXqrAielESv3UwNP/IrHuDmLqo3brqyIi+pMLEXmwL
0u+ZtsLLSBWkGbIlTz8lWEyDzlSnqPDQtvIxRc1YMBZhA+NvFsc6EIRJxeH7O3Ge
9ihaJnFCzADyoecKRVL1HAOBRiPFf9FSI+EXPYqvd1Z8n3Q8oQV1wqlleIJoen/u
9yOsfdRUQfrnk751fbj5mxR5fNkgscxwP3IWjUIS1wyg4WhJ9jm8kNesJUYrQzWL
0dC1b9/xetWagpOH4Wef8JavcyfPmj3ow0aooVA7tXUK3qqZ9PRzuC5UwEDsKM0T
pxUjuNWig2tW7xZAQkNoOmkznvcS2ao3ywpAyTMy2hIKWWzXQfCS7E+Ab5+jLZX6
Cd8Eu8oLfpDlSxzNon4kxWk2Wr3PSmt2D7D8dRiRVv0CF44sQcBVwp5kQtp5JF5i
YGLeibAlTFnOMSksHgzIo9KTpmeWrDOAs6ADRox/KwzVr8qxg/OjgEencr9rIDtA
galxZNHVDsUQmy43dVoa2uxwpx3pQUz6Kd2WyReEU776jxZD957JNN4Iy9apMKHp
IU+FC6lNPrIA+tQYkYqHc8qn5lXmduNe1wsy/8+CKRbYMT3geXGie11Eg71r5kmn
B2c392HVOVZOymtUiIiJk8V0oEoABNJG9wAcsX+cRUQbc4Uw6Gt1YBRvzFUrevbF
W1vqTWl0HHz0TLjKzxUrtmqxpME5+nt2yfDCZKkztBCkOysgpzIeon2yDSRuYJJP
hzE6J1+T/B1UbzHutkn4TjCZ0HQwNk+ur01P58JdeVGpOrPXi17fPml+lu9eQrDK
v08+JKOMVTxZISHcY8nLgccbo2oEUPk+o2J5YYC2RHxOivl5Mr/Dg6E5JPI6G6iW
ruECJgEInz+tqUzMYQ/bw+Ds0uCEANaWFkVoWxqiW5/2qWXw0vN/eSkZrmgEtOYI
aAdTOUhjwfb9t98nwPxqPTqQ/GFdBFTvXeU6qddalW6LyIW5m5LSBAFna7mhBD+L
VKlt5yU1BW1ZqYpeIfv51CSgmP88vSydzgei/keVU/yKTcv+aHnigJoE2KH+BflW
Nn8usFwbDD2n5QeJq06DD8js+UpAG2XrKvkddJhVf1W/B2eVctIGvzQP7ubWJshp
9Qrt3f2/iArt0wrBoUxkEM5YpO596FvnLgVLd4U7ten62dwDZ27Vp9LdqnOo5YGV
Xcsoj4C3D5dKYD6Gi9gjKbeMWrDWZ79nT3f+sr8wwzqi/tNlB+LppXlT0N9OdnPu
ycU+B/8P92NWlO3O6slRETiQml6SUYZHAMHrOdZBaxcTqhxuuhBwYG7MhIOVTR4z
6zV6QT9erTQpZxKPgbVb/EwcETluPYNwZv2uNr9/pdBgNy7F4iLLYWQaRC3TCVIy
fqMEqUff2GAUNIsqV++HrtWB5QIpVbB8IkVCGEiBGW3vwHCXtJztnYX1DkYaHRWF
m9MlKR0DHu34njVYtYYCRNXFiLiqJRKBV7bCimDu+n6aZED+WxAPCmrsLYxBitVz
a1v7KbDw7iPm7yOMj8fZcYiDJJnn9jvRjNp1hrkqm95cXNE2KII1JBbR4mhXp8lJ
X3o4h553mu695w06T/uz2N7uGrD3Pto7Yfnpttv9hD4xAsxHpUbzGW6IyUtgBMMw
d9xaxMk3U0BiGAIsGuKGcvHq8pfchOZqv8/jAPG3gP1VHVD2FRysCf6PKWuHISfa
uHhntNtE4wPjfR9DaSZmBnn8EBQ+D0Nyr3j2IzXMZT3QDIy3uOu/qeu1K6HH40WT
WvACbv/+uKRjt7rrQv1vDG+4RWrDDgokDwrVRmabTJphoVT2CLafTi4fB8ayTADb
OeY7jFAgR6QHV63vpKn1i4kGVWa+USIpY+KQRVYfnz3WT126abF1gFGy9kJqDFWK
yIojBSO3ogczTKyz7uUDgEaJylW3knY23VdxcfAeRVqNIVtrNOQQSRglkqTpfcFp
6cYboaVvyCq7sHVqEpH4FNyg199ZR1Z9RQh4ZfxPkkUgPZtkj7ilE6u7GFCglQDS
ZPHUIofDZLc5QcXUlD0rjK0u/OOcoeAzhjQJTMCBk/Il09HxgRSSRZUpixWsDwLL
Z3nUge11kOkDf6yInf/jXg46pdUX9LqeGOO797jopaq3hk3zGGLwXFgshGhlG/Qo
3PCtgYoAatTufNBmTGBuAL35/hlbRIkkXdWm9+SnZ/XFXnofUXi895Tvs4xOiFuO
nFBXU5uXESevZgBIgBT65jCaMFKhv6mzX2PqNVEfpRZA1SsnmQzBA9MAU1JNSl1G
i0HhgbiUnpnQ1dcBY8/QboXVmNye1l0RmsviLacB18qICIAbrheoXkN1UwUW73wl
7wf/v4zNaa4R+VhmVzWNZaIr0RDPcDd8TQbBtTvn2asIYlYhnEoPoB5ukGnqCcfr
bXj/kXL96zh5qXgQOiMZ6HWn+tuFR5nriFhsX66zkwHP/YSptM7MJAwsolT4LDtC
i+/ouC1kgr2IEpXPwSqyiUtqD3KVjeQzUKAYWYieyeixojQ6f8EJVgZ062Yr9gyP
QWy7uHJZWzUr4vSsbpeRTb02tQy9MsTi1nWHDvb9rQi83f9+0JuFvOBf+aM2xJuK
hU5la7fUyI3Iyc8gSwyFXspSOe1zF/DccFlsLdXsmgpXYpXHqsTuAwyAsxIsERLT
EYlo1LlHnaAyDx4f2ypsA7oAx/Jht1dJ0FcFP66O9lNGV+XTrPk0T4eJtdvXEbty
YiDZ03ZN/CSQ71TKgiDrTia6bUpSAUB6GDkB3jvmkNJLkYXcoui7ElE2JkT1HMJR
wNzDyAz0vSYcQBjB+t6v6yjJNlsCwGmfiTkfvcp0V/XEg9Nq2fR//P9RpyMEFotf
VB30c2eQxsKvZFalm4L4P0tf9BzcUNqnBU+xs9fMK9s2AkRjeSMZbVTLO08UJV0D
vRKRtkH79fhuM4VLSEA2TjoR8vjlA4JZ9568H7vdXO1FGrE34o5V6esOfCY4fX/B
DoIes3Wk0C2Qujp+P6IdwIifEkLy7pYYxq5IrW+1KMh7dQYJBW/4lRq7LDVC2AIx
8oXS/ZdmdvS+LjLom6pECFRTirgWsik0eV70/cQ0SWTUqI040wQT/MtfBCjAkgux
h75ctJPiZLeui6BZhl5f/1lUPzPCII2N3m1HwM6KTCmFB+NO+ZiaboJtLU6CbApZ
qcLDBHpgfdayKzmX6VrgZBt3p7sXDNcPuqECf2bMO7+X7/Ts5REmmMnMTrgMpKMy
NeR1KbG0y0bdBn5Md+IXvAsS0D8h9OdyrP/MozY/fklh49N6S6LX5HIR7H7/v5IV
Fgpq6vXdLJgpU2RBrgofRXK7PLZeX0uzNm8gUy6Fgq8lpqqD2iV4ZTfOoSYr3T6Z
IbYw0LC8RQTfSxSk5ieoaW//AwoARcqoP/MdeIDsCcbH2hmZlJdBbO1atoRlM7Io
HHPJkoi0KYkX3KxKgJtFhnxaNQUkFFOq3F6o7IGndPJF8rjxJhSr+8FhLUR+b0mq
1DSw1ogf93MgHN74RP7WWJW/IytVRSG4Rz/8mUCadU2LSHQ2/vpSS7//4xLdp1qQ
8T3hGTT0q2fbnjGgvZRLh3F0X1flnsg0hNG3pbFLoETvSuQ/Y+ckN7LBoipK1lQq
GkVOMUtFM1BSI6+saBmrUWtcVXXxKJ5EsXvSjIYuhXQoPfQGuqgNIVnt7O5WZ8Ap
PsM/q9TOtOtPtmjpwn6TKZzTUt5akKXRfGYY6MaqZgnLvM1ApFfJtxoDYX9q6AGI
bcvbBdqCq+kQ24jcZnpDoR+WSMAE5UGX2ymdIhOnX3FAGfgn32guFM1ogeBDm2RI
UE+IsfPeSymi+oBXsLKwqW0s0x++wjlf+pUjVRH1xHKe/9olXRvs5/Hw6woj73Sx
ieYDUGLuiGr7FnV5xMTsjl6KApwfsCB736IYLb3gdT4dGpKGSmrvMLOJOC8IRg7C
86QkmofSYgiXV34x3wOqzPtkRBPn+yySrZISYHbWdcvIY9V6GHoBjme57Q4HTq4l
psX6ZuqgJxTmXiGfa8SWc2Pzst6iHgWKXffEsA1MOKUu8hrI1A80NXXFJWts24Fk
ZwQhp+noRy5tqdaeQPxvDaXgq/xQztIY8mfaytJm63InQ/vdO1g/lo5/2iyBRVBk
hRmSythnX2FDjS+DjR1C4bGU0a8Sbbi9gcmanNM0ThwVMdh7KlCiD7UmgTUbFZ8o
8lk/q8EM6Z06+8lSB0hgEbyF2+MKK9myz2jyKJZYvvFnMSERfNpTwIGhjFF7ITf9
1bSX/sozzFsy5xveoK1GGR4ESD1nNGc407JstoycElev9Mm0HNHmxEohKba0+d2D
0CkiWiW0oZUXAyoqxonZz+nk/PWNBno6a0yIkInq3RMcqdWVkiCUGhsEfdkcL/ve
6sO+KXvGPckWvqr3TfyuWQkIzNoMba5uynW5w4VYCzmCmTywldxZHbgaxOM9bBqU
uEURcEZmdOyzDWANnaFxT13+rRjqpO9Cqtf1zHB0Gk+5sRug0oROjS+hyVYBIjd0
THlazTemtgsaLR/e3LmJxlxHqPXqMTZcdmIh9t1Au+K/GbqNbpr/5wXodmc8LuPo
0/U+AznCJtYiltN6knZRGwkbCo9n8pURlevXpp3JMDx/i8ccXFDNympkV/gG6CPF
z/MObjjIOCfmirO+iRULU4Gd+pVPb6SpRbQzCPm+zJ9hmUUSrM88IRxTLoTFHcio
RWPtKfAWFCoTfrm0wFcp9ZbICoyYStaVCgpqdh5z9hsUy4pM1vqpTkBbwoK05GAc
v1s93XsJItP1+tY1B1jCBrGWgzwZ+ex8qjjwkAM3t9RCCcYOL+wjitOQMO4NqYRw
ARTOPmXJwNHRQdo3AkNAshSwjU+DROzUb50WzRzGXh6EqM7HzvEPlLPS8k9f/4ei
0VRvtQvSBgURUyV+8utcIVYd/kEaX4f2WL75G0MD93uFpBsOZQJCaBBJ52XuDXC/
6aeqOrrhq+Fc4PoD0JVL57x5QIH4bgQRUnui9VMksgei4jk+D1Pp+RForwl1LjvB
RfWp/yhRY1hcKUx+Bw7Oev/UgOYODiY7uS+sTBbMOCJJtoZmKCLm8bj2u4/+aFv6
hyAE3l/4x/DQBh7sLJ+zBN9eKUYYLLFlvXU+G5C6GzufXIBw613VjC+MVsi7HlfK
VG10Rclt237+2lUoMdWNBt5bgramoo/aXrRJDu2f56LcCs6ERk1Db3Rdmx7w1Leq
3wZ7h25L9O+n2zrZ3bBYbk+b+qHH35pingD29HmGArlCdwT2YyMdKSqHlEAI9n5D
GPCRNIYPf4TugQS1QzHrDCM5bAZ7tHyisQVSOx2bIRPRJeLDE7BIoJ6C3koqABv6
yLhQP1UhxMyjw3/dnrXzJD+2J3iXg60pjqBluWgxehA6B0t9W4ii/N4cMKIYPY0m
qJrVqOVqr6XqQiLwd84MueVXPU64jlKqTeWMfYBE3KipJtBE+Y7AtPPYxkWIwv6S
pBlNOBxOsxSsp/aYiLQ1tKfa/s00aPJHvixCo1c5bWOkNykhNWBZY8gaLeFjHO1I
HB7vGDWxPezPGvPDOLVwKa37GCvtl3QppsoLdnQUTh5Qqdg5YE+5tFSryejHF4ZJ
6JcX47WfiW1n07Nj6RfW3Sr76qoGkCyobyE1KHpRRRGWj5kfDB6wzlBoNCdAIXln
REosOiqv5PQKAIDZ+fNImkgDRX+aKgZgPic0NKws2Ol3C1liqbbTWYtbHXD3LLX5
Kr+RZLGEnYGO95oDxlEKSOp7zyeHtDmy5+sZ3J3A8buD1JSosDcCQrmNXYrFGR4w
RB2b/8k7BON+u9i8D4/haRvH6lIZ00RS3YBRF+KKXXsBvff/KP9D43ivCXgZKmZF
NuAhSzut4LfAw6LZEIks9krzyo249OfTem5izgxoIw2l79sQxODqwBoQTTeijtaw
7Ymx8WgcmksuoRfGSORtUhwzyiaFn8XCT79NP4gOt0L8AeP8XFPfMRU7rxft+Wdi
smiw/wyiGE9cqMPQcZPuPyxl/7ZbPQQC8zIK4FGvizRZ43H2fez6+h/p9wV2Sl5+
19+iGZDJqhU/Pvi4eXnfufAs9hVFLy4YEIhIhxE8puSmzBzkNo9Z9VltpY8W0/HA
FkYQFGTs84vzU513wBZk5Yoxszb2M4i8j1pqooLHUbtw3ftG6CaMPfPMM6EAzdwv
gkupe4VTg8LzcbfXFounZ3toF0hihdGFh2a3igosEwoWY9RS0YevX2BDoXLS+qIa
RfJ20nitA2GG/o4rtFowmusjdQ2KTEpf69aKtXvScGwCVt2ArBHpOWtjayKVEGrb
ivvGDQJ9eAg8DiBB2G9dVHDHvHGxLPlp6kwOok9+aTjk5ZDR+/te6zl3/LxJJeqe
RfewY+JXSbestLfUNx2lPktHAu9pOilzH+Y9Tu1mk9hWWpgca+QQTCDjz75d833y
TWxTMbh83EyM8fZmVZy65BG3GMK3gGu46gOw+Viw2QnYpwlDzaICx+moNYuZe/GA
vm8kp2EKD6XIW+GXh8O2wY2YA9R/d5X7HHJNjgpaORqyITRhBJ/BObQilNzCufit
2GnST3twItSskfcGkRqGVhuY5MnurtC9Ry5nAeR0luuDtM0KIi8ghGkFUjj0Rw0L
O2ZGcsg/Q94B6tjuczCreySDLYm3iUWSvrIq5EcSrgE05gnM0CkkoGFMH7HN5xtc
E7RVx1lx461pP/1kbjXaDz23YD4vMNuTliqK+f4I8lqRXE1jwIlUb+6W6TwTd4gk
dC22Gzq3zoFskuU/OishLCew49f3Mym83cLvd/1sjHFHll3K9CSedMQD8rAgmNqT
PyxYEQ1CjiEVh2lFJ+oPLGgXPAWb6hFrOfrnKU+BvbQZ86HuHKMcmKRM+X608PhU
G28h+vNQ9uHZdFSbvWQcBZ6a0XkRgpW9//YbZBB8g+e1LDzr6utzEfAuIR8O70Mb
sU7w3cfN6moA7Hm1aG0FC86eVrYbwnkK5slKuz+jHCh+wvPeG5SWWbGUxp0hWKRN
B/U6mOgVu54CpxnM3GdT77a2mDRS85JibIBx6VftWw5p79YA277FMYvLmCpSrqs3
ZPvVXzT8684LgGXAprewuginvo9FTJfhQDtpNGx37a4Hof+h7eG7FCBycvJGYB3N
hVtFA3CZShvtVsBxsGtj2HkvuhrQ3L3pXbw32nH7iJqQ1HmI7beCM47rkhbvDLBL
9xBZMyF2z1UTFHh8M73Bb/z4bN03SmmizAddcT9pdb29zBko5LMpeSmTxPxcFCmu
f90ghlZGebSZFmRmoxhGVArBuQLNJFEH/fr/caiXdVkr/zGg25/aiBsW3raPYDjw
kGEyLRmfMhcyutPSMMpPDpdA7Ow/Vf1nA/nMNGXU7FOx5bynkrnHjDAi71oqmcb7
WWoNnn8KDECn+SQ5JZQwv8PxUKJpTkbZfS5pkdRzf3isg/BlJxSJRmv/c6Svc8tj
+LShMoUmSUaNj9WQS38ivp0Vsd06LDDtPmJUsUCE2BP8QxtU8IRm8PIvkEVIfMBG
g7KQ7PGD8QtSyupg5nPghJMzuw4hIXDKjqdULraX8Kcb7/6FSWw8xWI72fICR3yW
PKTlVy+7CFWakB9uHkS4Qc1QlJz8kUc4ji+zjXOaiyjO2ZoyHHMYNGUSv1kiEMwd
538zgCNVtW3VSqThoi9N4v9wKdVFN/RLHkPe35rgypf4mnJUYJehm9JWnYQyWiF4
p5WG1BzyxDM8qs2KOe5hyJ25g40uGWl5RcgWYX3mDtFP6nOb7/XYf8gNAdjlkNjS
HtD7fNqJ/1UPUNwYbq8wiYpMtDeNqGjFB6Ja/j1GjTK+y1OV7XN3qW/J5t/xQJuI
YbIJu5U0xv/N1xO1aH38JCpCgI0Y8cbx860pbdq5YOHaxRVesLotnN0eh9QhmmGX
V9TTs3THPoTbT2N9+uVgAPhuE3uPM5aUyfc/x8lyGyzKUcyYdIKv94nP1XXLgTMo
ZtatXrU+3m0f8ZU1xDOUk5yqe39GNQorYCPpPWKe+AWn9yVNGYh4yt9rmTd3V2Hy
itxWWA9vkNnAe5mtfM7+Rmwi2+SU6Zx2Gt85EiPUzIo9qeNtdAPCwjrtHwR+4jzF
ysCDina99rRKXFWbKHiI2p8TTUHK+6oUplyGJ+R+QPSOdzjiTD3ShOyTS6NsJIMU
EQnZIMrCdoEwMebpT6E/46yw+z5+S0jrYeftPGpRdxr9WhWRyCtd/q2boXvhg3Iq
b2XXrZTusBDGdNyQ/hzFsJmG4Rc2gSvv+WEOUgLoYYrrpbpVMkTpmYTniIFb8Wqb
h1xmIaTXogXu2IQ/fji36h+HS5nlUeNsZ3+E86EWP7YrUpa8w5zKII3nc9hclR5D
OUoOSawAhr/1mdZFnACCwws9mL1mrAFRy7gNLrESPySe19clKRuO0dr6HJ3UuvBV
K0FYFU23DaS+dDDuJLW6S9Tou6r7w2oc80Jd/jtTOFtK7x6jVHYlwTV0D6CgI8z+
8CDH3hEmw1Rrn/9aql6PKJsiA+IHItegmijzy4sRQjlIWWM1ogIkVRgoCikwWjEE
evPFQUCBQocA/RnuwHbpJJGUt5KzE+KPbcsjnBdcv4J7scsv6i2LSJIcycMx7+XT
mD/t+DlGnm1PAOWeQFUlrdFJxWEF0rq/xwQs+woZD45p6HHaVU5kOoQh0F9upbvX
rZXhVCSp55ZBuLuUByg5Q1tlbZ5jo7x72ZEqyMnk+ReWpn/lTOXORmSBZOoicbap
ikL9Le9HLGxOHr/I7CYIYsEVriscbFe+tcCwIEU0bSZ+2qFQMr1d3Dv6Eynzmzsr
1wnqxw2noj+OajWCKHhvw6WOGxsWD2Uk5LCLHoO//G10bHvbrs6XM6QMWYVUsb2C
Tlm//kFKff2w1pi1IRXgQ2NcMfbIT9YFIkOw1Znxg3O0DSnquTtvDkibQ0H4qpXp
7W9gY3BF5tv6zSNUlabRJIOlSnnc8+OJX4CpMlXNZdVObPJPhuaFLxB282kL9YKN
hZrsgd/7dnMwE+32sy+CbwpviqpWTAKmCVT7R2GVUvq6p3z4EecwHPWhHFbbDVwP
NwcTtjptfrLhsfoDrK46g0F58HrHOiuI5YNIH+rO+/1Q0/LXI7NxqB17EeNcDxWa
w5/gp4cFleWoMOyIvunGjSlFwEvtsSS3jsqoT26Vm8vL3fCdDtyk2wL5APcpE2TQ
lEKYpnNFuWcc/OgwZ/DHN2HV+UdQ3GrjTexgRKxVhmh9ZQyySzGHNqY5LCkYk/l4
PoNvidFTx7WRA7+utY8QCE2IB3SPFLTDpJJ2KnuQtSH3wW7hibl0a5TpxkdcpNzG
ugx8LsrC5Y9D2siWpOe03U5vGQB0OPpzWwelxmv3UsOfBh1O+XHv7vz2XvD4tq5B
04XuBVsWEwW6oFkHfLRndCO3s/AOlDXpAB1TeGP+7cFPIFU0xn7Ri83hvcoqPvIU
rhy3/HfKnMPFuw5CD98gt9OLX/oRAWj3Gpp6xVf9+6IIsvxVNklEzk59bXyH45yP
oHIFaURk6F7+Z3aatRipGzNeJ+lQf7+zio+Igb/NTb4o1ZoO70a7IL2Necn/iItl
wxO+QfVoog2pvwq4IYRKWkGAlmMbhxPVVYss4e/+kQ0zaJ+cTF0KgMdCxlWjGm9w
57611Kgf6YNidAlCHC/VVYicY9/yvB+I6KRf8+e2/FH1TyxF29FqTpdEMex4o309
33DxBc3wpRv9/lCklWeei1x2o/39Gze70APFoZDCXXF6QowyO4mA+2OHq4MYsEHI
J7qIoqLnFX1MxndBwJIIH3xcClZXGSrlG6OFZoG5414HlWqjr3JoQEDnej4Zd892
vGS/hxMVoec5MQbPkpi8HsdNDNmQaD+oBR5WSQnLA6pHOu8r2hGFlNTjssfdkOb2
ytYNgTdJ20tLfeLdfoTwR8FYlMZSvgSMMQmweOBdBuglKvI1VUsDhVOlPHFBi/WW
QM62cJpKeiWirQ6DQM0apmsotS4gUvLU3vmZtPmPl8pmMP11ggAv9P37RgpqUaKt
j64TXKdfgw3Q/vkKtnyqHl4j8xB/wxrNSeMzk3qcBU9X4gR+b8et+NINg6OBHyOW
bqPl3VP5kuT5F+I0Xpchx1H1mlrXsB2c0c171nMuLaRIVaA6WKcfr6MsQCjtPHtn
EbkpArI42+iNdTwXYkKdYtbel1qK4rNCHd2QDTcw/h46rw3hY4ubuBxe8PLHTsYe
XKKj6hzxLm0tQdnM2cuXY0Gvy9L9JzvMBWYlJbyZAIjtCPWhl9uf1o+9dcgJihDZ
CgU+U46zMNIGnBqLgPzifArG/fQWh+t/lkGYHxVS7uY/hfnPsQ2PB1FnPUwjsqPv
K0GjWd3EX+GgU/8/TbjKoyArEBVE5C8IRw60/dT5GRTbb9/CTpvHobid2pOQ8ONV
gpCHL3PgodoCRWI6wd3KApwRF6wj9j7LDfWh6TwKERDFMH84gFBMvINBj8Vd5fHU
dtv47d4Y++qjq6ABMu9rzsx/Opu6ZvaCfZ8/5Ji9QpG0cuABpbWLe4rcq2N0feLY
KR8egVE/utpSFwEZaKmdb0VGOTjajXZj/LWik8lObmxYXuKsGgBvK4NFVWW4eDRf
1pQzR6cUk6Kp0b0ZU0ISrrjue+olzlqh1Knh7v2VdLzo8e+7lJe/ESuJErKyfsO7
erAwxjKU7dqP0QmY/Fm+Ubza0VHX2N0zb09OFJgja1/I86HHSaB5hHdmK1eevKNq
mw6iNTa0e+9NdrJDveyeQnd6NEgoOjsXK/Jz6/vXZLqH9y//0GfVOH8pxVuFuyva
lKZriCpUZOBH1KcvJ19pMaOZbOjVOXJo1bBrrsvw4neZGwV0MAsV2byh3TJo/gcv
hIegZlzKVy0zL/H8KZdp537mdySPygRacU9dJxKX5aWC4Zb7M8+gVY/av30W06hR
b5X0MIpkZZzWLpK47D4HJmYWycqFyTIQtfwY+r2krqglQzfrxoKiT//WuQPYv46/
BCSY68I0x9CuEZFYyMRSIk13g4WKCfTm+agKbL+4FMOKzBYXq/mQmOGMBV7MZM2h
yp6sOsTPqAbH7EYWyAqZ0m9DFRyHXo04qhKoK4Kt3ApV4VEi3B0bwPSmITxaUFtz
L5/EimNI9IaG+OJbzVO8SjEYCa/5GI5GN7+0ZzWMFtwi8ymCoSrGMb/v4SsLg8Vp
rS42gWGNbtfqhFe05ntfe14YDeUtPngTLTqHkCbgD16a+i0+cdYId5v2Vv3xI6l4
HczfCBqvCTZisczJQGjdN8Egr67I/vktDDUL5T76APnheoeJJpOFkjKB/Fqhkke+
55lQwF+d+XEPo0HxggUJUsdzz7ocV/csIuO900u/Fy3oDXA1lQTsEKLkotsmyhck
wW3G4sGzUYfqO1Auu8G8lGz3mT0Jh1sib4kFVFZGUlYYMtmxs7P+MnQGfdl5QWS3
CC1AUy05YGJSBHou+GJsxrg4OJerBxla46le3I5n7wnrtvzDxNlALDi8Iq8WzIOP
MMm9gNQjDzh7rEPdjcE3fqZl3ZwGIakZDLHiBw5usQHVHwM6t2Xv47c+AbXMw6gu
dIjIEQXJxcwr5XAKHw1v3ht6ycE0ZeaxVueCe3zG9Zc6BB6pOMB4WDJ/gCR8ANQu
/Mj2Vtk2y8l1GPaYEcqz7NCWpT1nkwrHI8xU8q2ow2hUEbD//ptzrjW1YQ3MetYG
024OU9+c+6pLtV9W3FP7kapkNHgiP7RnXjD1ZP7p2arRqD4zJBeUjCtFMtFF7HwK
oiliOVzbwOE31/2V3QyI8lJuZGx3myWBaS5OAPX0PApxlVBSQNoG3WLqVcyQSROT
+wF2XGZDbMGlmyq7QPK/FGogbxhtPpgqilFuTmByQVEv0RmLjUaAiQsMJYdN2HQq
DoXLDfxpboNZlQU+vc4XHaTVpDU51s/UTkaMxVZluhuzHMByphMX9JnChFDbLd3p
2OfHDWGvHjFohTgobkgXR3Om575FZE4L5AurhTLog9UDH0IiADRdqaz9DW81E6QV
VD4PLW2W8j+x/UO4siNfyWM5rVkNcTQB0ogHpflabzyqlARSp1V1pIBm4eJvcYNJ
/HBsKLS/p3n9J6tZctLESpcLktybWGDF6ng5YPsrvivYdmnMX1A+Gnmsncsa8qvm
3rLETYuyGdXbQYTrYeyHzLnIn77Ssye9IJRdFQMAh/sxac96WQR+AaSEEW0+CGVF
erP8QoKHzN8Cii/GzpEIehTaEJMxjtmiVmSqmli9iVAgQ0da0Y8yuHWRVJEsGHL3
pas2zZnfmRsnytCyagjY89mjbUIKcdj3F1BuK8Hac1QISQm26+XTlIwxJm9G6Sdh
2QFLe+vZB499GSr95/iQOK1qvLBwWVqQmQG3M2RcaH99JRhACgp+a1bBUk8QIbGU
LCJD13nMV0lg+m54dntUGGOX/aXLUE9biLzb31LZSLuhBQzjqAafiSRxmg7YagVT
1QMlJ3Fj0oL0CiGquOs8J+br+pH/GeRsA2He/de8aQG27NfY8nqUsmyzmJKYbzeI
VQkL0MQdo28XfbMcR9WqWHx/aFhwvJ4hVRmuLE3wUYFerNQcOd65FngjNXw2YUO8
NygyS/p/IlmO9JeeOUbZARj68NdC6PokcgVAk22LoZXqQcE/q/1IdlGLL8s38/DA
kGF5hHmDABVT4UDhPgKdhSOhKJ+6zJgan1c09rpVdoiWbtUzPHc1+vdnVRDidOIL
mTPd3orYI3YhATCpvDvX/sjYdyTtTEVgfYvp7u7K6e0hONSzqyUzj8cyz+UWGIw8
ssfhhkdCfI1bMWcyl4JYBVtdzVqPO/77cYNmx3ATzYVb9Rl9lb5mFqRwdObdO8Rx
3jV75FUdUICy69BsPOvZqZtLZLlT08HvS7jcruc6koHjRAtRXsKKtF5sMAgKmOQB
Ugvqhun27BTS1x/JCTkJdF9jYSysInn2WGhR/KeI32AeyQLg+UC5U7LB5fdR/0K/
wHACizFHVAmA+186N3MgPkW5Y0HTJhNLECY5ADP7aEUKKmcLXosGidcEUiXHYf9w
ahbsZJ5CTRQhFUOo8tN0oEgcngUMFH9O6DQO5VVH1eQoyRN/LKAVyTQqqrAgAPRe
3AgYdUDgd5AY4B0oHfnDy+ynbATHzmIj4Lz+xXVWwTbq3zowQkEBEoJwGimO6CmV
YFHby6QpeBShaXGICpZ6/m2HpNjPwF9uzLYQWx8m8izftCdjD5e4WUoASjcRkDtC
IMV7ggyH7gP6pBUIHkxTSdCOnt4XzUDCU5VakV6joPfKuVVn+sDc+pl6y04tt0l0
HOogFbqwEX4qgabO1IANCffDIVoIRbrhvFWYKHeBtzWsoXG18gh4WR9QajpOwy4p
TtS3mHHhKswPoCXHq0kuGDLK+HD47Lixr3X6iJ0ZZ7MM4Rebmc10uD75DfDptzVO
YTBYKE2xdVUbh1NSKrvwzQuCcCTQ/IxGGJuwjw9DiZt9OXFJ59i6m6Y7vK/bZ3WY
Y1krh5YVfx01zHUYba3bm5MUC+h0W/PdondCE0DKDVCehY2/g0ld1aoCqPGKwB3h
mjy5pN4Xxn3iyYfEAXk/vZsXnLqP1hpmUPgQQ5+K8UwUkWDhq3J8JzjQrpDNsfEq
FUbzVTA35+ASq9KHnJmhZZO/FtiiRwF56dUSxLhXJT3PEyiGLaqrh3FJ/KQDnkvN
tCp5HJsvfV32drPVmIr4fpXAbGb4Df1AD9/d9phVIaay2ZkDiORAv/91q4fL+aFj
51kTMzRy8VCg5PgFgEsJSJpa0U/23xwUkq6fYR0sppLVCN6+vXbiebOA/qQXVvlW
g3VVCc7XY2/cUofK7sWomLIPh2r7zE2aqbi/EyXeLIoph+YcjAnGPsYXnishL9Ju
lG9LL0JzjOyM4k64dpp4mUZZTpYgyf3QobHZqgxqytKSrV5SiZ8J748dsHPq7oK6
pLdZEZW4RqyFD1rPfJcn/0VE6RSWaP6IGpCQshMQQCM1Qh47HO4zsW1BD/BrmoKr
Y9MccfGcL0654OsyrKsao7EvBmq+eJYDjDfERfs1i6eTiQsOOOgR2tJ8GEkug98A
bxUmnqKPr8FOsi7NRW5G6PndHlK1NG6yRP9wn5DDDzGZ0Oap3qbsznIhticXty3n
pz/HYeceBPTUV+kS7bTSTZI1pfXqGbO20OFwdeEBjUlIlDSc+Sq+5v/cxe+n2aAx
Qndu3RTQeRThD+PdqdSqsQu8gmpFY0i/yWFbt8GwOCaz8x4KLIrzch6sFK7ElhLt
p8/EdP/L9kx9Um6U1saWDYh32pF3P/rB0SxtOoS/wHVLVh/a5jh0nuawjJfjpAn6
tOdtSqhFdu/Y5Qam7/+ULiZpV14zChTfMDyChO/rvvZrJbLm/7qFPLG8dGwDPEDp
mU6w0nTa0MB+3wYrAl1RYvaERwfQNs7pGpx82hx+brLBbmbzzCqIFdvA6W4DjfVi
moZRX0VQjASDOLAWMnHcUylUaH6sEgbPomvT/YatY3OZp9JeLIbKE/RIZln1W2CO
ByFpg7vwZrEoJuJwlZxXxTlZ0iPP6aLiEhFFwicKzWsDRqOBKR+T3HvepfpUlpLO
0/eI0T6LdihlZzHqh3/XTmK79JksIYfbWpq4sR4raxfrsGx7W8ubKIDJqdl+YmaU
L/z46ZMgvGZ8nm4UJZWtGEVYKJ/S5b5re56Cteg65nahezKZE5rfPF1iqDX/kmWY
CV2N26hyyC31LnZuDbNXsWW6YWGe4TQFf1OAC047jzE9Nq1DdrSW0019rjqt5Neh
jBtn7KLx6zc+kKzXWCiK9WpgilWdM0FCdvJffanRcyksDx8FgrYjYvrQkId5Gz63
69khDwNKDv4fEJnwwGuovGGRLXlXYVyISOtooNFe9MzUXoUqq/g6VjpZldF5svQR
M2LCDkLVSMWamP3lixnDhHve/oOHYfmtqoqat+cCsl+vULy6lyZeEd++Ld81h+2r
Ga/CE2r9/8F690tRBG+IwODjSygIfsOH3eUKYufiQE4AfBVaIicrt48XEs3Jc74K
a+b10eqrjxxS+yq8PTZMJwVEsHDZu47Lx/qoid0XdoQSwG8/yrP3x1Ed/BZ98fQe
DBFQkJ05JwHNtY+qoCCDjHNcNzltw9QfxI5mmGHZtTWxHDuvR6DkSZFdh4VTEd6i
0H6bLeqOonCSmq5OUxXpHYjqn/Jw+o5c8V8YQmzUt7h/IxyNh9GYTOEqYr2f9aDQ
kAd+uYYd7/JEPBMJfxx/QKF5u9lupGh4O1zy3E9U6A7ruyrXuzW/xIqdNNQGgEuW
9/gQJ9vQJh0rzfgRKjnSfqsTj0wQrx0rScM+P+n6+v0=
`protect END_PROTECTED

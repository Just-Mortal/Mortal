`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nI7LBSQsuc6GrzT67pYNRFx6ffxM8a63cirR6UXXKj0Vz4X+y/NLICDSp8iX1LSc
DJUUQZvwuy+mQYAz+f4mvAc/snX+YnPkw5wyKvlfZsA+D3oMtGjbUn0iTjXtDICZ
LNkzTVOTIW60+FozvLYvL8v0rjGcq07nXOVfCOCAJU4QEqMjE+VBxUmYYZx5Ygwy
ByCJhRbBCHQQAX0bAyGbE9MSvXkXIA8E4ST56ueRnb0btFrN+oS7dEyKgWwHO5tp
a8Hq1nBez93SGQ3lB9zhSUUevVWqR4oLpjf8V/A61/etTssBdVWfzDdcBXGJbHtx
VpJqFMquVAN8E9xSYqCoUc64zTHfGvXYA4dPmq+7gaPFRcTR2vfkvekJ+Mq6Qh10
6wqxDu9Tc1ybu7en1WFbxKlO+yPBRvctaQb/BTopWZOPHOfDYYyeY9G5H7myijfR
vloYuNaYbm32G4EgzuKOCKXyANFRmZwjfxc9PYS7CFnboFSdXzOFdjB8XMXia4W3
Kmk+0DNCxfSpSIEaOtFnRzRN6KPu9wqeHwSxf9Ta4qcsT4nQFpo4MkIGfE1RNjtF
SE3T26gmxy+3c79TF09tPAalnSw6mHatqxapFK65b43HGbbj1Rt7tQdgdXJm/tjP
ihO6mZvZcn7Vw0rC6KcVfJdijMUwhTd9HqSYcvoJ+aho2Ygu4rTt++BabFbyI8Zu
duEJtJYwbY/CSh4sZBH8/ZhX3ynyKdZEFWBAN6sHczGPYPk5NCb1OzoO88LW5E2a
ikvDaNMKbDIgOcqAUi23vwMfR6dVGNBqULwK57wpGZRhPfGgEo8pQiJD9KV9+rGF
csNANsQQigkpiEz5BqUgYlZGIYUN7Lxl+e+0dt6f/QK4/ul1eJt7B/gGKZnHuA9j
SOiXwKW/OMZWEX6X/KshkYN34AhpFhLJPvZBlGMs5JMnHmkZb48UpjG6+3mRbwEI
b7EgXf7CrrHSu1XFykOTlPGkMhABXhEvuwS7EJiSy4vniCqUIIS2d5I3Spx3Fgmd
suewQObzDg4zPz00l+mY6MSfGiclkV4z+UlSRn03EOWEm75vqQ6rRrq9/qe26Hae
Z6rJTt09+gqex9rm6uUBEpECWkGHAyKOZb7n9SUsgMiaf/AVEc4cXkyobuA7R7XN
QF9mab5eySqhBMaMAQ8MMdeIgavw19M8XxS0oC7wQgrbCEsz1tHSKMgi3s0hTO7c
bJ6WzN0ZxYEoREe20UfQH5sZOHVktJcwDCpS+HupcrFAfKcWNFdrlt9yN0No+l5H
lKHFEBy35ArSehWJ+DHsuXDfGg6Vg8b3l5f/7sMjLxIvx3bm6RkxHvG5QT3CGXLQ
ky4mJ5iCk9N5jlzOL5RfkPjxQ8X+tV5Tok0qDyt8FC4SwRo4eIHdqZ869pWCm3w2
c6DHs1TGl/sYZYm+/hRsD2lrLbBNHkWXxqhSAynSqmTw4bfDWuso50pZDNQYvjLT
Z/GOzOrF98XkpUJ6FyLpsj6YLfICTVEeHcZoffXyLR/9qnvIA6R2q/MEu9G7bdza
62516u9jzgnd8CWoqyBZRIJqiRSeTQpiXph89yYLiicn1os74Vf8XN9QRRUJXCPr
G8+0PRuCDmTX+3bWpveXdQZ6VLMQzTc8pIp7AGlLubTCdfrgDKLtauafRK1CriLL
RWhW/rZAoA6lsHYXxbGBFWGcdeuXT8WTawIoTxm4WHJPvSPoR+PDyXSj4FbxqYHx
AbjXRE0djWnz4RbM08yUhzzOoPH2YT5k8bz33MoYHLjmO/WOZE+1K8RlFJcUpa4t
eYgFO6rqmT6UvmMM3g5FBKPjePxnlz0vdLIiq3oZM5BcFBbcpd0VjKZ5JRqMpiBV
4sFzLU4HT7ckK6ZlcAF3N/xR0AwEsB8o6M7UFIfVnIcQZ4ZQFPo/V9BHv/v/Ae3f
2aIF1WGEZobeoP2Aq4XAIVOAdNQRed6odTnD0mO5CFpx2RIZWnu3lvrezRd10upe
hvqfQY1CE74c31d8XEH8CZnHRgRiPcAA+G+Rp1vSqv3juvJ4kJoFUy8YHWtFjszi
ngFv1q23d0r76lsgd2KIu9scDthTkLT5yVLWLZZVqup5HvSltPgtY7349pq/OGn1
aT6NtFPHkVaHbGDsUmnfuQlQg8VjcotP2jVGsPpSA891+i9BjkReaLsY0xJ/tCaP
cIpMFYEm9+4/I7PtTGBisfVduMh3zvitYKh2270aktxJoGMZ65vjx5ajCoivKv37
Q81mdqt6tS7ej3JCbZoLI8WGiWc5DyOhShU606crXHyixPqhV/yaqsDXhtF1asRs
BgJbKDQny1NLTmFecMrRwjEsJ7IwY8BVIv1NMI52wvxgD2n/h3qd4/5H22uP6T5O
xfz7HYDaUyDZt/4Z3PNnX+UEN/63atDATH0qC38JASkr8g6EmBLcqzFk0eEFEtNu
a+Q15nex74dseXhTLqYlBQ==
`protect END_PROTECTED

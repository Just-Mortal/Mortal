`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iG2/aLvqFudD1YtysDo4Bx+4GINHnmmM4c5SgaXtGPivV7XvyvXbSH1gCpfR1Hcn
hvtYOo1WXBphctpJzuBc/s/HZJ6TLWQ2OyKSL4rAYq3/WbnPP6KFgKyxIc02aaE7
8ETymCwoYkrxvbi9NYla4+tzVPjAzRGZoNpcd3lzX4ubH5TDZyWNwgpWRF2jj+Xl
RH0LoKePmDOYJbidZHsqYocGmuN5BxObP/8LwUdOeh7dzQTsIxhEPUhuKkElZEeh
5sO97DmuKqtmJrLClLMvdLZllSed2GbDZyKUkIy2H7y/q8sXvOvjfDQ+7sBQdDPu
09Ctl0OX/mdvT3/kPCL2fiYiMeqpou6j29VvoI09WjhZmwcROnslAT73mLuD8l+U
/lFlLTqfXsst8CnoSmZz2W8JxV+mJtqVkbjn/zFqIZhlJqtTD7XfhAbZ7ozmqpd3
vqv95NCOvY3eg7k26ios6wNqxEqxzH55QqugvVdSpxS5CcSjDNHdWgzrh+5DncfY
vba7Vmf5K9ljK+mlVs+Rs8j4nVv8DM1dk1LUTHfbayj7XPF+U3UsKJCPJd/3ZGga
jeDtr2GxwxmtQt9cbxAn/7G7Mz9uljYFHFa6uvNnAFB4Cbukpo3LE9nLcYwPiJca
+qvkCvUyufJLG/23nqOAlIIBpbFSrsCEQ73p9MNqoFujfgithgvORZqPCGsoDRLm
tUOxPXscuZFhHj088INjxwFeSxm3RKUjnqCUNyv5+aVJqccL65ZMT8JJR88CJMDY
sozBXDPM09gEGZsTkv+e6GXgzZf88730bcgmF064DsHyHg/55tytBj2zEwedijbv
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9cR3JtpMWIhNSBPtA/NQrTiL41BZ55gjHmM3JKlVGk9284LIfqJmJBqecH4+LrW
Skg8b/PctCSrCV3XUcQwiS2S9PSTzurs0YzVWmM4yMVXQ0sAufwY1VyIGP4v4zea
81y35V9XfciYbOJ8h6CwUsbEDiPBm9msxpgYJFEyjdVLVmMsr0YGezKtv0QnSsIe
JFoxo9R0KrvqDJI9aala1ybHp6Zh1ZR0ZqWT4FcdgLZBa9R5r0qmcFWbc0OihPhb
1jAYayPmemdpiWbZsp7gTzmeYtuolguYk6EQPGw+Vn5/ymK1DjoT1MOfzN6cch+a
YKcEDeJSPoDzxWancHSlOhcDqTk1o4amgfl4bTyVND/4+thc09qSJERrRIy/ZP+R
KlXnoltICEZA8A3I46GwqKihp7kDwd+KKhSZ3tJpl+4/qA5TTDoH6Ig2rKdeFEl1
gjqIBL8GEmDVHESx/d0oq6FZw9tq/zWE6xRExpyTPmu5v3Nul8VxEUKLLCyq3zZO
H4W+rudna/QXL3E6pQt1ZIy08C8qt5frcTYYoLWRQ0KOCvZhESyjvDE1IdJE3VaA
/GMOfxuJOovr45j4ac3GNhfSH43817aDzKmQkkMOX+JvRfQLIgAWiDloUA5Z9gXX
fKASrtj0ykt6Z7gGxi7kvibe2f7KhAZNo1d1psLhBUzbD4Y3e49otdko6HoifVht
v/u+HM7bzqJvTghwozgxCmwAqJ3e6bYuYDA0QlZ9k+XZocC20DpRTAr78s8cjvXj
7tloQWKFQNz/K0wTzt9kQkC/Bn2tbSnFz3CVy0VeM2kpWub/pCvll20sWamoCJWr
ddGz0JW7A68eg4U2t7DEJrN/SXL610PpD02d4E9x394JGeZ4CHBs9/RQS8VTWafr
YPdfTL7dvSa6VepExZKBkxuOLGupI/Wn0GtSFbHhL8C1gCvcVKH+GDUeRkgTgicf
YwJJ6OwOl4r71rlrTEJQJJAKt80QeIP5cR6m2SmRHV9KPETxc829kJ247NKzdFY0
QJ+BIyAYX3ynLMK0Y4e+o/7PgKrS3FVbMRV2gpyQ0aRYG+xiMJQZMxt2ff/6CeNP
nryxnFgosL1fbx6PMAMx0tQzgu/xwpsrebUovpZfNcQsMWFrcokVkMfMCIO1QxN8
VhUGmT0yCS+b7mlbIYIlmnFKN3Bm8yTm0kqFdfb9TWMjuBpczrsc5S5cP610dP1R
5GqBrpnFDZed+tHg4vN/FyDZ43/8CS7/OUNM2gAW7bNt3zceCyPvKH6TcIG1DEPp
OOTzSj/ibo4T7FSF5EE/BrvoW4rmMBn/5mol0qbg4QMMn+lNHlDGaxf9n3ec+YuW
3VXpuxNc6kXXotLrUgDHfxAkYaKZsMY0nlQaqIf/AoDizMWiz6QZ4xBvBrqgPb0/
+TQMh0e3FAEHFeItOBGqqOzjI8HAX22fgAw1YlXaTJJ8iWwydZv7StkuZPmUD4B2
vnCV2K8ON/FGJuXhpIvCYjLYJeuZXlF6PUjIgltbbLb5OS2mJ95Ogh79um6odItF
nAy5T+XLhXqtX/aMDWw2hUQ6JBf/u1HtzyCz8vzJc3i3YNGTxLZG4zlUGoBUCpXS
TS510QZhCt7yYwCE5JSXb+KOVCmz+0gG/qOaHzgqEf93tqdad0FsHPkvj3PmUVnx
LGqpt40yO6PZ2pefR4biyb95QmHg0ayu3FXJYHtP2ODUo45oyleCXRFaOBzoX1iR
jSJ0Bj3sKAR33iacZOYOcmQ/JeUERDBrRTyo8umtsm+mBrTj0hfd0tLhmN8gM8xK
fT+sdHX2aYfwEJMMoiuup2P+Cc2kAmeF9Er8FsqGy4cMh8DL+gVD1Oh+SqmsHBYu
KnyLzIdKeyY7Ll3mOTsA0fcVM33NcCk4y0y4UKhgxLspZr3nSKo+96jC3tHzvSzO
FZQ7Y9Sz6+uE9FbL1k/IQdIiCtP4579V+umGi0bHGpOokwL/wZFQ2QUNk09Daz4g
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ecluyvAzON8rzFGHKeCSxnCSig8zOedw/pOzq00Q5hzXplpR3Qyhm/XW4liJrOSS
bpcgqE+mSihfmLHZeJzBP95QnIB0k7SSK9cTjWISdJOQlSxYA0KKBYrBAfTchUiw
JW0KdPIbq9vFjB5v4gpq9hUqsy10HMCbEjbEhMdCIyHRz7qmNxnemJOdCehomrKe
Xmo0ABk80A2/8Ny3c4BDYvxG3eDtSyEZW7Qu1du9PvxV8a9mSXJiH9RhUSx3xqbk
EDfdeZRrjr585ETQHAuvy8e64vt0R7KHplcK0EVpiwdGBZ0ys/OcLkdrR/uqhYgg
2rYGNbdemtCW/7u1JBZ21yUzXprZ6yVgiSasXPvAhv4aqIoeTLwSosyQsIWqywkO
CKlXSqYVtDznm2FrE0Red/E7j0q+Zx8Pt+VkaGwRJ3b68pi3HJPSnTm+xd1VvCfZ
eq+zLYkN8XT87xCZdZ7q741QW3U0IYExJ1kI4wreNHj8U/zfpX896mB7Ma5ZhcP6
NvtcoUUPMQrWh0P00Bl9VdhtIqxFcxGP8xrR7YcTWWLPKR1ZfrNZWFrC47ec3sPN
ZYEHkLHkZTRC9oFFt3aoEJ04MCdK/evlZ9OkEyCN8FQVHKuxJodZPHUf2IP1KNR2
G8th+ll1u6r9pGSZwIoYe+AWxYm9iBUgM2dVBTqu/zyN8TfrsN0oyb2+O/4/+eAU
BpnBzb1QNjuao7gJG7+qVL+m9+LbO1VScBbjp9NJked2Vf40Kvs4QWcPBBxx7TD1
cTpZTjESkBjK9/eJIrYzac+V+7PbGfs8g+Az0ky9vtozzb9ngaaKCcP+8B7z7dns
TlDJEw/xjiysiThvIu+YPgZHAvSW+OuVGKxjGRc64jVD57ys3+LrHfJBNy/c+KeI
2YGo67c+Ks4HxEP3Um04YHyuIgeS6/2Lennq4PpxopLsUHCWsJQHN8m7qcPCy8IM
FMg3abkcWQNBgJkFf5xGMY3boKbL9kbZGzQc28YsV3gt2j9B7hcBBfvyg1tYSNmD
iDO78/18m2wdFJ3l9KB6onLYLbNvJH8IOnk1aErXbjZP2t0ye1xEY9glZOcI7b3s
Fx2/vAD6gXBywfZY3A9A9QSuEJYDjYMEGUbxXMgP24YLOeLLeefaBiqkanaTIHlF
/pAW86M9f3NPn/CJWXf0B8fHC60f8lzAR1aIGA0YGHfLFWFpp476kwAVf/2o2cLQ
t3qXevPD+VqozZo2r+2Y4x1u381CjVF6U8oLEcdltpFKzw9dqFLK+UDdUqL7krM1
Afzd4UhaGkgql9iumP6wTN799/oUAvQTxiI9/JIkrLnG47pOcBw1P8OqwWYB9z1H
rKotGS0s7+tgRGEOHqHn9NO6mXnhmKz/VFe4Awho9wu9oosZngxNMvz4foPyXxtR
/9+EVXE7XF5odcxo5cweJH86i2eHdbUrPZEPi63pdzJ8mzhB8dpAHRxaeVTGUTWZ
Y6Pg3rEW0L1+/rCpcmL1pzz+lV5liw48i9iWRpYJ9S16ugIaLDMb/eviocuMZHr3
L/nyJRROSwNgl/DRIB3ikSjf6X8ME+VDq0/Faaag3phREhu+FuHST7snnPgEtxi0
IcJlHWUx4mL6sqIZd6g42Xv8odTfSfWo4iYH+9HjNmHhBdMDzLfLyGuhfcfXZ1Bt
dHtwcZhb88+kMK1GuBXRT0Yu/KEDyijS119mrBcjUO2jJ9tOpjMs2fJ/uvuMMBB7
YMaO3RjKpSwn2RcTzruDJRYoWBYhVUH9y2qGe+vsMRBXQwwe1uRdFSsdvGdK++gU
GKDCShTDLlE4zcQQJiG3y5we56hDv5SZ6vcY21maik2YKzvF764ftT0KqYdPteei
+kpWrPbJ3FE8Ee6yCfo0mNOLeDPdQV7xwVITIJpK6Gi06vfewUuYOMRQosIzHwUm
YF0eSxqTJGaxqv0h+teck7vxhx78LIzU5zEIcw/yktXIBTskXpMzlaOnRVaQcTbe
QPv5UvW1ah5UL3B91jXc0c6c7e/EEJfgNUSjtMaPfER3z3s1axakJSjuA3M5R1xP
nH3xkIuOFZ9upcrzDZEvnDt/7HA39oHbm+gO1T4hOG85RxWXjuXd6MSZZX/2NVHe
I3s95eVo5auVieBS3SxLMUPLrQerZuqKgdoEZXZNBDYp2AIDtJoFinoE/GSdwwTW
H6uu6b8LZbct9TO/yakP93BaHnuGBgUzsOJKM28WEgV4YTDQQAi1h+bHUVLVtce+
uCDkX30178Yc6pFhL90Bbk6fdMBkQ3lBKrbZ/umSEcqdxbSrdUOmB0vQTTvsmiGZ
/+HYtcTw/ahXclX1LS1IkkfRrw2YRaBd0jTmVuOEvwySnfd1gHmtWCpYVbm0Ctk1
AvxULYZhSTZs3EE8cP9DD+CSM26QfhMhrsfXb5USI7krwjcNt3SW7vdmIxh9HMGV
p6gEuRyoL+ILolMQ4EW/mzpbGrS5L/il1Svisg2UlvjsApQLc9eyB/XmplZF314s
n/EYBtNG2tOINut53BUpQgwmzYjLg9wQTwNfA8JFrut9qlqZ8pAaxlOe5Ea+SwY2
kTaTdGrx4gz4xtW4AU5oNK6BmMf2y869FioXNJXEAKng6nlscptQwP7JmF8OZVW8
rwXbqaS8dnbsRPPaUwAyhm+towYpsJo2m6Wa+1PkCoHLR89Xmn6kaNLRcml9rp/m
pzX139TwUGeBnN5+85+j/kte1OyCurBil0/Yh6E46zsXMbnykCGL/jKj7MqaaC+9
tcrfdcVEDHLSG2Ll9d5v6z1D1ynZmKzugU7nbgNDNv9SpAeRFAkmXKECzo90u5kh
sl6nr7Y35rtcrV58JrLahKoIGa4aW3VLTut8RP82gSlnd5tXVQzICmpt+XvytVsb
mqImY1qbiWuiTqtiar7mokP8Sn/cEvtU+8J8V9+BUF3UslvCt9gmIQ45X9BSLFIH
yAjPvzLzwfFlrkaYUz8hcvV2TAFmu+sZWzQjaDFMDlL0pfRLbUj+qFDM3lfFDpVQ
LAd70xM8YiTV8uq3Kxiw4u514ZaMrFZ3RlRui6ujMh37utVzJhRg29RnK7l6CQfc
xZqobPT1iCwH4f2NA8Ar2ju0rzlHsGrW5n5PUrRWVJ6nd9pfPV4K9GK8S8GoUcRv
AC7ZVgjY/a4I3hsC6zxCP5boFo3hqhcH9esAZO++/Mg5/FJ5EU6JKYKLgvXtOGw2
VmNTEe5c6anDf6j5D3zEMShEAc2EhB7ia9AMBil16fl+Ovky5tRDnxc8zEJxhMh6
/e8SngNBC2ggruxFOv+Tv1QmkdcC3v91ex4cwpekQP0qXHDx/wgWZXcSFLYtkCBM
UmtgKsgOMqVxcMi7BXjpCtD9ihywCmNkH1oQhH0MfLSWEpGEUyiICNGnrTdPDBtX
TjcqUXraL0d8q+cY8ocQW+tlmIjXZ5HPsID7pKJy4s7VRfFJcZzbZZplv2SiC0p1
0rtlZ7iq9RTTrU5Gq2+pD74dwgkHzMVlVykqATVwwOOEwc7RNbS+YPzrQy2rRcqd
XBBFaf2yY2oBAwuL8oRahL5HC9/PZ0WmYNprIP0bN/NEFHQLfv5bKrZK0DDf6FiQ
B4ViIOcISyINgmrNERWlAJfPAGVoXbd76wbQ5rcHFX8FDWlaYI5NEli5baHp0P9U
8dYtIqHHxAtLTwqS1+VFHEa28SkZOH0In9M0ANw7Pe5gmc5iZJfmMWqF7CK4Rqjq
c0j78iWLdzWfwvH+VrKVnBmtjE9tScp1PstxCMtwcZQvMEbaMaFgyYtPOFYQGc1e
UXHRIDpq02Mm6WStBzBPFq/P+dc9WsqE5ooHim/79ID+pBEGaogGis4WIfZ2mQX4
0wHKzI1whL4lPSR+w56T3vjzF0g3thaV02YLhcu23syhJsrW06vQGhAGfl61j2s3
2JWNuJhhIoNxndC5IyRpoSmZ+oiGxBAPRAaNNgUUebX281aMYss6X9KGqTZkMkVA
j20MQ03S6ViH9fLstvzU28wfinmYoFIQ8CwkATrE4R7kyiIlpV9QUvISn8gmUB8R
TwD1e0agmbH7IqvwzbY8RsKz3BK/WWCbQJw5A358BIG9mIseFQ42wjnFFNwGKQ8C
AR3NmG0StS/35gZEDFBa641RuPC4Pdhu98fSQqTEFbjFPIJLPTdMRFoTWT2UblYl
AgQibWuSOpGCWSsSRc4IKer4h1EQx4AL0EUVy53iRvMg4fHJH+Yt+v/uhcgvQn+u
1HX7c+2JOxDFeL6VC67lT2mrq+rlMebPozGGD3uUs/b8tTZ4pegWIhpck47u5WYa
NfOnZzqD91Ji826MJToICL9EHWj3VGchqfNyoOMKCy6sbDaFzXiVL5QkGE9UNYXB
lxYvdooMR5/ugP/CzuQasx/BCltG5hkBUeNe9pYZlitiXAvIyOua+2QgZdnP3R9U
lxh5TXj9PUEkBmZg8hep8b+thZmYx+3HVb8WQZ1JQXoyXZA2LZ3ScFD2Z7HeMWaV
PxI8iPN95q3Sg4I8+MGIPZ4xa+IEB0L0k54kMzA5G91Kbrih2oedQ6hk8B8sGK/r
eiMIOwwrGq+ir69w7AClP5lrE1XFA6GKXNGUNxvIiKHIT6ViXMbyeDMNYbROaFC6
+0wnNACzSm9I/pouC4AVi5h0UwQNyuXuOsq9e5wBsju1nV68HG2vvuevcaWehE3o
rG/zXrJ8TLC9oUztzz9DuNLhR/rsOaa8AwYEvujSh3B8vGiFNnxoLqxmReH3wrpN
W6KV9MoiTPzfADMfoZw2igzXfw2OwNLD9N1TahzP8H+TsKHyf49R7v0ZWKa2LiVW
JnJCjM0B/HLHPJ+tGCm/u57BGa24vbcwBSHkhY4KAPXfqnkfBUJpMfepHx/ONquL
k4yn4a9SJKKt4igCPI4BF5SaLCr8dw3vr6w018XYcedpsTZy9EHUA837588JPpUP
4KfrZh9Dd6CbYDO5VLhlTneUfqVA2HF1bAQ3Y6NOHz4/6eLtX3m2NF9JuhUrVqrS
WcLQM0oSLQFNpCQiypXTxcO2GZwvt+DnbO0RumH+4S1WGjuebYEOcFT8QG8v1Wfn
NUluaDxd3NibrsjlEkzbFi2iOEHnWTjP2nW408EvZPJPGOHgcPAvyr9rV+Fri6W1
zY92UrRMNH4PCXsN7LzmI87ETGQpy+VN5hLI2FXIAgyPBMZkVp8u031PIVSeJgJR
llnr6zObBGpbzfNbZ2ZzDE8PFD1n/pb7ie9QuX44N5zqKu01FJqgtV1xX608bGuI
ExFuoxEkw+xlOrRHqKtVOVYhh9ns7qcJ4dZWHClkyaH2g44a5DxQCrL3OG9G6A7k
dR/gZwJSPYSI+jrrGWZnZ3lXE1IC8lEYLsSu8TGODtMH8N18/C5sdikGNk1kXtZ3
GyOGR5vEcZCdEbiAvME/Aa5QrVY4kQk8o3q4AkFtLXDnNHL1qPS7t+TR0ihgg5sN
gJL051fJCrDn+V8jF6JuGcnqbBt0rDQUoEEBrXG4lftc2VyqjS68oAQ0qFjborNJ
jtAsfHj5rmVi+cuIFjSAA55vrhbrZF5yRD+17X/pjBUBT/3UDllGCUywOM50qQM3
uF/dYKGmxJ/krcUmHzB0IZgaypA/GDOoWET1Q7IuQa/+eyjCPB2ORvNfhbIgXSsY
pBgOV1HjDwgwJ48adaIFkJ4JBcIrJosVuQQ9sc/1uumyYKyRtwNfYv726FcYQB78
QV4w7PUkD5ThGECz83V4mNeAlZ+AyS6PwHW9+5IaxvEKwi/qcSNZD0+YIl3emCm6
3fZhVIKF9NyUu+6loUD4zH2XhNGWx/xfmc5O+UTcywtkm1T15VVcs9i7CmqNYo5e
bFBHK4FW8VNZLmM5MF9jmE80487CVQzw/Z7J7NRHeRk5o+rM+hC1/u+SphGkgk0F
k83Dz9uQmcR1lfqYTTG0bu/6JN0SMyS296isFe8CJIamCk157jSn82/1v6HHK+MM
m5vDZLEVPgcPzX8fZReGQQkyVeoTGCZteIOO4N31pRmwOd+HwaTl5MgPFqSWw2yk
/ceNi5Ousw/8fe225W3V7t+SaTP3u7Y1/m8Rf3/IfpH77nn+8+JJPygh5tXp4wCf
eNYTkVuUoEei+wRWtmgGleLpFgqmDem5Cm6i0277xjS1U2OuxnhUX3jufLH5x6hd
gszMOvDSv9TkW7gOrQv40Ul5yP28O8Qw/ePm3QNN8A787nlej79WhN+WjX1utCaq
xCpNQbjWYWHOmKJYWI5dPX4wSS0W8NN+VrZWRbXWcMopcpKInGSqSxpq6r9lEJYd
h4AvPnPfWu+InmZ4dheVyy8o91w6NcthtVg9uGiXsWsUz3FHHxncUeFf6NcEap7H
KjwUiJV8b/DXjDuas2Ei+EmSgAbOFIozmHQyVQ8gsNMllwXP0+mO5QerO53oRhX7
6nO1BsCBDRc6ZEUcECoD/o6+5WR3BJXV27H+gnEe/lyK3QerFaPtF12KrKt7HPs7
vwJYGBg0V6Wua18k0FFbKAQfEtNqqTx8Q6P+m/Fq51CyJ2eysAW7P9hyVLLNbIhU
EIvW7Qa6FJLwgRxuaORje3VelvTpMDCEmz/a/1zgWvnVHsXXhHzn18Ugfd0VMhwC
c3H9/TeS3gHbNrz5MTppx9O9Ai7aLczE6zu5QJp07tiajL42A7OgDiGy+j6YDxx5
I9obSgGdHwypp2Lzzyt+EJZteG6FBllfWJ2hIOgrtbRy/YKPmLEJmRPZ4AVLpH1e
xij2N+2Iv/Macz8w5DM450aKBbojqitnVt3XENpoLU4LTV6rdhmA/NJ1xPw+sDmL
OsLS6Yki6s/SpKZ0gb+wu1Vnu1p5ZKALKmwCWALK5DS0+oZFUYDpINuFych+OPHI
Y4J7ByFS6ITbcI4AW/B9i6wgvdYO1na00ljzWB8cg/m9MAhjO6ZLg14WNmvpfen0
fJIeTNk8IZK1EHY9bODeJ+RlBzT5wrFM9SAWIB1v8cxREGbdEkECAV8RQaYreC4Z
Mjg7JEYhiKyU2We0GqoYWhy6ngOcj0S28sx8z7UagH6k89/l9SKwa50/G3h4g4TE
rNPds+fYZ9jn8fd9Hd4O/JRA37NGKQ5UGrZveNiKBkMtwzr5th3ZSwQRT1E51eID
HPyoIydM6ME8/AA5m0js2Y40zasu7gq47sUsMqwxhzHiFNZyqvIfFAx+9aBdBiB2
/iINBCTB1hqgbN+BBvU1Pe6BuzC78uxSHEa4QVSfS8Tsr/yhUBf2axFOY3B2eryN
97TzJdQbbe6zvK/rfK8dN59NX1VTlhclgDUOCUaoOe83dpqEvL7ZoWMMdQ/B3qdY
VFNG3GVSZsg0xzyRxYto69/udKtDm4pwWXz51P5zHPKkBEZ+vrghc9GSCW+/k0Vn
fkma7ozQBt2O7FOAbeQG+DCl4uq82wOylbfP5SE/MYW7n0phAZq8DOBAWlcFRTZW
BhqxtbwXwUjL0x/2jGkAFVKJUG03R54rNKVE0MmKrhCeV91B4Bkc6Ud6539h3H0x
HXS3pm/6GijRF2r+yITFIHvrNpXwp5pULesJ069SVyb1mAH4TDENhK1PT08SpMYd
ud69hL7hFKBeYUIUqn3cl1STc2YdSVvJemYGKbVnrJVi1M+fXwkr5IUzbHe7BQh1
GXyueErIyrLstnw3U22jSE2W/ESc4jkN0r9mH7dsTnD7yUivtL/xWxVF0Fbpo2og
bOo2NJO60e3opHBiWRytdInGjrUfdt3ifZDmak+GAfFSEmd4HISUaNa3LtW5Tz+3
S603WmohZhL57hN+bcZIgUbhDbqhN6fO1JvKyghCsE5SwN0TRLvOvgTuiP1pikxr
Cdpx+JMXCrrJJ8gWFKWiHpr/TV8aMMu4eCpJJivB1tPMtEooESPnGAeB4zJWmBWG
qjknl0MQ2KtUwpQsS1IM86hDIaljlJTNBNgaXeoUiV7EiLTrS4wTWdpoLZ35Btz9
Ck89BAqE3i7JqIIY0ioLFdrmLlZfEl0t8pf+0JgEB1OFsd1J62IvarVJIzK7ORB7
He1C+koJ1rRvZUp0Lpk5MVFtAVQ/4olYFW5HnyaiP9mRZFhtpgcLu+GzifYLGU9o
u6AaKjGG0VscKAFF4f3+Z0w4Eynyg+U+/Zr7Z3ydBWCuYJm1EKNSFnMawDbRgxjr
vZCm6qRl/Kd7GeXop/XIlBIF+eKTMk1ZqRuXB4RPiijpGaH0Pj79iz9qBEMnrO5+
4WwXjhLIVxriJ3IfhU0zO6ew5lyxtdeRcfVIkELPBise2dZ0MNqo/yuG+zdyw96S
HI7uhZRzuR3EhU8oZ9f0Peei4KzNTZ9HxkQuJx5abTovKYFdD641WPrelvkWv9bU
JWFyx2TTjwlvM/11cZG3yQP/1YYXsP/DAgLOcQvy4pUX2fAIB0JFQu0Xi7s27j9v
ZtYUlyNY+Sx70cvb7aqgpNckSIgmpTEOr11LHzyCkImw0yu/xN5DZyd11kvKJcSH
n/bWeXJdx1bJNXl5p4WZWnfN2g4VxoTDPQenOgIqqedNpNy/Qw7MZ/DeoY1e2ru5
K0juYuWt2BGtgf4oBPI6OweceO+hQDk6NSvHH/suFkhIbOI80aCwBg9tO1SdO8nl
o3V7DDeuuKJbZn+9H/d5iJvvZuSCOL1ewhs0C3SX6u7VguFn3cTlkxFfc2aJmVSA
QKeFvkMs9NEvnqHx2XaAGY63jtE1syv7V7ohulML677hlj1pOIvtz4lLQcjT1dBU
TCH3XjpTfT28HuC8ClkfJDCP0l2Xvuw7KMUKcOny4GIXHpfWu5cg/Yl2mlcniy7s
rRS9lm4Gew7cyIPfuDaMwE0dkT8+eAxdV6NaWJ7Sgt9hm+HsI3kxRYf5r2IuyvbC
TyGDpPrMMJu7RB+k15miTI71aDK0u67WFGLA954ErPiSqpXE9L2nZO/cIMzR5EG9
3TfOYjndsVbtZQPRusGBiqKuOV5zPiqfDggu0ae5XB+WtW5Hj+nZywh7WAGU5Fks
vl7RQsTqLJefBg0dQrkuxMyGuAQih+HvnKr3bg+wwwa8o4MW1YvUpcgg7jxAJOt1
SWLbpQGzEi8yNMe0zOIXu5jDnj1TGuDKsRrZWpv+fVr2FvZKRVlGwZFyeLZ5n0qu
tjtiZ1jgxdTjJQgW5I1pXgTHSn3JGbaRqXMGqFYd7LzeSedlV3H+cWcYYAmZoFYw
cnKp0hIVA5MwvV/gxIOe4AtYvapiSAL6jGb42z0nUwwCnyBKIuyTiwsBCbaHNyEA
9ouemmiB5rWUqS6Sb+jkBs3gr26zsuHcUfUtrcb/NjIgFcid8b5symRtZFmkUFFR
3VJOnbu7BA9z3CP80JIzNVh25e7rihji1fLWmNeeCawh0J7+u9YToH9ag8spBV/n
yOFzVMnqvUSBdC7gGEUp3Y/UlF0rwMIYHX6rChfzh6kxveDR73jkfuDKMrzkB48q
n67kTy4aaeebqnkjtctlhwJAaxChEDbPOntXqMzM+lWJ+FIflIBG0ElJSOztTevR
3GR1NdDm2WaCtz4ifyjUzfo5ly4YXe2CuJ32HZ/4y39Xu0hCzhCrrZlac7awNJ2S
crIAo3k77/ZAGl1BaAjUHbfV713FGXgLrXDtEPQg3w/48L1l9q/22yNv4jfqe7bH
7+lT51tPiLsM7/o7Qk2wwMLeQ4T0OZx8liu3RBJZ7w+1vhuUbS21y+hWyjONNboA
2o5xwCRZuCxsPOLSmh0bBW3qoRqT7skOeO5F86jzZ0RjDnsoE+ILy3z8kSLVj/++
GdLPwmQpwQVmwqbjysBAP+yDCxHP7g1S1xZ3aV00z6Xv+HW6ceR/Uht0Em1BoPAC
lCWdaOafONo0kskSQVnwaCS9eKsf6VVaddyVmhxAZgr0e5N77SapuzxpphRQtQj7
uG7ckiBJtlyGiuCLn6pi+nLbdtDNKmzd9zgTCv05PCyj0Y7FMv7pK8EkzQ3k2EFQ
ToJ/JcAQM5+AkZJs3VnTk4ztVV5f2TdjcbHFyPMksrY0kg+dHMKagjDgoEaLoNGf
I1np6kxnlusFtFjZtH0LUkF4kvieyK1kI/ByzkiJEjwwQm7yHvDek89BgBUaXdOX
PvsXkNzjyPljVQwzKg7p01bj2TSZS+W70+FOHHmFS7L+jOlzXvfGuwXRxOASI1t3
wGAdg3Kt7Ks5sx//sG6NP9ChNvEpPV0JC1QWXuM9lXI/IAUbeDv5jQmRHJTw3F9B
KzO3FU3+X82Py3CUZnRgoyzrpy0Im3aFR52Rec9gX8TJXH81tumlQAikSV47j07T
b982lNyWU/62M6tbMIN1kS2DXGlLgmf6Ev5nBhoMfHtL6OHK3JhAZXWyPEi8Tsf4
R4SXR5x4FdruzQaAaM/SykisZpBpYrSCAZKflXHrwiJWVxZOqTf9saz41JN4Cx5J
7yASTOaNzIkHjyRNkOLwportuBwmx9U4gddsbt5aRWpQtP3TqDCZhDzTB61F+pB7
k/AmdKByhxJPPz7dMQQ+KkR3uxgUONCk7fkw5fC2moNj5ByWaP2agMAhe5qbwYcX
N2czrrzHcOqMPADe6aRFAz5EWsHLk2Mx+ExzEPbSm6PJhnIvk5jVZGZ+2EKR59I8
6xi3gQ5YLpMY8naiHoQJB4Xj+aLucZ7XBwEg3DGxaJezWR/nvxRDMRiKCkDkxFCG
qyU7c1Y+Fkq/JSKBKMStVDQZHuoXdnDIFK4N9ug6h5RNinMY7lnm0AzLlq6wN1xe
UIrKB1HrLHf0BiHUge3ZmD053hRlvkh632qHlv+X/9U3tM0w7lo84E12vf1QEbeB
83cOExJvC+HKZsBN/tS+ITlSDXdx1VaeWDK5NvpHaxk+ysOYTEqj7EJAa0uKfQxJ
nLrU1L54HRiiE16lQ9IqYEy8XOJbDOuJdswaDqGFsLRIA/y3BIq9graEA8frlW2x
4RgLfLtBIJEZF1lDcl2K4FnRPiGAmqsxI4J3toALCei7+DQtEYtVLMXY2lOhL0Mw
bEZyL1n8Ss69qxjF25L1ujXY+D3pMHpYkf0N8/+eyIut9AaQktI7dSWJ7vgA2ATS
qbIBK+/076gwFH5i8W/JgW0Xlr7eUS2YbieThsQhTAW2a7MSgGVd4WGBAbIoa/1W
3Hd+sp88SHvIBwLUDuE+AaKbEybzWF5JiWnf3ULwurv2DoXw22eAuWfeJOUOqsGw
pdgKbFqHHSHxU7IXwda6Zg32uYi/tZ7Js4mEekv5Ugc95ok6a6MuHafBDvQxtyl7
IAZgkXoPisqxBy0luE2lW8Rl3ZIYyn0SIyu78KL9FNGjCZNtWjfPJRgd2ugKqo9Y
a2o0lpXBK/koDnjghH86LPNbzDa7cYZfM/dEU+o3JVQpQkpuVhpQF0LIJhArij+x
VRea9xFqDOp/Gi+cfgwR8PbG+pmItIApVr2MB+DI1rX6RmQyJko3V6Rr6d46FCXm
yDyfICdqSzy21LfWaVwaGBPgis4FnGrf7nfVOonPJVfdDDnXNO9M+eokTdjpfRug
fha72gH5UVD189gT4zsfhDjzkBufjKiS530/5toZpU5dfcloKgMa37MdUwxRjIkQ
r/g5SlXYmsKNDY4hbsf4rREnqPNPqJn/B1YbzmAZL2y7GfdgQB4Sf8heG4+eOi2t
+UnT/gLnrvdOcvVLAktNwbOEag5AAJ3h6j1DhRNxbnEUZ2SV25/jRgTfDD6NclLH
X5oqKn82WjViwAshW/Mn3S75O5ztwWvN2UrzKWx2kgTrd/r932OPtwJtJZDcbd0t
JJSQOPDUyaRg6M3aOU1iPe3doUf98Sb80MX0iAU2uVVmO3oMH2aJbRr2x1vf7/77
DmoM721bOBdBp+W/CB2flgBE65yAROeGH7XvlO9bRmhEQq7oC+q1zoPsq7jQTwPq
YUc6ZP3t4iHaBHn3ahGihwYucxc4/YbhB5PWo0XGizrEzf9DV4xZLYpPUwKFYsgd
nwFbwz/MyQ7fG7hkK7kq9mVSuxRHmDO2MVH47ZxrMZbVxfy45iFNCCbZgDoC5tsi
w5N00fDwgrvGGfqTho9xn+IX1iAGJ3N90zlnEvrkcjIF+7JXwzEINP1poSnAq/AB
r8/RYL0MXgMo/JWM73b04c2+IlE6ry0ff6vC2/xWF6S8nwXETuyXOiLCWkYqUvdT
i02BYZRbKmor3se4+y5XBzFXL3awUt1bZ1k5E3tqQBmr3kB12ogbcq5I6vzAarBz
qc1H6vK2PgRT3Qzo77AiWeGLUxL5bQtiTUdS2jnnKcDAWdDT1XHx9NnHvQvupWrN
iyMR/WhZd6FJBqwNj9OlQwGhMStKB5c1RBv0TyDDLdQYOKf7no95dWLqOeffD6Bw
z+Si6QEtmJf4LdT9PBWAwJJoGVWYWT33yyk9qYdoUG64iXRnxU4KGmQQbImTbH26
NjHH8GUd2NaQgI5bWggxU86dcyZ3UVAerj6dlHQYQHg20Nf2VHwR+JMuBH5wcBdp
DzamewNWvVbvsFpuiqdj51LoLns61BwZ/3crN2M2gpkyNfsq7ngCzBTdHN8R9A/k
ra874WkkesW7bXzBOP9g6LClbkS6CSxrK/wo1PZV/wiDfnaeMC4dNJvP3Z6w02RD
CMj2xsyRmTdPpEe6/ubtTskjExLCR3cmphhg1QEstQOm7ZAG4wGNEz3SfqEQOO/o
xHSm18Mnnp5vEUXJ/RQBhosd9Dfvd1trwkKiOJztWO965SktAWumVrmYw0H+fGkn
OVFI3w2JYL07Cl6airF8AZBhJdgVkn3rX1pdJdCyDWI54qXodnJHKbI+bTujDFPm
wuQPokl528RGEGvjCNyMHonWvkGs4tMYTehYVPIX0hUKqRTeiMza70rPXecIM/6R
GLUfMlldp+rod/08u5uh2LA7RglHx+vNZ9zxwWi3tVU054bsLJ5fjpUFM4DrcrsR
ivcTHL1A+bySqbzlhimIQJU6LrG2XPSc+QUM5q/xPDhqmjiQT5sBab/GwR5MXLzX
/P2aq7MxbTaBU9o3ID90vZNu4PRywkKiUgLUstYzvjhBiQN30Zl8WzZJ2fADB1z7
ymfhWHEpODCQcd9ewyDdLeNbcJ7A3KLmqwDoJ40RgsWbY5cpQp5nTArD5I7eEaSX
bB9AygEUPh4eILEeE0iEcubFO2uCQZbOzIyis4YUmWKelld8ClCezlRu7AVpcGkP
BkmQqI5qCp4FrMkuhezTdcDh/K6NobojfYU94bMTSXATEv2dHS8gXYXqNguMuzYu
tocqLuQh61smN73jT/m8f8yIofcxDJKeQ+LOyqp3+Gr/c8OKvK6SnJa8mxs36QVU
J0pG8lJerXCR54frN/DBOH3tjnuR8vg+7ATQ0n1DgfVBMuheXKDJEjpUbOeq+zz1
mpolbwcNmoDSjNnat9cdCVHdWwRsbO7w9ZQtB37X/+hkk+yCwlSWUaaaUGvxPF/w
kOXE6eKMhc2TE1L+88qvJT8zEtr2xFRxOkMJtJgM45VXhj8jAjEAz9OkAO+/o3PO
cr8YzbaStYTdOcsO5iOCTn48/d+evq7o98SUxhHeYIl7Ws0mXBOnVMJcnRm1fKzG
7YAmLeRz7rVY7x7twcyVbzEksG+JdmeOV0VSQxj9pFH1Oq6Tqixhw+R4zbx6b6Od
G32+7tN5Qa6k7sezNKnuj6dNCryTLwMWaIELRpWzRiqGgBaj0EgftPWktgCYdTSU
uRVXrYiCzCCiAUn/q/aRWWp+6N8r+THklMxly52NIbBiL/rbgr0A6hCnjHm5oh5K
pZLExMHqMYEZt8v2nti6kZDRI3RgnpHqBPtkSJmIHM7SlfIKgXCoCZP8krvsixKG
lcEOQSwceSlJkqe04RV6mNvus/f7EZih/etb/7reMxTo/qn3RYQ4lzOGSwfF/c+I
YaITQIyndaB4ttGOqJUH3KdhqHWbe81sbYJYsfuCIB3VwewAtxuOprbz0z90B/B+
gP7LSkA4BAZxzZ9lsszxl2jfp2nrb038n2TTWjxhj1Z+1TdKlFYDFmOxRJmaGJhW
twt8aUfExuA16WkTUYdyvduxfaO1cJie5TvfAOQfqO1EOCVtIEhl0Z0IzVFTrq3Y
L1bSTlr+P7nEyoQyDY+Hif8iP0R/RaEWaoPUn8zz/vsjR3F/zQS0M9U6/EEX+1Mo
gtmtyeYXibRPT5+zNJgIYSytMixxubHCyf8yjRK8/bQHrRjp3CVeV5bnMXVO4vIk
1RjqlQctIn9gMFUpBzv2+7Iy7O9VeOxW0tGccdXKmMxwsAi1e1sOnpP33kDgsFzM
Ar3CirkTGe1x9DD/kuyW2SNtNdlLVGhCGngUufdi2JFxica1pwI4c/7litXIMcz8
g0bqDfcC8J3s5sV7hr5/3zqJdVoQYa4r+NBB1mszZgIEw0Y50VqhKry655lyImej
6qeUV165PoXN0LTms3qa7rcQ31tHQuGt/PKStbRg/Vw9WJ1Jx3LstxiZT2gt4v5n
aDxAtapIKjHuZXok2xXC+6B6CxJ7VpW0pGtyyntaSCc5QDDTyjPbUr8I6itWfWs4
w3uldzXG7QkVOnqDqAIPujM6m/iTklnSMBXhQnlghDTY3soEz6sNEmGJSV5SlLbT
p3pJL8SwOglqUBFzX7BQjfCaBkFGDYNaKybTszaeTOZdlCoF8C5cES4WI1c+qHet
B0OYcdD0T/yrF0FDtGyGqvAnbDLi093gSq7LwYAPq6MMm96mYkOjn2wOovG2GQmz
FGw45Zt51oBUhKmREZ+gbTMiTfqa0XOzmlONvGtbSqlsOKm803NQPb3fyPDS5Q0O
9r0xVLPaNGjslITDbPCuiVbmI9+q4xbgiNCJGwwasVTfz6RmvXXNXVeKqyG3wjIQ
jpKBqCctBhxDxsJgsS6VI3arR2O7AfcmYvSCMT3h8fv9sBrUg4S5dkmuTyI1pYUw
g1J9FxkrbugePP77sdSCOgRpUDM2ZIK6cUYNKVZVbrQ7ZBoKEWFH1EqFV7C3cRwa
yqsCh2SekpX1B2QJRdUChSVmYyWPwbFTgzj1XC4vJraAwDC4gfwdm5lL5+8fVFIC
cd5H9SjNm2vllt49uevafvAoNJsNWhS5uROD1+vn8dLeSMCYPEevfefAATUrQsGH
cGXgHIi+iIC7yyvn3OYJDEFBclw1H1iFkj2DKnda0gZBtXSzYe4H62RgBdtDHNLw
32FE40EEQAdPQV5JkhxzB5x1nLGv8snH/77eeAe1vRBTacX1XIa1y8mF989a20Lm
BxmmHUKujT20mM5UARXpghuj6U5a6jYrmGZcCgoqg7WSrYZO3Jlb0qPphgZg16cM
nnJzSdb6Ub8pGxlxbY59MvA1g358wDjK985wZ3Rp53iswTBzIVntS4XRIPzA+HRA
hdKjNTDjuSynGzLajh1N4nmhkvHAerj4vleLvi2ytEhAJP9vMFv8hk85IAaNvg69
Rk0pt+7UfDrtpu/fvh54zgOp4Kx9yliSj3g/xhVXF38QlcpZqnZAh+LZb4xjqWA8
f2eSUeggPSylC9wmvcJhJs2cynffWMEzB3l1hDBgqZMwSAg1AR9VBvI1I39tq9b8
iGYL09ve3T8QxJaK6Algjmqwr2996ODUjrJ89hwBXFNXpZdBAHiOWuzGAO1NHnsm
aVm+I5TtojIQCq3188GTIrBjlRBltX5LrPR+6dHZSWmERlfw87AW8pTkAxV8LzXr
+sK4JSpCLJ4QOONYxxIZDiJQfZ0HlpVOjaKnTL2WYw3BuYDOltpMcgMSDAlTmX0e
nWus+66PcrE/feWTNOvOOEHaZoFg+7GkxP+3ergo4rZX9BAybUhhOGdeGzZ/JcAJ
S6Nckx1CKlRK16KKvRwKcw0defy2VxpZ2XmUtzYxdWjQ3wm4NMF+EKddwuM7REhU
5nMk4mgMbT8+2H3/3Wz5DeCEwPrO7Tr3+nF5rEkTfyxx8DzqSp1fB7OCQnQz4RJp
LKgXrI9vbuIgjV1fBHUExbFPacEVMkgLZ0f88Gchx3/x0/86DPnfN722GEaJgqyC
yrTeH/wbwf63GHhPS8EOtMXm6Ij8LFV37OZQG1tIj1voWcL3ztZceOhLFVDtOf6f
OpUFhG53fPMtCYnZUyB9f1wCrbv95HhqjeJkljpyA3KTBCxOX4NuSgLaaqZ5lIkT
CSEs2R7buf3TNG6Dl+M78Nw7lwrwuSrToiltYa5CUfG9xWWbzRnUlV6l1F8SbH3V
FHmqiFt0OPbDkhPKcBs+kmEQT2F2jIubBamQ0WNa2cdmBfvQZmSoI3A+aKyYx4yB
32Ml6XQqzlvPY7Tzz1YB7cdClFKC5tgkRfmbsES1H5bXEEDOAcId3a9OhT4PRPuY
UOCyjhM0m0GfrqLOhq7e4bVNdmCvG9XMcgqMuZ41oGg0TgjbwbZN/VFBKGN51g2X
SguLTEuiyjjE4a2qfewRRuNW6iVX8XkHcmgPy+opIB2XkHx40s1fbz8TFs0xccgu
ezx4VL+a7gtyz6TzVpqqE7KVDCSL+SfFam2u2SGPt4wNT+FIFz6o7f4IMdl7JI1U
S0pvN7SV9GnYftpZIG3eYJk/qU/+YfvPLrALBMtjaC8nfAAUAAml3sWrgBXY5rc1
bXmVBZqy0GfWJf+3mXx6WUCutY7VPOwXno2TD3zMhUZp3fbG4OUwQ5lF5I7IXkoO
7O3jFL8EbaIE9+6ORT6QFkzYCSANLJhhHtHA7GlGClHK1qiesmXH3GYVasmOI/SB
etUiFRrgDSwg4ioCn9S3heKfCiedqcVQ0BMj6jmEXocp3HiT8t4NeVH7NljXBQrs
3Ct1pWNlnUoSWaOpFcya9tbUlmhk0n5M70DGLr5qr573aoquFsUTRMa8TxJvNej2
6Au0x6ynC7SffjjMy3FjSx6nRtS3/TM2/qm+bYmsT58AQl7cbZT8I+rbTTrQKOBM
13PIk2UKyEgaevsynN6WZNuGMIkeYF6zd5nSuv3DURIA7bYOYoxx7+xfc9tJpgwc
svMKyYdg/uGFiy9YCvM5ACacVZrnnFgR7VDqP4YotWsfpT5oWXrverK8u7x0OUL2
yc8/AnuisWPJ+0OzuUKyNoEAKQsI6Y1/APxb+Hqqo/DQ0vVfuGPd1MxsOCRU7Fu+
J2emduH8Ld7pBeJ+VqBPSLC4tOfDCsdjSh3hEVUf9SAre3xgNSt4UdACU/qOBapr
XaUsoxjch5LhCS2oIcpz/91Rn3dzHGqkylJ8/Bx6oqudaKeeoWJu30RE8EmqxC4V
Umq+1eK2f4erfU61w8ZTcTHEO0y7i9aeeNePKMOwDR6w3NZoeZ/fnhhRgEn8z2hQ
J+FUiNE6Q9zzxOAl76uAJdaOd0qD4/vym3yf8eVjnDZyIBRurK/OXVKfr0sFWqfv
CN/pMuOqDK2a7ovKA/FyF7dISuCDQ4FJmr12irzGdoW22XBUms63qKuE6LNi0yfn
IEIwohXdZuoUh6jZIhKQ6co01n6FRTSZMhEpd2CWXuKfZztvB1YOqYfV2BUzovig
3OdCDZN3dWeDgj45s8iC14wEDcg2AQTkiHgIB1dDCtMLC6pAKkZiO0YUncP3D7Zc
cDZH5jYZaxLsjA/4LZ9Dhdl2tB9FDgVFAvV+B1WqR/V3hHueXf5n0VGFHqQUYlPJ
dtEy5cMR7bGeERQZ/RlNu3zMFGbZBdBBATjSGrFtYR+5sI8WLzMRClzulCO1C/zf
K4STgVOBw6h5cue04de3LP5eQIdqNDyPIPMbfZVgt97rr+Dz16n+iqABL6LmNULu
jSy2fz3t5oDK95Hfg7AQDSAmdW/WlkglqiW760xtwn0yJtfif6bBlbh258f2icZ3
zX2KzLNLY3qjnvhGHzYfmLBRM5rKyfhFDtbEUPvEpNfRWkd+H1qb2P/B4U6UX+a8
+w4ps4+1rpA0RmgKKigEqizeLE8J57G2iiK34NiPsUA7q6v+PylPAWZBh7ocoy/+
lFV1OcumQYpknvB/3geArz5YzhsUa+enkSOy1DyeIrekVzJLkH+SGQYa9GwJi6Cy
+M+EcowwuveygLQaz9Ryj1GOWEzroGATmM9uTZJLSQe8eEMF1l6Um+An3vv2HjF8
DLKPGVwaQiJUHQuE3qn3znWDoaMokBQ1IEFWouUEVJTWS1KBGNewxTASXVz8lSFS
owjDIp+6Hwz/QKotxCCXTYclVzgHPG3LMmwg8G1GkYeg/MZm1SGlnjUYU2WAesTW
nW9eLWeKZEdhbOIuR8a+aR0doqgtXO5GGRCNnaDx+rGgvy47DOlfdun2tB58YHAT
jBgHAM4tSUvc6obvtJtSo916WVx3/9NbGMnlSJIO97YZFJDRJmLmOOa3qHke3TiA
XXmvixy9yQUR9BueJdNGhss718CiyGexQEzFKUZiIxEyhNt5BIMjkaq9dSgeHC3Z
bFm7wRcZjmGVz5zMaVU1Lvn3+SvmjlNKL2JnWJtkyHQY7BrvQ1gU8Mdiy7vJAB3i
/WJqUkA8a6ailEbzAdSrvjopX0bDW99ETF6ZERMXM2QMYpu7tcMGJ6aXmrNCJ+Bm
AXARrnzI1s+k8/MMe9vJ7RUWMuQocnO92OVqOsINPhIjGjMq5EyqK51QPylxgZuk
8bx8B+FIN7c/CVMKmYV9fswWsqKNAkglpqH57S0xXSWH8t2m4kNzuPPMI86XT2fc
A++43GcVXO/J5gCvyLzPPNkG2YYr7B7waM5D1gUeWlAz72i2z/z4SZ19Nfv2q/Lm
SSBaHCq7gMh8lpfYnKMa7MGfmYzoqb3GCtY1sGdJzaXsvT8Rta/6XPpV7DpKjZcV
fOSrpytTrRhLYB6hG46z4Ro8yKu3xdPKRg/t3yL9EDfy4jWqpUGIumJ1pGOLRuzu
Wx1rm7kLfgk3Xa7MhCKQisrizEG5QKTuxOgnK4H05AWzWfBDAz0dUc4rJ8Ufg6wW
s0uoMUfhIjdeYMB7pn9SkbhFa2uZlO2rMYZmWvt/XcpiqXQ+PkzLR7dIrGiv+GJF
TC6atREovzzI4l/MSW3SX3rx2V6ty1xNQkdO7KpbWgwctt/X1XpiJFamqIe95YDj
Q716EBeJOtUPKG0l2bJinnPhRfG5hT3GXMb8c34+YeyXw01Aaiq41N82bZSzfLsa
7xNS5uYmRLt9z98z8k6L1xvoavXgjcsAhFAm70m/9/xwa12nyP5EXQ+PnYosNxQU
FGkUS3xPZzmqjYukgFOFIFYLpPAyATwFD3pFcjHhBZTWEgDncDD9th5K/pVlWBLJ
sNn5aF5POkJ3D17ZdlUNHefJYKZWbwIJRwHj389vtrlPJeqiiN/uKqhtpp0tsRcS
sEajO5imSWrV7qj0KQIE5KkwJBVi8ajHOj5Nmu3boiHpaU1LDTePN44gQKOehfjH
LjNNrskDHt9dpeaEWTiBrkOs8LjlvA0YhlKlYd0E5TEfzSs8p87fDMGXAgIUiAaz
6on/RYoQPXQt4OIHHB/0NbPXTYvbN5TMDDh+ZkzfYB9IkF7RgmJEfVfWfj5chUgZ
RBXRWHsvUJ1Cra9YIOsYX3OVo5bK/GU6NFryIUG4jHniKI3pT0sTvOtju+p6RNcj
BJ7N7lFg5MsxnfvtjkTMLrausWdiCExcudGeUjxIcZiMHRU0VKHAHRw4WFlbVVxg
uEEsAIKy+4nKQBW2x1Ar5f4PEgoRfg67Kq5kC+szVZciaTpxwWTTQ3t4UzIoMEC/
DfJUSuii4RoWWwyGl/QjHe9Pn05SPy5Fl5uYdFXAgEvIBZbpfU30Rn0vL5sqVOef
XoXTQbEkcxxyWa3/6kNgc+hVJ+EChiWyhYv03Oo+W9CUlyloHuDXAnxvHDuZgcyZ
EG2q/DcVl3k64rnehJP7eLZJwcLZ5cIUZfoGgW/v84z1g91QRoNcqVNaXOoS9WpR
nU7Oek7R0CKqzeCFB3h3/MlLumr5GtRgPOLgIt1Hs726Z946gnd9mDXnuNO6GZNy
`protect END_PROTECTED

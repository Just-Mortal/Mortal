`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1g98B+APejqRku9or5Tf1tMbvHGyE16CNFI8ruGQKew+zkYnTI4HJd4IkNi1g8Q
/GaAkv9LRsoBTSIo8pfgbrYkvl6lvrBOT60OjrK0DBqzncXQxU72Z93l4Yqm8OHt
azXTQEIi0Bmw/DdjUof2TGZl8vik0H9l+/m/vKw/Q8kSfJ3ChZSR2Q9nesiKKvJT
lELkIQUOZwIi548B3xLnJoxmV5tMz2ISHu2nzuLTH49bncViqyWMvAfmDdVFho0Q
e0S4zqdnzEyiZPEfK4yjfJp9Cz588+/ut+zJM6pYlov6zkZFxfhGg3wdZkghIrkW
YwzNR/Qhm7UUY4xcVl6Naj0MgqrsMfQQGa4nPaOvH064JqGc4jDyRuhMUuXpKhvY
YjIBH6qYzCZrxFrIEggOBGSQBx4EBrTnC8YSTPaL2fYdCZO5T36N5hoz0jOh0hhM
0y5xIPaNbhb/OacqDIDUU2BU7iJZ1/+kwmTwWY6lZLShlmRJYXTzr9lz4tyK3H6B
eSyKwhWTwAyRyw0uJq4SOS6XTwBAuN9yIsUgiEGRqnDVI5rBB1vJH3ZqxsaGPyWO
J+S8bPn4dJta1dzq8ozl5yrfDQI7g3i9ZqYEr9klCJG7+HhKDAewPZlCEEnkjI34
BzERVyT0KGkgI45C4yjwQdiR40ax5siKzj43+Ud9Luu5ylBvGCUgo7TsTx/CcNG5
2pOOxe1DWbAmfg5OkrYvmkCJc77/CHZ1qiejWyyvyqhaWkRCruV73zXQo2cY9Ixg
rSMvy6dR1ZgSl+MTCDnN0BwAMQwwks0eoNXO2aQA6rV3QVYOrSV0Enqsf8qLg9gx
CFa3ypGB/X7bsOE1vdfTBAKjZUl+daDA6/KstivWBschWr5z/YTmux2hGbOK3BJI
NClIyjXbTNRwa5/9C9NgS1Z5SS4YxWVwtr13OIIPiNl4N8abhcLoH+c9bBo5pzfx
d3yKpuKQZGnCezmJK6+l+A7Cx8oor5lqcaSNu4aJipWztMb98ARY6ZWAzQlr9r+a
ljtLF1rii0GxyMyifDMVC6MPwG0iR0iAHbiG4cPKCwHpWRV7gUCETgB4sZfpqtgq
8168kfT5WPxGUSdD9bqkE5vDFUBe/EPh/QT0tj1OT6TyC87o9ArJo3ba4CeFB7At
5v7425CGngiuit3cpsti7vDL+KemKH6cEbrXcse7nDcHvPZ781kzMLPN2TwD4b6r
qGCAbwMcP5rbEHlWTrLGdfh80JbIevnBtp9mMlzijIqO77Bm5/rU2dBZ9tloT/fg
bMoudNL2zD3hrJ8KjkuItRbpS6jJq4vSbTpiMwgP2vdTqmCoZNs4u7e7Y7oMXWxV
vfW790aFKfjlaokWl5Mg0TiNqpMGBLkAhjoX7dMPYFIAE42PF7+V801j0DDLZ1Ua
jMrdT8J+WjMtS011XVp/YeV7FIdVfmzIod/aeJD7SD0uPCQ/VNntvICsDjf3P+/b
g7T+9b7vvt6ARKuKS8SkDoOFh3F2ale0+h3mMnNQDpnAJBfY5oqLXEfzzGFTshug
T4wQ9sKfeUF9dRefRp93TvCQyskzLzNbWR2H6F+z3FlDtqUVr9Dob+c/E362ZUlR
Rr545D5xvNpfnhGxjBrF9QExnDB5opml1CNgcPzGIGn3xa17QrMcno7YP2Bxeoxu
V1+3eQkChkhRQWlRu1GOw5Fg0fBEGV/Z0dg2o1efy0pfo9VEQXxNC04V6s00ZIT7
H5amoUOUtXYNIvq4Nar8v7y4c1HOEe8FSdYKnaitMWxoWhnYm6YHXRyttB5cXsiF
nj4Y+wfL9lS9bUMNKG8UgGLfz/oHE31wU2cxe/jD49y97Z7as0sVFvQTW5s+SDgX
q0ohnG9BB56sokI6GuCD4078VJ0WC4+SpBKvNUB2rDNh6VbzVugNtQW6fqu16JnL
40lXRn/OlJUOiZixl9ZVVRFH3IYjuDSmW5vlVTDUPd6ZJjfjj4kxPkWiz5Z+UOUE
76AGdI8GuGw0LeJ3KtS23UyOSBbwbspwFrn1MZB/HVoYaKFvUDSIPE0eC/nWbysa
3BmtbErj6KedIoVsztSKycK+Tw/lyKPJpVeN58OmfrM/1sxd/Czjbl3v68C7e9eY
3Xcy4/VFB9EyOp7M/UI16tthOXufur8idLTt/n1ydhJ8ikUlNUwub/31d+ZaDADr
NNZ+ArBtYbix1STnWTcxfFyWoItB/jWLJdssLR4sQuxVvOVF7VeCFHITzm7OP5ka
qv+nyQkrcIImPMvW1lRbTEO1FjXMDzi076jhOmvdN+k7VYXvjr6N78sBiqqVMypE
3Ji7NqiOAeDi4jEEOmHJ2hPY9mevryzaV09XC2XUvSP6DsKyR+JT2BWwBRltVtlh
E1sqh2BUKzMoMq23ukPBMtiPLFrygdHsa8gxPtH+xoa2HH9hqHZjmuHDxL9qUTR7
vsnNUf27y7XO/eQsEA6KQBqYjb/IuAjrqzdXEtXZLFN8x7WOhyZxPEuwFVhLHHu3
WKgnMyx4aRrXvXaE2hn9mR9qSs/+kI3OWGQVY6mSizY7Rrw5kQmWH/1TbdfMkbKh
gwk6dPCJy/JLE9uw8GfrhoWU8wjNh6BhICDR97rJ+lX2VPiaWJ4Ms0W992vrBdv4
AY2LSY5BcMycmclh0zAJSWNXQBX67GfUhWLlbwQXvEjj7BjAWoBJiHZfsKOLScxW
aJJy/uSI/O0VmZD0dNx5urN9uo3yF3l9mmYlyZg3nD3WyJE24Hf6vMv/A9pO6IE/
YJGCleR2r5fmA+/nZujyhM/UbFm5KAnVIoTMmVYk+3SCAsXrRIDa6hTkpzIbFzar
uhsQGVa4YG5evJ+NwdUsimOgLWFzzRk1VWvHvmBvoyQSkhNAqGb3Oyvhrg/H5SvU
KCwCLHvWyWsSmBsyMBc6rPUvgPYp4zPDwkSzNekcBevK9QeSFUoU+hWTv6XiOVoM
VLnJi9ap1OGWwVQpF98R+Wqk20lU5m9bf9OJEeMyGvQPnufe149TkBzCjPeCKd1e
9QopawH/csze3GKp3KZX+/6SZa0tqIUYv7ST3EzL2ZhvWLF5KPjdaKuUxeZy7Jqb
84SapxApuYPFQpyc5I2ohf4pFNPzFuLRjaZ5M/nZpP6YqVFHnvY9iH/6lbijFuTX
4wHIAS1aMGLIUrbioPF3i9p4vYDkAqvJk5cRjgVNYm6O4r57UXQi+zit28uIlUdA
FLVRySUqAgxdw4Y0SgQX3/GvW/mKlp6MkTMHUmGMmLRj01swi0IHbU5W34SEI6hI
MK8XhQiESc3uB5x71KRRyYcV1LBTc1f6ys65kIoEv5YKyZL03CBEebChKsUlrFEV
hNqiYz21/PBjWpfciRQyiPdqcg1JLpBOV0GnH67gIvaiHXPCc8iIBmvD6eRyosPE
LB3OjphsZj/sa1G09XiOemY9CrUCXmqwfG2P/0z+1hRD8srn0tS+43hxsojhwNc/
tj139u3Kxa6UpC7Yu4HYf/gSV7I59z490xJvJOjhevP0kdIT863UBvX5MvJoKLzv
gBBCB1h/S6n4Vap7OANMZPyuR8A2KUQVwZ587RCjZi/9gGjxayk6YfZsphZYSoED
98iESd8/U2aRNa0Gt5kfIHbrnaBvZgxKhYR1BQlItJfyauOyAG5uuvsm/QG6YTqD
QF2q6802TP/cak2Nhb/K8VRA+dLZdWmUmHcrRIc593szk4onHi5w7H/svNH/BUiD
Hyo8xrTEwuge5Kqlt+Euv7ldrTIPngkC2iRhcIuaLYjKY9DLI9/KvjMy6LvqAj3B
8zuAc8jyRe3UkfC1X5GlcmCiiwFoBF0o0GFXy0oVT9rTdYqW4ch6/zWv9oeaMQnL
urEOMNeDIiPf/99sQfuSCyLnmMdh6Jn9TsnabcO8qGrwukthxKVoVZGpQ+dJMkx8
NNT3p85Nv/+tfnenFH45jCQmP7PVeT5aadxpx2n75fGp2rw6Cna8KasZ97RK6wDU
Oebo6ebYiAHuHXbG2qeuLB5uJMrRJal7dpPldiT4PUuH2hH1yYEPNo81q+D5avbK
tZPSCeFvgZic6FVXQn3rG/2SS24y4R4z3DjlOkYFP+SDa51qHlcMvfqruTxKY2X1
y9kaqg/5t6jdHquiA0bXSO2vLfM/qRPGtZ6K39X5AIMgNyDfTs/Tb20C8i681FcN
MIt8peQF4is+hvmg1YCHu3WBeqPzGc11rtdm7ovzDyYzoLEsL8DGwds8F8CNrst6
68fO0Z0VCqwdH324zdgKmUBFFrga+W67cNWFIlwSxKInNPQ+ABgLzg38CFeUS+Qk
P6HnIK4Mvz4Yevy7DhhxmPumfH/RnwQKt2K5f2TX5Hq5/9xl/KyzKUoGIqR9vC/O
45Ulep15IfnfcHduHvwl1lZQW4G8jMxyVXkiwnsJkOe8busgDyd5VGfIi1dOBdL2
oYoWSj0PNmndCPt78vdrF1PbVjzEKAQG8CIj+htqnw9LbwmIt8h8ZTbrGx2Eleku
n2YAq0/flbf3ApI3ploCMLtu+6LaH1hAE9hdOLsy72+Jj6QneodOwPhWxqtYDvII
y7uJKjasotciEaSCT7MK3LfRt5bZGAxRiG8hZljP9WbQPZ9twA2JqDCwN+5R1XIl
71joPlRmouJWgiQQKzmeN31fvYsVt8rwiNRZ9hFJgHfxNGRdRFybTevteVrXpj7n
lLA/co7K5sAsNxqjcfaJ5w1x/W0kDhnV9cyPSaZhrjjgzpo98zjd3YoLpftfn3x+
ngzDncFzScW0ngoXmSoFoMOTTJDoFoobcN+/iCs57dqlLR+btyMAaeceo7WBAcvB
A8GOnWW/g+ZM3k5ClxqGmeXN7b9MODdPyAjtHIDdnq73ZI3rtNKpICuTBZ4B89df
0nURONTK9ZH+VAPjBhUrZSlKw3l9iCkUubCpzDYXD5mikGN9gzoEpLyB1kHChW1Y
4/sRCuU9ZqZArABGokJT8W4HCL+jvDib6eSRZRau/YXVOXPd4a8gkHUc63i1go0u
DoJcxUH2hg7LdicLx6ZUWD0Ik3h1lQNrZsg6YxBxXcsnzZlcVzk0AtX7pZFQL2jd
swpKqM2y49C5mwjONnfYVP6uLsOibVXBO/MnAqPTWpJrxvvPNaLq4d3fnSzn2Nhy
jIdI7pw+REIUzixCXYJRp79ySK8edGC7AGjq4ke/fpvGD3gUPU42yxo5S62P6eF0
tPRwTPCi/J5Fdq5/IC4NmQZVv91NvMlQxcMS2GNMfGbKnOYyAqKoyZMuLSN5aE3M
VVwFBgoXyPIoZAF4sKo2mIHd1GGJnbrTB7akM7EwHiuqsW34mu1jDxY4C7xTnOSq
96a1D+4dM0niwsCOquh+U/Q97BRKai6rroDNjV3N2rOrScIiPpqCJ0xB7f2X7v4d
drZW/vinmxKC3AtHtca0YcVwQbANFRJbMLM7Fub9WUKbHdwzgs0myEy9tgxcN2YY
coVAMKF8HggkSJExMTtt3+3n7JbKBqzOr7mZEqkJ1fVQMYr8nAs7ZDFo/avW64oi
50+D7ZV15IEV2D4xmk61FYbAnK4gQte5MmOZdcZbsW5HLwycmLWReBSM13Zyxmua
TCBLUPLu3IplT+1lPdnyLwUYq7iwRF+6/uzep2PowklG7bEW/bQfLpcCjUn1GAaO
/8rQo044DzMr/LXIDpSHlf12XHrEvKwGxF0H16XU8lriNSgZkBF5LqhXy3wDvmw8
cr1naGxFIzKYy621ueusBN/7f1GFEseLqE1t00n42YgENzHDR+PqnTiw9+WZlYKU
awCuf3icmgkYHNaA5zzWR2HOFNC4WCFyK1yVBaHSaIF4tpUFXz6gjOnJw6gB3rcg
qhPktEqCe6JSTQAFbClHiQi70EcBf887cArVhTjwQhdgBxVWNbDW43aJiu312RGb
SMDq9YjWbmG90OdjR2XCCwyANmzJs8AmN8aa4zsV5nA+zSWAturraHpeit3RDG8n
6WaAoQ99U8lafpAtPKyuHa8NLWM/MTaP+IypDlAr+0bogOdxbht2Wou0mfDqXPZ1
pPwxU7VqRmtc8MMgPEzyAoNWzJd7VG6j8AXMkFOuYXEyar1kCkPDlApAvg7oZK5R
HlaYo2BwpWOJWexQsJX2aNZVJZKoVhB7qYqf045X23HOfOY+4Uq31Ligj0dxL8sr
TOjOiZwbq15EUGqwkQcsBba0Y8UyNoni2dRaleSSZfvgOoQKEJmyR4U3H+7law0u
062ddtTrrjq+Ghsjb2+c6Pr8ti2GCD6tLh63Lt82IlwDUPfK3V3xVWzpdsf0OiND
qw9bT7mY1f9QhiYaEfW2gscmc8GpZl1t6Bl0kRp4pAWbBNF8XpjV7ffsofb2QKVa
yiqAVre8MtmVrFwC0PQyJHnW+lTOvIXPg0qA9zU/Y6o=
`protect END_PROTECTED

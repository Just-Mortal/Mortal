`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/bcwIKL//I34yfraKUcO1iYagoeAPMFbMS2TepA1R+Z6Z5MH6Zc2c9HjN6l4HR5
5qJoxjUfk22qoxS4rLFyj/uSvkol/t3UKtf3gGlZLe/nOUdtJeSD762Sd1y31PUh
Pu0FAWwSXm8ReZbNzOX2F1Tds38R+03YltLO21KQTSGmfMSS2xJURqposIHe9ny+
cS1qTeyv7dDwqQG2UvvXqse8Z54jK9uCx/t6eenRgXHQQtLCdoA/kIHIY3dgpel+
01aekHGUzLAYHU7eeOXY+WDu/f3m1U7OOvlAZaF221qYvm3IunXUfI/SQKvVseAl
oeRnUsDAmA9djcMgwL95MVLSrO66mXJOcHRA+q7OKjgmOCI8LGSVzu//F70mMWoV
FhPqGKKcYoEGFJ8Bpp+jOr/OmLI6h08CYy9Xu7lhLsMS565xEpiBOMTvvt4reOFV
QzYwZTK4veQrOezcw+MQg9v6v5Ufxr9ETmwifw/WJ5PjY6Jv0pIGsw2YZDBL1S6P
YUTklQO++oofFH3uiAynAWE6p1kg67mH40Rzo5yG1OtNRyYBtIfxLOmYSGxH34kU
/N7iq/OBjuaVQ4bjHBI39V1bKmsBeZHXvUn6Z2XLzXdhbpWk8byzc+p6lFGuXori
Pvg5cURdYagDDxCJw1bg5pWsi2UPcKUFpR6u8Lrd1ZFjJ1F76XjK52YtbWNGJI0c
T3v7Eg+52m09+UoD9mzPdZC7vRR0mTH6hHJIBPTK7wtnNVq7FThxRGXa0piL0wXd
ToEqorrtiBc3jViQUQ2f2C1pFe4+jyLGP6HYbOYJXLn0RkZB3Egk87/dX3/0MbJw
jrPT80KVAXcFYcMoYRt03bkBi5SNV7O1E4tTrZD59wY31EGo/2+9jB0ZsxSoCycO
MJ//JNo4/P0DHtsfmXh4unpu/R47ctAouketnAxX2C2lOpotFZIzmwMdL+F//+y4
++qEFCw4iIkoIrAQvGGr7yq+TT+FABYAHKlH6nIHyn2VaL3RH5UM4ZBwNK1nP3bI
i0uYoHTiFGGU5WZBNXbAWp+ZB1UgsYN6/Oa1lG28rnwJLG6BOdbEpsUzuImCFtIL
2AOHLFTQyZCTtJi2NxSqN7OCbWNT3bAEmrTsbRDDGfn3teoRkO6rHwNCd8ux7/Jz
2/SfIRrxH2822s4UBMP9aRvg3qHc8dAmT4Ww9wQTZRWfbRncHzeCKjIaoFKa+Jf+
fYw+rtv1kEX6MpSOp0l+n4M1t/oXBmP7dpcVZCVFL/QMLeKGQ/R8xlodp1qpdw8g
9O5l0rIF9oCY20jdxVtSqKcyiF8pUvKlIe3/xiHEa92iVy+JfsUe2GV6Js6xda4m
tqeDul/DsLMnIyvbN2XVULrrFkWiOvJ6SXY14Eh9j4FBeMNXHuxkbqTzTaVcJ5mP
3el3UQQOcOfuauxlMmzK00OADQclmERiTz9B9TLqfoooumGsV9Rk018WOEYY7DCm
/VBDpSf4185lRaoL9WS8toS27Xky4JKbFrs99TkGpr0rCTnJWdpNylta98ACtMZc
D+AMOu3SSMHWOwqs1bD8y+FKLE+55skbcesp0DjNA0Ww8nDHPJwVYRro6txGD2XC
jf9LJo8Ba/+PhXgVB+4ClfY6LWO4WPcoE39FRbhaYB8fGsybFnbsPYvsvTyCjriO
4SADCOUNh4tNojpg1jI+n8/VoP8mtG06tIPIeMeBS6RtOX0p5YS7kf+kpDTGc5j/
f1zoLAFnTg4mElJnRksFaR83GGEvWhTENw6YBqwYgu19YdOTEiddwcFcDrfId2us
tgMgPh2zUi57LNwsQ5vMh72yC4GdWDtZVtss7WDkKFZP+vCFhWsT2qPdVuFrTXS8
5sAA5W9us9FCTAYrCnRRAVVKt8Vr9PmYE8ZT0yDj8luJDD6y+SWz6oaACSXVejtw
qJwiyhaGQzGw4nL+P8AMIr76HA9iZLFlcXnHy2K1AwsxcFuAFwgQ4RHHmTCbvJsP
jxT3fLPoxPhxcCMUWvPHTZ6cUn211/gOdCbDC18xZWzbfVRhiMkQBGERRB9HtTn8
bVkF0N1ojGeOsWnmnVJ4a3P+nQYZy7Ak5VbAFtZZTsDRQvDicHRmRmLvDpnTN75M
JhQ5/+aYqTBenPxVkxZa2uGUO3etTZBmI8nHA6USP7O9nSbyDDJmiNR3EazK6mCo
PtlD4BjZfbAUgTOEHeIY3ZFQ04+zHFAFsR2D8fC0b34cZkdVe+IuXJtgFVSlWb4a
IP9TM2H8iZTXE06jW5ACtuUd/TTCDycp8xmUVdTYu4ww9EcSaXVY6pYlpa74f0Bp
P+v9MhLjYaUZMYfZSj98S3oRl7dN4+RxR1NMIWxjxRDOZqECKsyZ7mguhYb9J8CM
bXeloZbvo8Rf7vgiXwlnDlxd+BR5r3Vve78D1zzdlOk9nLerUr4TyatKhN9rBaqu
zQI/KkxH8oSI1OHOBNgOJ2u3MvP4fvKcGFVPhWmUoZWhrnoP32brjf21qg/AfiNP
cY3G+Zei2iKiRUQE1mN+HCOLYMtAp4Sb+tHYfBHzHPQLY7p3YwXhD+qws1KGbexC
Up1nKdPCB7HQeU40e2ipn/CZf7Byd3hedxwhf9/FiMxxeF8KEjsJ62/qPESgQGJk
Zy0tRJv5Lfu2sRagvwDYQOQbrwo4SJzXuq99zB3c9HM8em7Qiu9MCSIvSxousWpd
Okm7s8VM8G6W/rDAnFlR8WTeCRzLuwefjybahsXHSWcecY4qTEtvLYWSZdO8SgiZ
M1CBePmtKYc004nDbLcXzvGWpuQki2Xk6Po5lEblQlZV1e1d+hByK3nwk0NiImyE
bh41zajJKMBV46hlvH1ZphezaPcIQO5tiPLVQkH5akFyMnkONOOB7YHR64/lQlOl
oKhgVP4tbmPpRp2/3s+hMdGGLEGg38AxzcDCyWY5hTFfsz4PT+kFfaPo0IN5gW3u
MyW1dtDeoRwwghs7BWI9AnhzdoIU6JaRsRTTlGnQ3Qm8hy/b7kTHIV40SuJFnhiD
Yv1WO5aQqq/q5dvk4mAl7LvWVWYeZjNk3iNWfoY+0n0i9J2UDjzX2i8XBcKWAle9
CUACHtvSHjolpbJqk3FroF8GIM7REeHLzyXitviJ1ZF+s4oL44mmTD65eshZyu+H
TXm10zKAHBG0rukUZE5ZmyTUYyOnuG72dSMeL3xI0gjXCNby3hmtHDuN8UIbaYZM
3nQL4IynZTP4g7P5LdDNtGln9pBjtDHEJc4WgXULyVVFcig00GSz0CSVUDr/BeO1
n+hEbG3mDJjtbjl0+udgCzSpdMLLOmrdd7Zou0glmoaec0+NGRPDvMtFMu0ks2xw
YQfGQuYB1Vft/2Zs108h3sxFRKq8Kkgf5X9Dj5JvwNNCS4O9xomq7jMbRaeVNfQz
pjn0P+l4BwwLa9chTQoQdtXuHYXI+s9q2fskPEZ5AZtlR/XncwM/Vl4RlTDs9+Hs
8j4LYgk72DASGbmV7xVzqEZWFLb4sRkBG3eTkkwQpeJpkiQ6SjzKsiPsQpU+Gmo2
uTYay+6KA+Talg7yAdMbevN0N3SQZSdAMijFvFHjv1OrEp9i9FZCFl/YIdL4r6xF
gOBpgbR8TQ9NHIceAO6APeryvK984Rn85CAFYWOoMC2k+eBGPo8Xf4sFU8UDoCok
6vAWbBfJyGg1Xe84PKnRY62QBwexXrbQyMjWo6p6ElZHPsKXY0F2FeEhlzFM/pl3
Ho+atZKVfQwmEP+ECi90JbsF8+kUL4B9G3mdcRZVtVDXbFsLO2NCuYvStHtQUlno
IzCzJzQ/GbuTIPcBNvCm6URE4qwNTE9Y1ZYDtE13h/k01Wv8pV920NAdY/OhU4+H
2pan0FfkfppRDatRLz0J2YSMCdM3sJVxeuu1c23G/9tZDytA6vWEN79vOFSDoncE
FdFAoGjJ0Z3qBQJtmMnhp+ZRj6kKu8rw6a95vrpacG19u8lRU9yFn4v2MgAj2OF6
h93xtirZul18nrr/wQJbt3T4Io8Y7sWZuuQQQ5rKQDAItwKSLKe2M/Ctux2zp3t/
7ySIgPS0hzNjW8eTISIsSy3mdscU9oRR9rUx+XUsetWou79oZ4NFvcjooJYZV0ad
27tI1gmxJj3zQfNPir8+QGHNy5Vsfw3lXeB28//qqzhbn2zNEqGI4by0zvlGvNKj
keYyHV/RH6FDmOi6fak+BcOpN0DIEmjFqZG1zf/6R4F4Hiiz5XIhRP2ETYLq5mQv
ZRwi4g/80oC//A4h7Iz4HrrdhjqD7p4JoR3UIA7TP/oKv59QgzkHRko3yLEWtw7W
M0FumHNimNXLrlRwI3DuJOo8ddYz7Kyr15wufmp0vXcd+tKlHk6ghbPZXd2BnN0Z
ZlVg6NujA5JaWAK+ZcYFPeGaAuicjTeDhYwygiE5KF6IiHEEMz3gfi5Y1CrgmkeT
fiQH0Lq0I2Vv/26W1vIzc2UzHDRnOb53F+agj7UmT+CVOK+Yoxq0VGiF2ID44y7t
MRMuYjdo5zy11pgP0Brg5oCpaTJbQFYBSeX0tqoCYVmW/PFJjapW+gUupS71lsEA
94RsGD3jNvFzTVonWCdBy1mcqzXywkVuBBdr72h9k7EW4Vf9A+kc5p3p81zJ6Uor
7Z1I1actQ8psOMHXrv0t6TXravQ/0EG8OOl3pxz1mg7A/6QOF+ncWN/hJ9dsK8BQ
BDFVt4v8ohIW/9Iis6MzJSMh0NCzgcUOarvO2sc6lNODBZefJLysmDrDO3XNhbVY
nAHExiL3oOsC6fmgXiuibIYfxFfiFTqeweHm/TBJJedNRtoRhljgh5aZPvsZ/VM5
7Tlwepqoyas5Fn8wbPC8IXAZ7XZ14nDV0PeInQGduGmZIKyOf/NNJoQ3nAtW8b7C
J/f7y9Q7E0t46FseaokG1JJzO6q03pSW22Nh1XgT2mNhnJHrUUGWq+opp2qFpIjj
DpZvzy38m0B9OjDP1dSSzi9dCCbfHPaqGnyZv339VCO1X3GP9EKhbAR4RNcsuoFJ
22EH8jJaOIOIHfGyU+KzejTn/9ptQjrxPu7oVi7Jlz3e5AAtaCbP61ONl3n2ZoQU
H6CRDvRXpabxz7pkJYwCpwB6M8fSi1B1/iBPTNTKHMkycYD4SVBn7qZe2uEF0v4p
O6BtATm0zyzU+ggN0WvGBV0DTmNzJVZ0ebyY8SEZGu0S2kRhOU+ay2TfT8FGJ/Ga
6YI04a7rdr3epCs2kSavM/r0JSe5ozBHb+o3a0Cqvnh4gEyCmFXMjFzezoSVjFGt
hOPJdMe7YUofo+HYo+k6K4Pw5lKR7omB04Zr23vv3dUhaZLWh6LtM319iE1B64xW
Nl+PgvCteAI5uDchA51JzFdHimNknpPeOPc2lM3qMl37KIsVgFWug0vFSlkD6B34
1N0vn1f/KK/mBM5YHqFMN1gYIthvqSWHsnuw9ypL45MltM+azjLBykszbf7/d9m9
YXifmGTNYLv54ozgZyg0uprQqu8E8MXNa/w8lZed/VQY2OAbeRvfKUZEPnuyU8ld
hPKoGPrcWJKnLy74aPVpniz2poMx6RsgGVssTxWulcQLkWME1sshHmYZ/daZtJP5
H4DGA8MXpbZm8EIETYvr/vUxuDikziWGaDrEulZVRgXRok/qvQL+bK13Ve2guGdi
LL7jlEm27OEql45XcmdpFpmYhUGZkxWtT71Rlfud4GI3RhfJXR3910ovofDtZIPx
hNkywzK71CXvKCu4x5oHZrEWn08WL2vv/9yYj0XW+8GkjRpxvBg0y16rspjNvNla
2F3JwbVed9F7fRfr2JCwr/ad0tJ1IKsoCAO2cYgIA/JdfTGVIiub9hjcwqJ1gEEE
nurvp/HzQ+VRiuIJEaGaud9K0cot/XIEu+MF6Ju0SIrXhEYqMPnbFo1WC+ZftoEz
gv0FKMgyzN/bWg+X3IZzOnbRIR32oppqyGd5xCxJnR5ZHmXCsfPkVXRj3jgquOPU
wJ1f0lCJN/gZFSRL/uaxNHkSWVMYp20QxdZ1tK31KWlSIpXwlR4CSDOtB4qv8IVz
Btw+X4mx/wSSffQ+MO1pgS4aZQyxymb4/SfD9ehB52c=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hU1NfyOjOEwyY+mRH2TUnSfgPpcNDzCgbSxXIPZ8WokD4O9SIEJV3fEuEqclRJ1O
E7q0Rms/FSftocZvMAdaCooR/xSDC/ve39HYmBar0uulaT/Q4dhUtHzMOD5D6a4H
ILVQDiHq4yGltMS+RubOqWdI6HR2zXLR3JqNP+yMMMDe3fgm47VFIBc5ttdaQEhw
6I7pxq8y6Mc9zScwv7E8vYTEg3bLpdOQexWDh+e+LH5E7SLaOMytgULiYBOaQW8X
k6mJMx5QgonPvlBGWSfvuwwDFwuU6LlIM70xMEV4MAkFnaDbbebBJcCiyDLJI8bi
kcs12e9kUcJN4L+rOzQbSmWLY449StP1ND4PeoL6oakkRx3d5h8xhYGnzNhA5wlm
Ao6ZEB6nP0bfOWVPHnpoadeA6JQKHaxq7EORa9dX0a0RWe9Uw/Dymh5L1yYDnS7i
bW/TTMnAafQ6+yqx2TA7Ctt1W4XqLIbsTfVI5cdl6QUEXfmXwBGnzpyNqB+AH4sO
JAkhdE9lH81ZqbRqUsWS0s+JejH3qBkkGzWyJmeliGzGVVOX89CtaQ1BwfyySuAa
0OisYaJbxtvgx8QFRlTIPLiO2z2vdF1+ukGP027qkoXuYdo0mjEk09XeMo09UH7/
mIOKUF5yg0g3OUw4Xtyl7CK56pLRgeXgvmt797tSu0FJeZDIRvRSvG9SMGR3vcYf
22j0/sVP01QnAevp6Krnu/FSjoshIPhUQSHl/+b3WKs1fQ6iSpSj1ZibaLFUxZu2
5riIt3PwJ2uv+NZN0zx49LwxOdvMShcT6oFsQvOuti8MljGmcamszc79T0A8q4E6
hyVCBR4XKwnFVczJ+kT9Q1EWtJPthCV7oT3F6r8LLNfcrN+b+vWTUBDYo2ihmzgQ
OocF4T3nJI0f+KDL7P9eckWfNeXxbLPGYxxysoXdEtQEJXS2g3OGUJGHzPJl1b0W
wMoDv4qaIDg5ViFFj9ra7QyBrmf9PGNz+EjmCmO9Okt0UuYXB9st3Cigl8TgAkqb
O0hiRN4rrm2GgAb3i3rdm3XYo+bVmIS/WapfOsG8OdcjtaIfKldElU+Z54FZ2/nc
PyVwVfPQg/1Tt68YX8eCvuZPhQB5DdAgWfmPgpECcaClqQSa9yUxB9nZbNRhPRC4
Ryq0dCm6VHeTB+zxbF5SYcPfO1A4SHhX544FHpmeuis2nU7lTZlwbiO8VXnAvQbW
aNxPv2+nRtRndPYxpMxBxkSCVbFWqcfTwz+hc+DVXecPDrDiGTObQ9XqDeWv4dV8
XNPrXhvRw5axXJxHJgRzAnfx+LsRNgUhO1AbhlnHO/+iRc8ShKvsxKOfai08TQbR
TqGzLZVgI+qZ3umFCbRXJ/MKwyxlSk2Sd7eFFnAzaZa6PzScGcEtNsUmoTRokJyE
jdCpdQKQ0Gu65O0NjS2QeXNFkEAeXhK0oVRGmHqKX9xsBalT+N1h11bWS6sqXLiA
iJtTOGJ8BHWmrRKxQUnGT7G/YCO703a7J89G3oUU+djopJZgCdOgsafpkf6Y+Zra
YBtsdfQplB/WI3po+A7dvQop7OlscPJHlxC5jKyR+UJMMAkuV8RtEe/ZWJXbYN9y
GqqZ169pKT3+TJB/LSf0Bu2wFK0kjnRVdGaMbxU4itwkAxn0g0kU8DO3DmXHcjMu
R+SqJEUzRBnY0UQKRYicN3fySeapHKTUCWMApqWYyDmMfzvNBSdgPhujYSrhWmVl
xOIdcX4jaGNz2zUCXYGV8GUp7w+QnxAHXjorGgmjcN2dGBnUFJ4KN2cIZ/VIl2uX
T56R+v6Me5ZOXgqw6+KOZE8XhGhdjEfSBTUH0sAClgm97thAnbZlzP8iYsrEWhAn
OlYTev0WVH4VFT3SXzdNlN5MR6Iwph+MedM+JfF3mBRf/e0hL4mKufHK1DlSFtwq
zt2YxHof+aEVAjrs4N0ncVY6j+j9SM5hLszbx3dXl0xsQRpsRifXHBvNYTNhV3fW
72hAHXctFSeUw5e+FdayGEwGAK7Lfnf44UPzeWSOBK7iEGhMpLXKZ3HTq/OkD52N
o7IPjEI/bpCHMQoPg+xrF3By7UcIghKVlDFqhaymTQ1cUIHL0CnE0iuyzgO1vuNf
958Zah+5GLjPiA/rGgNitiGGgQ32KjjiMFq2tsMQHkiXUZe+JVDPvmC0joUeg13G
8OOnP4MpEJLjqNLBrQFUaTjNgfwibSLn9uQTJTktRg7gTb+RmRHX4kn1x1A9TOWh
4/MlAzXJXWuCWT76wJiJMaWHXnnakUJ49wrel3n9YbBUJvvQC8SZFzED4nLRmfAq
8fddALLpHENf2MG5XAxACzXrev4KYQFmfSAjNFod0zyLC3AS6PVKuGlMflr2llET
Ine84kbrBKd6WARKak+fOeBHDUSytim7UWn0MKV3WBkiwyazJiwRuHOkOdUFxiT0
LCRJav5IoI4N6SI8pBey/E99relNxv5M4vIDgVIjPecjOTNoNb16Pwx+Kj2JnYdW
QvsRSOAvV45lbMxAUMIXOU7UZLM6OR6Bm5J+Xq8oW02dkbo7QcKu7z0m4SRsiGIp
YZPW73ULdNcVSqO22ugfaa6d/vNVqCm1l7/k75uKCWtuLSlVuObHFnG7daUFsaEU
1jmilN0+ifGboW0WdZbYwOOBIllvm6TbMmBFLC8wB0RAThJgqoyDiALUn/hrzlde
NkPmaLp+/P41Oa1F1anuVxdUVywNULK2LNm5Fsvkolt9JMOWEvV2ApSx2nNkAF4f
lQTyGr/BcvUpAvcVcVOL5FX1f5GHDayapbYaRm9egDIVIg8N1gohazxp0zxYNBkA
BabgRu5o06en6BxgyvstZilZWR/ZN9QeYRoN0ybi9MYC53twP44ljau4zE/LKROt
5AlXGqnNVFb4GoFaDdz4Z47NOwIbdfnP6CKnp06RZltF0ncvYMs+LkqNla7pJ2B6
JDppbEUFnsCBcXlTFb+muHF+TMCJMhQrdE61BrvazDeSotJLqfeAt3FgLiFVeJbV
+tOn2vhwgnFkAWuy34a8eD4l3XsHJRnbc8jWOu0pzwpdaoPd6AoArwl+TGlFNAxT
rXwTZt6r5YIeG33vhkq24Xf7UE/BTwtt0+RP4gLv4RlP6ZIC1cjid3/tFv6rwUuS
kHKnb+fV0rAfBW+JenMBUt67fbxp4d17YnYvpA3KcQfvDgUaOV0Qr9/3x2J08zLJ
jqxW475pWZ8OCSTdyr1CJrKBx8j6JeOfe7+/XVab22XsaM53sOZB5+2RibyEKvB/
HLJrzeu9yM6kyjy9ciXItHCOsikmX51lGGAFqyn3OCkr1gB+HDFV70HUQAc/OHfQ
uHhPWJPCaT+CP09vGV9wHMnLp8CdYFwsnzE2sebmhpEzNcKeanEV3jlT+o0Zb8Kj
1VVKWZQJAPLEN6Q1kkHWg2KmlMgVsdiCIaANKJrFrF0cDZJydyNHSzzM/jbk7LSM
FBabbk4pgMKmygXs33Foig==
`protect END_PROTECTED

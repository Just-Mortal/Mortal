`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
okq51ZMJw54q6J0/IvzjAyYjHQ9y7xmzvBpODk4A2vkHDz1D9CAyLC7xeeRQuLOX
x3V9zZ2pmfGmTjWbDeMxZ3WEr0VWlBrMYKirgk7fDWww5L3D2tE+JBYDNuS12uX9
XWuxlyNAqHKPj7/JYu1mc9bjqvRbBbv8cRhLa15hA/Uh5wrb6eRU3U1isVQy+dj7
nsqZFJnQvPDZtIcOKIk5Em/rNOKCShxjwmS4Pf/20m7xMVlc0nu9sibykx7waRfQ
wgF64z+if5nN4RfD35nFHIJz8TM7grD1omqcU7NiJ5rdIsAVEDbYBjk/mBWa3EQX
s1fjvJDsAeA82QXQWNte0DjuH6KbcZJ/TpwyRtC02O2YEEEloWG01+YtOe4+e2yc
07WzBqGn+LUsNSp7ucI2tgUuzAhg1TaNB+DWG6tWyL//YsYiLMkitIvP+z2FoVeu
amomKshzYQWAlx9kCHujaoTMy1mT5fycJITBzH/d/487HEZZfUoMX0VSv61dETa0
e0XYVmKmMfhGwXRxlT4ZjhOmvLRgLcjjT+Xds9pSTC1/KDbGO4bDeTvwuCOMEGFX
2+5aYUx2XnL59rllj0C00U0iswH92yw7v+pyZ5iV0YDQ95skP8irmKAM0vYCPzWF
90+GSu0F6SbkntTwrDfQ8SEi62H4fipaRnbDAzkjfytrQwPuyDMI537GC9IFgr7T
IdYrkQPENgfL4ztUdQOl+K9IILxz6fzIYVD0MIyBtDw0qoQTTCsSDa3XWEhV2rBw
ROlFH+ENr/dbX2PNVIT+L0evC61SAu/Nj3vdjMVrw2NjM8m6faVXFs6pjWamqlDW
K+fV0zVWJlkKTYyyksS9q9kr8BCF5wVjgqQ+ZaQgN9eHYwFntO9usfOPayEWUsz0
i4/iuLBja+WMQpTqB9GAwpIowvtk9sZNEvaJvZrIiwN1DY5z9aqGCJzW9qcijoZ4
5HWnn+XU52XXfsZWUwZQDcMLruGM3T+b2IpoXppuXylCE9pv0Cx8kjmIiqAvD6Vd
UT2RlfbFu/XKmbAC30cSDSUqQrlwY1qMUibdzUnwTWiqOBBPD5XeoDGls7dkv1/o
GFAA1g30VYd+DkcKJEXGUaborPNVd7YBZkurtLakHtXgwNo61fAG+/PWwWTXof7J
sBavw/PdCxiiB+iqupSjk0qIA0LqZtyDhtGPe/KmtDD+LHySyOb3k7JFRH1ornl2
4pbvVMHtaT4eOLflgow0D5UFUMDdX9mLgBlYLu3YIZkk5P/ICKr/wxdN4NpBRF2X
aVuYg/Rp47923Ug+brEvb085FJ5F1p7KkEV6fBYuQSuDjsbff5pIIYoqvGgF6ueG
f4Fl8RBt2eQxaYnh6igK0b5sWTHGAB7X5QUgNWTBUt3WkDwGx3Vx9N7m7V7uXezA
wpLyxxKMwXvbe5vw5noO70X3HNkPGUVX4bwr3i60bA0Dtj/on0lLGlCw8JmSsEP1
V7XZ1Ujjx9EtSa/sU/7rKwBm7nCFYuLbnAYzlUJ4fxPdrS/4go5qp7faZXUg1PHW
3jvIFS7Ei5EAYKwtc1k5hmOrvNLkRTUOHumc90QWwVejRKP433i/SAnM6CXu5SEk
r68r9fUa/SMSNhAtcUfGgKhQOuZBLolXad7/2l8tpbCjuRmE7wDWLlhycNDSlDzt
ir2V4flBlUJZa9nh+Z7w4k7+RSRaUZsxnoImj4hh6e+mu9zo6yBPFOYaXPtfugR0
4SnfiJb4aG2Ub0l+D7T3teFbIIkAvf0qnNtpx1JJKPT4JPWONfh/W0RHbvguu26w
sAiYZzItozfIXu9a20Hnu4u8pR+IdlDP964Gs3o6QrEqaBdPtrE9jYyYwkcs1Asj
ZUmia+4kaPJIok7YX5LwzP0bNF9eZfihfMQJdHb6L7bxK3GisdupuHIDhMw/HivC
lOIIwScrsGYYcqQFiYdIF0J6nE0+EGwz7NV1RFJVEJqDdhQhxAbN/sTGADyKqzJ3
qk1wvHvOTJlDmal6tZimWbYsu/XLGhrlLE5FZ0ug5ZmoGzdRemPtWYVUFCJPSsJ+
+LsnBMVWsEh1RVO6sCgqtQ==
`protect END_PROTECTED

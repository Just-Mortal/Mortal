`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xnhCV5X86BEpdf2x9BDjgUumqsZO3PDNgisXNxTBB7SX2sfprAQE2T7QmASoe2SX
bTnQuARk99vXBQ3/uXz70AdHEY+zVJeV/KUL2hOELhcuqoPwJkJholMG5ilLtVJm
wRi3vA+uAA6+fjHjHA3zQ87emwQPYY78OnIT1cg00Q1NzYER0rTamIu1zh0cADKH
+fNAh3XxjFbX0QQP70kx002iFLD5bwpV6QEgXA7Of/3E721O0Zy5JpywZS/3di9i
477atIsV5JfzHyZ2mrvSO2nsJFbli3mmPVv/OxUomoIEB1/eVNmIh/hMFNTrEJYD
9YOoH1NjNLngay9XMra0dlH4BmTbr78s0mpYp+1gk4YvscqsdMFIXUhLDZI/r9+D
coT7Db6tbkXY1EwuZ7Etjw25OMHlcq9++EoFJO1bwUJsnUJYu7Pg3E8caplCSSDX
GsVm3q3v4Eo1Vebw5fuNhsTVTL6Cp7PcKZDaJwUO5/DOXYUTrqgNahShdp8nL3Sy
nO7JC2Ay6clFB05K/1Yx23E9ZuHL5jT570Hxt2UfQhNBQKkI5LEOJgsLLzSD1+Q2
TQZGadwlPxbpCsv6vcPUPAxSpOn/sr9jL8qh3PUkOwLQaSvtd7+WOqMnFEWSI0n9
lc/FM6ZM31vjFv3aIy9lWlL1jrTLCDyYpyCxylpUEHUAOFkQbu0Hh3+sZ67O1lx3
xonQCUO2RhbC9SjyaG65ldgGOMgjn7Zmlalxl4fxw4pB9leLzHU5pIgxuXtrJGOJ
rA5Z0xDYZYe6zL3ENrQhxlzxepy84VQNUXN2VCjJtssphpsE1VcdmwpsGXkpJ6Io
S0Rxo56lFQ90N35vw1n63stRQrugMCJcqxZ6xEdIgYTrxL8ocvlgRXLmh+9PPcXo
po9JWJblHT+DMsydF93bcNC8wErXUsu7m18f5TRisIzVZt0N9U+FvI8zU6QDgkUj
dbzKCty9rGieT+rbbUhA68H/eL5oi4Si1Gzz9hvj1s4fKQGwZd+1sijzC+TxCn2J
fFGv496hulTR1d7X0yMMtzjYT4LXgLXIxC6qxYULhE+hnnQ3bdko3XXpDPlX56pp
apnJHv8FtNxANxD3phADGkSpE0JcNhc/FdpSUl/Pzdnp0AAdTOJEcGOo2rExOY6B
Z7JVjr6AO7ehA1dETQXeI62kppeJK71/fllB76U9eVXdu4viFuZdxT+3Fb2FDrJE
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UtBGB6nHNXbxCz4wqGx4f8pVRD3yHmh6W7q8X0FUBA5qrPASeHHHMUpn8AGmSuLt
SgeA3KnQSUAbsJoH9HPfoCpb8Co37X1VzK1aLY76J7DjgYdKyE0rrRn9vNAjUJOs
aO8oqdzZJJieZ+v653IMC2jpDsq5fBlF0vsFl4r/LiK5vSbp4/E5FTuYrvinqXSh
F5H/9+DFvNh1MtZKgu/YM/JAN6IXLqF6mkWbcQKrtVjonlqMQGtLJPtkkN3j80Td
H169KRPnmL1r8Rga23pxwrho2TRB82KdIJta2k4kbXYCNmmbWVnb1A/uRaD66IC/
N+mzhRqcJrODlwtg3bczbV8+W4EIzRAwB3E2+EtoBcQ=
`protect END_PROTECTED

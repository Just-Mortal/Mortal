`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdct9W4TnfCcZNCxGmnoRjfVzGNtL04G/Yi0ev20y4A1wugvUlNcSSscQh7zGt5q
8KkLrFHvB57DxJm2WRwP32XgCFCop0G/qEBWDdxI6RKz1krRP21/GbFh/Gg0I5iX
0Nd7AfoPZRHvDoyfGPH3Jheejatgh3AZtPuClsyNNsEQbY3tSOZeX7PgbhYsMFVx
ysdqeFHYBmHcVobVX777bYcUY3gm8kYs4lhtHT4Gf0bbCeyxq6KCE99zzxzTruX3
DTmcJj8v5pXbH4OukiJMKHXFEQq7TiA45HbnNHCaoLPRRR1qwicjj3GZNVUE6R81
H0H2OnmZSQ4YnOeihc23AS8Yrv4abIvLMDUm+0oWVdLUnwgcpgA+OeCkQFeKyaZr
wUSbgC45vK2/TLZ7RhinQGsP4Bm0vGcaEqbDZwlUXUWW/dQlDIFH8GHkXmoD8G63
Iy2ouBFxgFISBXe37fHNmnv48Xym6bqwOh3fxpcS1mq4DsbSIDZIHvq6awtq0lw/
vtv/bv35kfN2s6GvT7N0xSGiImuCB87rM3YcWW465hGWzCrDXWgFQ6e0C+J9NnF+
syLQ8vYnmThxq04fRC8/zp/0O+cYLeh9Lv1e26mbKKoh8MMMylxsY48/n4JJyR6R
c1gK+F2gwOxBvFM7/2WnSFgd+TuNruVS9pe76h2nPnY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fj0mGTMs/kDb/5hJbU3iz3US5f+1lct2WmMn9J5y2vWxnWCKhxTEgF5+SVP2empg
wi7G/Ot5E985XFL3u4attu8uq9keMYcsKzKaOd2PkvKJyhtFYt8Jf6ySUZiFaC2X
Bv8BZrUUfc7f0grdbasF6glNiUIbRjDn4xmypnP+rL8xpgRk1wSG0oSH/JT+bGlx
fszJsSZU6B4F1qNGgPZKMNkHuU/QioTOHolqzWEFFjmvbHADen0PqWODXbWulWBY
DgTJCejObtl8RoQM+N44DaZWZHxqjAQ24O9dE6Ml3+GkEuUUA1gwiSPe5ptl85Zo
ryoaAzFFY0BAIHlkBpSQ80p2ui0BEoXdODdVffzMdL9C9fGw69d1J3gwwIu8T3ov
RGtSznqEwd/YaWwfpPhTqeKcU69DSixEGCqc0ocPrXxO12Iwsqpb8OaYTfsdNP7f
hrfLdZRXnx8RUGY9odTzORwS88rjfBkdXAhkNv98y1+QP5Z3prKbA3Ml3ZLzW3LF
CA60m2+bs3Ig3XYh94tf9FdHLAgiiMcjt1dqPJHyp6F36eC1g10OneOQCWCUwZWF
4QzSsgrhzN+y/1QNdedzq/lS/4F1+Pc1jO1vF9u81ugJm6oANz9ecN9GyWXelKQu
IosvvOwW8OsdO3zoWTYsKZ8slhqLG/7W2HEmhshwYNXP6FgSNtNfHtYox4JLCB5y
2xUjYxcQ33twI2xwD+Xrm8ZBo307g3FiAaAcJwjDdr8xdrh7FfQ8cemsLh0mVtq7
wj1aEnPR9R1unCrtwGLaZd9IM/XCLJV/kGRlsCBWnCALK96RPPtDfp/SL9jkJaQl
ElgVhPc4PLrYAR45/v5yAFoszQqrA1Dbe/JM6CNM/6nFBoy5Bv/27iDgbir+iysw
1XiM9v6jPtnTDbnJkjzz2pkEM19oxr9+nUGFUo5XWBddhR6s7l8iRhI4nKcZFH1e
apI7FG67d0WDxa3qkgU65DaK3HHb5YcJyYYK/VyPDhMUfvCVHYs6ucDmICnghGYh
Qu5fpmgSCFy6QuKdW30aYiVRNt/KPHrqFthTV1QpmQHt6j+OwRUfKZXg++3fa5qC
CCEdBCqJ7RZBbLLKQE9ZJDjrOgmTTpSEFI17cK2iezS287JCAWBnaaxSu29r7jqN
fwpX05MQz1VypchtqLaQQKuVfdaWo3wnPwrzWVZz38sz9xn/gZxfdFYhqELwbFbc
6ikS35tsusBkBM3VP0bkqjMUivQUYsNhwLY4WdDgql4LeJweZtWH9czZ4Av7W7Da
pXAxLlAx3I3ofjtu3jmZFFF6MjHOUxUigdlcG9oGuHL8A+ZO5YC+uC5pNq2oBj5y
exv4KZqnvkC5L3YwKQ5coQOBq6e7YFbgRHTIEQoif52IiyF51uTF1Ty6IoxulDEB
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9aOQC3QrmBypOtYCVIYjGTQd8oK932Pl6sEbon6HnjGd8cZd+1xCmeZM44y+JIj
//iLTlOY53VzMzJWQ2ojBmlevJ6qvYgdXVOSqZi9XFSxxsbHsm2nvF/ONWxrjbSP
wYmjwlJUamgXarPsCVHxyZUBaM3z/L8+iIVB9XjpimH4YVhP5fOj+zMufNBdbUWc
1YrNj+cawqrwcLsdtjvsBWvCbcDFMmIVcoloL9KjmqwhTRgbjnW41CQTfwwbRAIj
FaSzsmf6+vCnjyHr3wgrghugJv4dd2NXwcSdp06LqtTSnQTi1SZpzl4OoGCG6MkK
kut0jxTLZGSdFFQ7g4rq2bHoNI58Wi53OenlKKZ2+7AvulRsQ3r1e5WreoVvTMTx
JJKPHYwdqWBx/Qps6kz9onTz120LIsTJk3Q0j3twoBoiqFMuZ71P9TKbyZZ2nytd
CChZ8XPi7UgJeX4hPeiRqe3OTEPzauxySr6zwNJt4qIgl89FuBMKJxPV0hRFvDiw
I9B30XtCnFrkfEKbkuOSEeL2OubpXS+9tN/QLXdOL6iyGKiobPUilJpSMgxbIGE8
tFoVi3zLHiESFAuhqO2juhjCvf49xUIyPCQ4GtF1Qp7x7pSJaeM/NHYzd717evn3
ZX/B2PEdQDlqCzCsHNulLRTRUgAOV44KTbaQotWZa1GumjPCuPk6avBDq5ivxGhr
TLycwrzXhQ5ycmTqydg1wDwLZerMseKIdeONz6H7mTraLQmoNPw93WHTLiAhvJd+
3ZCv2YVRMKF17osamk1WFFb9Qjpa0G4zZMQ5d2KUCaevGI7pakG3RKXPKkm55Gdm
xcicBeg7F1nuGR4y1a5ifreVpidQdQ8tikNlyb0RBVvD63Omda5+59SwRhaCVN0s
qHShd5lDWY/fJ6tKTIK5bUHt/4R635XpHAQ+QeY4kQdxLDgbNBX0Y5Qz93lFNyRP
B1kKYDIf+FnERyxOez4LYCDvazzAoKVGprGYqNcm5sSvWWyZojCfLwdMrAd47otE
qKBew2EY7NRfIkriLnE6w0GIi99YGjbI6gP1R1AxZbU6d7H0DDgQHpVpd0VMXlrf
vJPYCyZj+j0nDgipHV1Iaoqk63QVIyHPnPGPUanSwpdzyGOHEQTI26K/uiXcV9+J
rsh+uE25KxDZ8Zyx0uxq1mugr8SoCTvnosovZatf1y3sxrDaKgMz7s2/pf59hDVB
sDyQWl/Up6j83Dp0a01Duf4Sqzf6eJQPcC66NvOzR94Qwpweoh6nK1mQHnP75QAs
nx61J++1NPYa/u8g+PsdEO6n/m2rcGSa2Qu6R0SMzOxRU04Pt/jsVk3f9BndMdS+
0waEg2mf1Pre2Ud9XmVvOznmMGagfeUu+CQRIwimvfuGgGKqIgJyReRQB2hE5ExB
uicsgtiVxtKWl9jB8Vf+Hd6SBKdW/2jNzjCG52UAVIgFnc/6txvBfWaiB+SmrltP
10ko9lU3bb0ZMdysfTU047iKfMiyZbCuOBy6i2mYarlZ8Xv2s4hS86uOjOafZGNi
8zvU44tOyHCfJvyCdWkxEQDyg2Q2cvkJAi8ggt3f4ReTKRGMoFkb1BX11pwGVZRl
7weO2EHFtspQkiUDodvrrdTQitpA1a7cpI7JXncEc2UYdPoIKIQ+tovYmdgpNDTX
E74lhTVLp7ABRstdEcnO0pifSATBDdWiwY/4K0z0E4iDbaEYxcACQi4NjwN0rris
qugcQFRCdUbEszVNKOP+WsxUdBWHquwyaGcyXTMqrRjaV/3YmhJ1oZjtV2iXZJwK
dQB2lCJzQ54zmq0Oh3y0CCnc3lLWsX/7Jks3jVZqy6Y7IrCIQ8lSGTLIOvliBBYi
wI+9YOrxeglbG7qjylxF8ovsQ7Sa7X0ZVHPqkZ3cUasR/SSVYlur+wSJBWRxY3hU
JYzNfE3oGYNBJ7oaTgpcRTGb67Qi36g/2naolit+TzFoyI7AVlS/F71FGORn89yN
R6NDDd8dtoMWj3N7/q/8QRV6rHfhdxLGrVLG/Pnd1ku9ohqbDnm7ViXL9aQuDT7a
RffK8olrnCaObQSqy5Wk7S6KEeDVZA0rFNBWGkMPxsqaBV7JawPjLK2abHr4ZBa2
ukjNjs/rYZjvXk5wW2cAopPZnHwaBPWYRqDi2PD8o9Yqn0xm+JCCzpFjqrIU4Ba1
OvHYC7KOORcnLT6CYw8P/OLEHko9n1bVxhUDaOFzGdFgQdsk6cwGxflCeUnHDFuP
OQv2QNG+Il93hZfS2hLhc6cCbOCjgcf+Zgzp9E6/ZTKjqzgoo7yrPvX+fQdI2oKQ
SBTEj+gdyD2+WRN9Km0od+Xwt35ob6swKg3YEtteZQt2NP6RXkO9imOlQqKL85WR
ZWj1pPTbe42qeXIZBWctIYYrlgeJtFkJYT7aFqzUbZnI7DIjWC0e8HLstW2HYvsB
e52crzvMScH+zpPDjU3a1DiSvKZ+Up7QTmO+B/UkxLnpePdKY10UFaYH1jUfjrap
7EhRxpSON0W9RijXNuCWTU+I0bDnAVxG0q4EN3797qocGN0gXGYXJ40sOHdi4edO
j1AFm2/6ZmJS7FsvA99A4zlVJTEQnfbn0kNKrgJfmGqzID9mEiH3fAHzUqyi112D
qe+CQC798zujm/FN3fSdGUlsnYr1UQi2NkNIwUjDcLXqwgVGqwFgnpLS2J8fHsRw
595+0WfX2XWKakItO1iYNRXHdZ3tq/woZrJyRNoUxQ8rk/ZtQLDdwWgYTmWa9pXX
uD2okZM20IeMuioXCGAtWWxDSunKu1T6LXWmQINWEJKV98DCm7PBkSRzXUkxOgM1
kiaUO/Bp9WzugR5EaMcgN5UJLHwxl3k7K4hADteImCXIzw24XlNXu8F5VmZZqvTo
5/p+CTDVzKhVjEkSQWXIpkCo9ZWEUEk0/HQRdUOWhqv2c5ZvNPkkBucMQ+CW5YQn
6M9raTgQaRnPvG6yL1Jsq70QDXiV02QMbGXom/l3C66Bc2xf6zNrcARs7RMSaTCD
SE8jQ6hSLHO4mNPeNvIOdB82e40R5CUIC5aMa82nZsk65fX6KHvTsso8EPSI8nmv
xU7TFZlbFGQYoYONwDQXHy3S5kJ4RCfrCwcQtQQ1HiuxTf+dFW7AVdBj+Qod/ZCO
xEzpESagdFermcBDlUXo1pA2+YcIvLn7abAQA6xGEq/28qSRLh45V9K7hIfSPAWW
9DkeVE7cpzPh8Zcqtas7WDhWhHcMPZAXAGmffnbpetqiubQZvpzo4nCAYKuyl9en
uuvpJzK9qHmz5appoQafUIuJJC1/0/3jr8jm3Y5e3j0xqLbwMHQJb0qjo6tDz2h9
8BCQvkZHENyQGJ90TupyIdsKcNI6iW7315ADdhzTtEDGP7sRm8nty7OsM8Pxu3Dy
qaEFsNPN3R117vV6JLREvWSROzJp02jdK6ZqRxQd96aen15iEiWeZyf7fT6KVgC7
WHxIWSQv+AIUqgsdRe1IARTcb46Ejm0N5xRoWWCDRnoGBEmQUXerq9BFWSpKvdt+
PvER+h+RvYEm1aaIpS8ZSfjhZ1EKw8xLN6o6Id20d65SX9rQSSQri1cxgvRdMGj+
5XqvjiOLuSfHnbWwbLYv2pqDbR7Z75xvliH5/XbDt5o7Jrq4j8zCG3Zx2HAUflqr
zJAs5KOtn6WbdDzRZ5RiTL+bwevUZAeTNr/XHYJmM6PF+THVWaj0lPoiJFzGBZnR
Yo5gvh0J6zYFf3wkcceq0c+ZJDYRtm+EwtNLBOkOF+AnLLqjdwZoIz2p3n8AIyOB
zDukDUwO2PKx0c8ilV+6c1RUeSrd2Fe5y0TjJWP+LL6pU+O/UDqhbEctvEsgkFWc
JOV7b5uq0l13HvkdB6hkKh5ucNPoxLg0S69dXMQdUBfjqqaYWi4yuVHMunFviyIP
MNt/KooM7PfrVvoi8JHJabMmyjJnOSfJo1e8gjCdw5AaCd+LghSAjmCVgsMCo/ij
sE00JdRzzsGngvE2EPg8g773kmcp9nJsyR7C102KkyrSxPQoObpTvjoYeZ9jAQad
lnXc9BlyiAGUYwB1g2W8Uv97LL3UDsU6Wr4baGi6JT+KrHl5m3uyIWklsrqziO9r
IekcHIYMyKFfWTkdoaDLdfNu10aIpP0jYlDFB77P81XNPej7UW5raobVpJjVqLlG
RPLxdLw5yCLuTtN7KBUvWivcpjPBWuLXw09I5N23bg7IHYY9xMWKq4KUWeRbTZIh
PSMMUCaV/kltKqkiXILu0EJ6h2kIaAbB5pEJ0tWh173q7cWA9OSFAswxcsojbI9R
ewlJufATn4e0drCLhGfM7g3YSFBuwxyovov2vn02t84QYe9aSGbknSvqX7SbXNbX
O/PaHgippd14V+gVfOevHOf+s7LRkNvPGQZa6t6Vss02X8G9W4rZQX+PRKuX4juc
HyIIfezaxlS0cV6lm5LQh4Usjr6DRMdFTezZu6Za2kfm06Bi145u0nM1qSu8aWI8
m7M7FOcqJ24Nh5VREZEkP6nTQOOmBQ9vIZYz2rzAlIOSYReSt3BCLN1h4mpW7ZhI
gu7XKMt0WhTN2t0I/a2YxQwkzOisr9CW4u+FeOQmVLCzjLYTBfI0NxyR9yaFgAVW
v3T5k04lUzEPtZvDhnwdEaBFAcvUzqc2hmujgzH6OWkysyYm3/06ZUsYh3p7tZ+O
Umn3918ac7Q7o6QaBrZVomWR823OtySwm3qOzYX4l9ch7QYEZP0LGeSpxhomcU0P
X2/ZlhpZigEttOVQOvowagwevPkXu55VCyYlo+z9urs+wo2FNmgOMPf1EyUL50Q/
kT72/04jVAQL6zIhU1SjopK1QgSCi3rhNIDvemLFxqZfb1bumhFfO1LUJkkM5VF6
oLligth7V0vbOwEBP44kMqu7vEi5KOPxvD6SNgIY22IR+2XVUi9OqN7sOzekDSjK
UtJGuvsuXjAuZjp88/Ta26DmlM2RAoxKumQVqil0pPGpfObjN2/vnmIf/OAeGwG8
DoZZ6jWXKD0Rv2Gcn0OPOP1MUX8DBzZUBrwH31Npbxlp3YRrLfMMKuhimpdP4sc2
+ZIuTbQDZdP+H/lsmPrfBPSpe2h+3IGF4DD40O1DAi+sWmC/uuR94SJcoijXAIyW
DIZLaweI3THihfQ9tNwWwjFDH7BRdm9kFTVeGRgCvJRvLu4ENsOKpf+eWm5/X1If
3h7sRjkQ0dV7AF73pT2kUi5w39iQy5W9PJbCVpMIlZ5stuC6sH7SI4lGzGsUml/h
TdMouAeyXC5flapfjGgVDl5y+T+XHX4ZlGra24ibzhci875U2dHfruP/FtnOVqlN
Vtl7nmRHDAke2VZyFz3JUrAbN+Oft791DLFPHp0W7PivLRaRBQWVX2wOS09xaAmy
+KtV4SVuYSpT60/Gvdc36pA7vWw4/G2/gU2DxB8w1wuKkCGozn84A6NNkNADcCeu
QjB/y0ij4ToQ9bkfSGNGLjWebCKKy79fkVBS6fhDKd3UI+c16qZ4913QIhnm8XRU
BCg0tQwuZ+kEPXF0/P1Go6zAKHkF42xdgc+Ep/1AHRH26rZLA58DZmsbvs86fV9x
tVk4jokWlJcHKbG4ptbxU1JXFULZR4a4aeYqCDHg+xyTOQ+s/PL6EL8oGoaVDO2A
bUQkzyDP4GGLPh6DpOalZ2CgIurQSdKmp0/tnS/lzoFCDah0DJpU8oRiwBG5dbQb
ZRItZI26eV/tmFRa14443pY6ftccvZ+2cMMgFNmect4ZFJpcpqfI717jm3PUS5XY
oed5SXVjqxNXyQHmOTPNFSw99bj68L09XG4m+lbtpjNMzvpyJA1uGhOMyUroEHZT
1BxipAGuQDQo2EQ9f9W/Sp+PeKg0SBY5gqW2cSMMopk/BOcbD84l0kSYYQJyykFc
ZFjRkwnmdEeDXHCgiP/uRCmePcG3ZUT6ePQznOESv5U4F8kubighBzH3ff93WreO
NlGhdSQXeqR7ZMNS3onypAbws0Ib/zvbabWkZHS3xWeP9QmcPVzFopja+YUufTYW
Bn2C52N2z8MlalWI72H+N6ZsJbhrZoJus5LSAy7YVbNe6ehdEWqHWO5P0FQs4uFR
bVrOH+MMF74o0UlO0VdU2gNBT/ZglpJdwSWLpK4OLSmNHYbBnVl5HObx/VlDjxqf
ebo9cYGjlhK2vXol3HqGosaEKNAGbGRO32Wa8VyoNc7ekNvSSUj18uIhCWUc7qr1
xmz/87WtmTQh5LVI1XVDTf5amF6MNxfPqY2H63j1XUFfvRnnSnR+TtQHu4ZOY/3B
uorEXKg9Qq0Ze1PFQH4qm4moIhrm6KBddVw5UrfdRta8nIZriLAoVoZLwfFm/9lM
zPSAYx0hp6cWwJJZN6pUIDpFzDA3y+xEUgEG94QxWX/9TwcxQrSbPJL0UUJOV1uf
peYZBbzng5osLFd4YqEMAZqTaEvpqH9Rp73lQ7V3EfHeUIkhdoZwavVaIzMAXbt6
V/Ea+MC53O1QpK76mNbR6VFncxfsENcW097NYpi72TnXekazLxlW8Y0zBi8jqwqb
m/sNzwjNHdilwfIHpzKEHoOAIdehAUgPR5QXEFMm3PFcgiaHEV/ZOMPAMJ9ZTMRw
iWapLwiFVksvO0SeHZEzqEFI1u+SDw1+yaiFYww0GduiQnNsxyKY0fq1A1pJyfSb
jfd9PJBxphJQcGTFFOgy+Z76SrPfn0axXs4dnHTXaewCDkPriSm/kE7nwBF/iuGG
rwLABCPqzMUFNwNBzwaZDeTIe9UuI7cldafnhULYuBBJqIoobbsz5vy/CJtO58kL
NrGv9aHn42SPI8y121FNsa5BDVw11TAAFHzJza77CNMkcNkVmyHHgx7F05ucqexk
PLqxSMzD5a/FeFrVlgzUjoCN+R+5VpLgYMM0RNvhrTvclpY/YVZgOw+rxXTkqv7R
GbLb7R3ayqz/dPr/3GfVdS1bG99PZMy5gmCkXfaW0z3Kn9jK9sy+x34f70nlmzAu
xXlRRxyEdYIG48X5grNIOFdb6ngdhjF839qcZOkpjPZQ7263b2YvG4IRVzrRKu6e
545BpujiNsW58kslmP7FOwD8bZVm6ExneMSSg6ohWcsa8Cm67AsrMgUmlDNRqJ/+
I+TRFic0vx3h52m2KxJwiMMNv23COQt1zQksPR0+phrHNyxqSqd6bovUU6Ofgxun
jfIeoYsQZ2UIN0xQ3JvpGaA4bAtpp4LsageNi9FUfYZ2SqYvKg2ljAP5n0Ebenx2
ZFR2xh5sscWDgLTu++qD5UwvCrL0PEJk/XHQnK9HdVD2t9u5J+su09WmUNLstMww
2R1ioCKsLwXVZtQTV3S2I0L7qcTbCqEF89XUvSzl4vqmH+ETOioasYqViO/wvFFp
0eoPpr1l1St2kS7naAg81kIPTmwOKWgerK9sAlrcTZde9u0qdtC7eS5C5BTC4QmC
ozobbMcB74l1aiDkeJoeP7pqbc5d3TtRT4HEF2lOK8v0d5TDPUfnV7FmQ135mfOY
CtZQV+lSctq3DemazfBnB+UikXIiwOliixLBhIJ9rK5yRA1dVqFujpsmeqe5evJs
ozBdi30HNl5aaPwt3x2g9L7NWMhVOi8PIako3fc40h4EM4jzJQ01zKNkgzQe/uB5
YpNq/aYRCoNABW+I6kJVc5dJCa1dusvMxFlmgpZUe2cen53pXfscQDDQgQaRcyqq
or4bINRFYNbyH2ysvzP0oAKSCU7rDHQgzNW0MH799GKeWtKjfnW8MWKk6+GCdEJ1
9hnvoAMHbG4ZjkL5Zmo8kXyIfA5dXIPjI7J4wjm57YOSKXcjmwD6dNk/36tIQ3UT
LHoyncih6qVopYvuW1sh8qVflC9aKkfshHOCz2vl+8oLt5KMPvh1do+YhGDFajxf
VcRgm0WgRZhbPNuKIZ6+PyuxWEfhnyiIlT/qfhMBXW4UxRenHevwqgasF4NcUP2G
B74+HPDQfMsGwnspFx+KUucBiINfNLsFfTS9vcYcxMc9UO7n7QmOCktkOdikquhs
BlDB2ry47y3dDDSxyFmPk00ekj5z1l/dkW8iu3/luYOfDdfUbHhLnLacbxs4TxrT
zARoHAdShq6PIXhioi2NULluy4teoNuQCNxv0/4AqIIYB0F5JMSLqx29wvo7GdCj
n7v0uqkc16pJ/yzcHxsTh335h2Hn3oLSBHBGzKrHkhKeEZvb6yI0A8E/XLTVp+3v
gnJtMwVpQyU04Jv4rqnpHjJN/yKd+LnXYljneH4r9VP7Mjwtfyss1kYgAGebCMl7
Ouary7Jt+YNCkYTqjlE2E7vKQs+jsAvOP4nX88xvBGz4SbDYa8iOb6tu9VIZVavS
O0ecs9Cz9jVAmBKzyAApcacmgBeY21wOzUN4gQSfkowIQgalqgh4CoO+34SjjIBJ
GR3/DgDCjfFNM0esz792b8m8dI8pPnHOHOUzlBIYiDCRUnM2ykH0ZC0iuSyc8roQ
/gxEs0g5EO74byFNOPqwhsx3KHhuWYBDL2wrvxwzU9VQKToZMcwZBrd9O1JfkzWg
oYDN3/x+LObojmXGs+I1z2c47dVyIiBcSmUZAbJJQDqk8ESuYono+FN4I0/F+V+l
qPV8+p5y43Br+/i8KRAwE2MCgWY3Oz08oPoi+3hGe+fQNaP/wnQS8DjM0v1DGwLF
XCzQHjvfuqqUELTpmyJWY0FVmqR1/1NcgrMZ2tBpTZBig80g6Kvgrn3muB6Sp2Xe
5gWlZlzSefrwrPW+AbU4FY/icG1ix+yHZprRqpdSttgNnOkRgCD0kTIPspMF5NDH
aGmOMnD0KLHZNqJqqmKTFvRWyZ457Vu0f8WkbewHoUv1XGqbgcZE2DYauf20+HOT
bjA8YaxiWaPmUTmqoOqf3QsEqIhZtM9qrWSHYKnEzoVCdhOLRL2N22ZD0HLs+mu5
LGmuV9FQxy6YJXN9gi9cm3tunrLdEgj+dDB4SqamambohrjmbU63mv2p+GeyHrOF
V41hgrvNnvSRyAEkP4KJA9q48Wi0gynl2TKHuEmxsA+xSAowwgd2u114kbsOH+HU
jbQxUFbP5vMrUTmMg4uMLqLBQZUD9fXjQZYCz+TAt67QBzA3b4ldvX4k9kWG9E6M
iCMCZlsGwAxdkN3TO/kFdcsm7cRnZd1bZdj/9LEiJx67+OfpCYlrcRFO1E4w85nN
CuRTtfYqDQnqF/cYdBCsHOu6mM5yMMRzp8tbmc4KFND1b7016RjgOa8jZK4iZJpw
XijxmyIKT5E/1KV8xIj4zN5pG/LipzdGeC33nZfSbnhjP8wVTC1Xxaz+cvtAI7b4
OftBfzSiuRU5u0hUMYf16F0yKsi2bXSisB0PiODRVhxcetVDZp9UG7JvbDqXhrsT
1vTP8g/W4nQvqJsVzctYaI6//EuMCcsPLbbXyPxi1I9o64YiUq30mq3z6CS6+hX+
S+wIY1k3tqvgyiRYgL+LOMSMi3Bm1akfWRBjLDrAh3yqhmtTVLInAE754semAfa7
v04/Tlsyvu1lbrtTZhvAvbQxv2LEGgwsTPLymVPqfAoComIUhkybF1nDmApmFXQB
Ga6C+xhlFq7jGF2oaJUXVFqKMW11KTgqVh5oZeWEP0ZsytyMt30kl470gH4BrEXF
mJMEgQMb/kOpdR32lp51rmzg9WaJauEgAd4WYEGkxngNJisE56a+04DWyM5cy6/K
9ol7oQlQyDiVAMoE39UR5tsfOfVcq+hDQ1oR1p0pxtZhwME5NzP/duTZpZ7mY+1c
ka0+Q7+0B9vEaWSlMOko+VasEIMbCNXUVwHDpxgf9kZcASs1TgjrUdm54T7Fl6EJ
K5/HDc1Z6JXKPFqdrpC0OEi4Wf734qm79esvD2yCsgIgZtGIf5WsvInq9MC74ikn
iAIgbw22zkUS62mH0FxAXtYs9Sk9klTEAN0ssUg9Bq+lW/x+O4yGhmND8iqeUHST
uhph/dmBAIW5BK16yFX8PtalsBLN4T0cruO8ixeWiUQ6d72FMQmrJ9BjM2/qxU9u
ieWGEzCQENm2dGnzAb5rol86rwhSC00ya1zuCUq+fJnjvuY1obLJw/3YBnBlT+OQ
T6MRI6h27a48NI2TrZ2FbJRJ6PbdIKz/wMkxLbmCtz4ORUwmTYxIc7cn/aEe10NF
bxAqyhPkLOvrjNQui7xfHOmLIen2aD/6TRZtVaE9mXvHoxxiwCME2Np3xZ7eqUUo
HcMO8RBPl8FjSsU/vuzet8J/5pVxqj6MQ48yscc/Y7OqrZq7FDPW+9bOu25X633X
OfbDLNZ/vCn73GqzXUaR4aDQQC4Ks0WuRjwE/LvBUHTql16AMTWHq94Z74/ZzDAh
Muv9ElACBV3cq0EpVEK5RqY4S3tHtYYFflJYiVVobR62KX4yiqI0eahfqeMR/vIM
K2EquVOhuZ4drxQNfX2O4auVm8ueopQcBPos9OeSPKezvAQvfgAtRXjC7g0ES3cA
FyJShve11813TBCtRj5CR7xCWslg7Tdd+oXJFd+XT17d2EtwDxtdEE7ds1tin4KB
5TO/8aMe87gTB1jP/8xqjdN/tYBVafmc8tg1cJvgmr6hDs7qNG3Xo98Q+6xaZZf1
jS8mhHyc2/5di/CEORIN70AV7gNT+JrzX6x8N1E1ZA9T2uXDMqD2ZBNLR0T+n7UW
fYoEcM8acWuwvq8yjXeCvt0KMUcxe8XX4BXlpnBBwnZbOnOLf23tH5Z3FSof4xZE
ARZsF5QV9uzrgV7ouNRcWeOXE6ZYp9j3cCeLPT3wy5WHNJT9yk1scZ4K/up1Zxan
JHXvcFaL2yjVMLsIPApZa5ysz8y2YYWNUyajcmFfuzRg9jXS+5cgjw4LbjhqMeBQ
8O5vtdL350YFm0PIPJS3PZqHXu06/nMTVULFpbEFBoBjGPyJhPckX9QOf1/KvCBq
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVkccnRfAY391mNNCeAev/HAHQDUxt4mskTvtGjVNkfBU4zljMAyeRJxHLN0RQCJ
4uPqiMbWB1fNKr8U+j0c2ufKiwSiqX7+3IeLmXt77Dn/MMZOeI84lk7l+uKbqWoN
qGcwh7/IJip+3VG+1YwLpA8ntTLQ76hp9WiMo35k/PQMLq/rmLn/heHY/81zWKzf
IXr9px2+astFT+XrNJ/CqXjqaEVO5mnYDfbCcdxYnWgIg3IbKQZ4vspk9voqm/6K
/6EXJKNJI+QemL1puD/g+hwbVkRTjhkFZPeku00zbMLDtSKM7gg2iKJOgYoqovvQ
9GRoBHsUVomVvMH4I48bwafeXkVu8wqBYsomYig4Rveo4JpxZ3F9ZBTBd5S72aT9
8wiXbeRdPGUgFtJrGVrAwX8wRKbtDeHpzQfpA9DS/IV4DZ0G7o+Rz+IK5gLat1Br
LOoW4bsza1RPPBceFa5NYg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkzJKrdfJBtN7wuKY8mm6bkSbHQl2ndKoT34ynXo4AZYhBVpUt37AE+v74tZpx21
7WvF35jNkCdcweN1qFU9CxSuxaVzZEKjtpMs41N5M2B+j1IPTbp9nDXYW0NCLUw5
V/KtxvbfsaR+eucQ6MtSD4G4OJUstltG3DYZkTY9yjRdwO0bt47+KMWpehoRJrLn
JKq1KSFs/q+YqJX/5oYm3a9ub1xxFOm1qe6jSb7BS/Mc0k8oyRRS7f3bmq+dH9pu
JN8ibtc7owNPoBTjw2UenPhlFls+2nQq4FdCukxvxJZAyFoSJLmbH6UoKnSaH0Hm
NGxPYhxtRAtCFzqPPaKnhHbalKU943oftkvvfKRmjrwOia4trRFGTsEzVMQkBffJ
HQCCnM3nSFL7ZfRt1sTWuCzxF0OxRz6DgmghifjyLy4V2Tjcg2dx75+IWi9VrmMy
EQhZb0GCU9aGcbEPVl/BmLTzZZha8+Hleo3EsxyaIDb6J0JKfmLQZvHfe8ZCGCT1
0GQ/ZJ98jOn5to2D9K7vxTr0tJTyEUj8NAa5U2r8EMcf8/y7wI8cxJBkMx7guhvY
JD8LLgEr75I5KHNcH8HUBuT4p8jHs2TNwVKCBrWRt1GKXNvveAfJPCXWRBImmkNX
eoPN8PyaqyhESpXROwKq/m32DqA45Oyyl5fsl1tVQKXIswx0jOQzKWZTq37avEKt
cdQ/lgyfhY4agZ+qmMN0+CV5UTpXOZCwQYadIi9YsT+1KtzN3XrJBEWEIXeey3+8
ZX9MIfugnkZPN5CHBUEGc2wkxQW+CXxoLrQsh2c6nv4fyT0S6rP5Coqo5xM4vNWM
WMOF4moN10shTcFJTMMwUztCP4iviY99cV1l7Cic04JwvJQTqQTJAiLjaMypw8S8
A+0+5f+GUpefzKbWmpOHG0YM6TBMW7mSGjkKufUMeImLK+yvHBGML2dQFpKiv6bL
3KtTvBgcJ/A7Z7xIk8CRnsIByIDLy/GeFNV7mrXAI9WWqUygr/6K5dw7W84pTXK1
5g60LjW22zhlXxh8W6O/ugZgmmztFIeIGPScGLZdmQU9oQa8PTnPMrUu6Pt1aaK0
wZq28+igoV9eA6pZ4lrC/OJ2scY9Rv/U9sJYoQGHza1smQmg4mFt18sgI83jdqeM
rPHyGN+RXOQBaLgavzRbcBdz8psyEr1AKTi0zS4ns+fbbwzG/rD0z+gxWyJW6MKW
5az+Ramx+WlneiNL49PicHgb/BpVaQKU3TQydH58HvWgoLDz53s+wLvbnbWj/c32
mfSknjyA8FC++lyGMAozWJBmhRWoUZ2S3eIpOWdvD1SuhODczFJr17Zjf6hJ4faE
w4c9K/GURzFreoTgSWZbIghVeStLd9c79yBE818k92KEmgnlISvsNE5ZQ7IIplrd
oeqakqqUXCwhLdyoy2kVzSCvrbAVdEXWZpOSEoICCvmiKBSL33uRc4LaIKoapEjW
iJr7/2xt+ABwxmnAta/b5bMf9jM15gHcV6xJ4RurttDcH7KMq8w0DAQolHqgUf//
7PtFEzCObwKnwQPHa/d/0xwiPJF3btr5dQ/gArQWUJQG46XQv5FIaT7Lywg2Mb9J
JxO0DFilpSXp5IdVzpufi+MTOG1rF1ep9HmIfBhD5x3Y30KA2FaOgKXC3cdDjU8H
VZw8i+50BgOjrVuUNLPUeDCeWyK0h/vN6WEtizU1PARjLjZRsTCqKNZVq5mGrbYQ
yqOkfEe9ssw+ujRh1AvMZWB/nBhrp6j6R48aZk6tWNxVLVxGrPVq5pyX+xI9734K
/wHC2KYcD9N+QVnYX9UM/znt6JiJgvj0sD3zBHmL9MPKBJHsQrvYIi+TkBV65T/y
vs89bIuI3r9wt4G17AlMAWiUwb8TqnzBEQSKqXz1bu7kZ9nsrh3ev9PjT0e340fw
H8BiHOpHia2/t9BTfzyYLNi3G2kuQqg4McpQwiuognj2TDKeqFIUR9Qct8Kq6Pt+
g3a/j5X6gm4a3aOU4FesZSktMNGFO//Gorrq538YVVKy1+VuHJeKGoT0RSwz4bOs
nfyhXTjNXuHkD0Gos/FBddnQMl0CI71FQ3f8a4nF2lMx/5vW3lINDyuCzVNKh/A8
I6bukiFR1h8c9inTjzxwopUmA1BT+RhVDEkfWdE2ZHR+1Uyo/DHtUPDq1uP/h2+k
QgM6HfJJLAE6UBlPVU0xjeEM2gRr+JPddeQsLTF2pH4wGirMsYe7uDzYl2aTXSG4
5419LWcPYsL/09U6nA4bYzLzmuBqaNCTqlYJaNoINDwcQ7yEIiskpj4bYuyWrpZh
rkxkLf7/3+W3mrS9UKbKpdJ5Tv0/EqHICV+UyPlSKmuflkBhToeSP6NHt5guxW8q
KiUn4lOk0YCJC1ZUZcGW/6tjQ1S0/8RgYsE84hJQshDvHYV1EhHZ7R9mrhG/5nUV
V3od7LIo+HCrIJFJfEmbe+PEE1+p9SBF3c8+TekQf00BSoXFAbXrqxfHlpQhxyrG
nx34a8tSHx4b1SxFe7cdzHf9Pn0711iVlgSTFgTwuweV3aCM3za9XOtk/+nmhn6f
R6/D8UBZYFPS7l6VwN7NY12EwcLutEAZUPal5EumO51XpcALTCZXlL4yagcII9PX
2gxbVBSC4F6FbXzTi6zmeZ5MlWT9TGzHFj+OBH9JgepcphckVgnGaJUD+eUt//eE
XnuAQNStvF94u2HpiTo/XtqWd2YvJQn8rhwuyZVG0ByOsANP5hRkLDjbKy/+Boa6
QsFRQ2V+whRLGydz3OmZ50LLJ/Md0zpCEcRx/eEmnnG0xKYRL6THJkSsXyTscz3y
caHHGPLDEWscTZCGb7zJ1oP+4MdV/aN2JGjIUDO7OdPIsnIqXgHvJ/pao4TN3Z4q
FGWGAA328E5THTutVLPIFbgZwGG1OnMrCc402iSEfWhvaBCRzZxT2oRRS+KSTkt+
hCzqlhMU6n5NvzAoJiBV5qeZaMwgo0xz0EBiEthgr7pkKQDB141QjNVNz52qu7r6
pH2Vdd8jPMO11mCR+XOdv3FbmEWNk2tx9xAh+Ec88rNrzP+GpFgwAM62kuKAS//2
b/9ULzIrsJilSP1s9mKwx73NhJo9z8SqIrfIsXVXCnFk/qBn4IbzOubByJ08BIiN
J3blJyh21NVL1tivB3WaLnISlwSccl/uFbH/4Mw4JH6mkl3PSqFJnVMVmDm4eajF
NvEhXOft30rf4QK3UgCOusctrEmVYlJIwi4eCxMdcQwpCXNElSZoe4CtW0G0roxd
hJvtH3i1hcM2wOXcyAuGBwThkpS49TtqJT3KApl7OSNBwYaPz6VMHdxCJMZvCBCC
RaDp7f/uZZ3KVzFK7j0oruPvVVd1PeLt01vXouTGawKzZkBGXhceYLuvYLqz3t8P
Cj9oqFueJIIDTu4T6cnIBRL2AzshO5TymZ2ISBzuIaZp7fDr66oBz5Kb/Kyjz0y6
NRCyR/ypKB8ZLvR6X+93byHt77UzIBWv0j70JZSOCD5pkhqtLJcQwL3xKsBJ8iCs
/eyiXnFu08XPRPP/mEzAXhyf6JwOtM1w70AGnNCYXrB886x+8iwHV5UMPsMOXKyd
8MNrJzM5j/C1mUKBHTUBdfs3asG1ZpNl8Vl4vYg4xGw1BR4xXF+8ro+mhDd3FTnV
ICPIhecYqohQDxkt52OiAdyqwjx/zKs1iKNBUGF4kItR8ZE2CHi+mq/xOuKWtkje
L72pcVo7eqwPUkT9Ckxvta6NE4KUV2arGRKosBe1ussig88jtfXyvgXPdj9fsWHn
wrQ83Mqy39Y73w/f5/4VWmorDrlFLvgp8/qD+6ZI0ObzL9ule23bJoYFXH+2EQY8
HsttCPhhMcSUqGSC64Ckvtrq0Umd0qTYx4yxd4D0iq0howEY/7DFrk6+Md+yzE7U
fxSnJmEo5YZp4uwTRBVbUiMd9vCmbgvvcCrGt4xbk2lVKHUzbJAeDvgFhjOYKUZP
R2EnNK3PWF6Qr8Hz3fw2lHMvAAPPyhtF1/JDhQEW1t2e/mQzCyMwNZzzeBPcEii0
sCzqqcNZcvVp8/r8e8GDsncXDHqZO9pvZiJAhzKDXZB8Qo/RqMcQuLw+iYVY1r9s
gJZEi8Vlv/9cHQVVThXtVShghM3yp2qSKlp06NAxsGmA6GUUKdLSEg6js3XlEyt2
x0vBK3br+r5rsCjkFjLEat8/d3m1xA3U9pkN5wIm/CO47Uui4Va2td4m3IJHNQAK
qZCDZ/7Sjx7BrHuWps2W4i/RMwSYjrO6xBvLJKainfGMaQOb7m/3YrlX94T5LFC0
NNrUW01AlcMCcLZIUtgyTs1qaNh+OcTV2mfDkf0cj+Q/NEz4jmXT3NVAeo+FI8D0
aRdJmWWt4EDxNLuWZz4/L1UwWJygIgSFwMQr9iXGLwaGFJz+CnfaIxuYQ/L+Nob+
v42ddN305zLsAQGrITAjgJxgLlwz61fGGPMxdjLTvnOPUGCXaJAICCqgeNAz/Iqt
czrgI7wQKqd5Bh4th2x+qSxRY4NL60m5E6DMecteKDJb9EAweloZ6+XGutbwHz8k
kPR/6HQ6XOXFJP4MvYKHq0Yur053rHhJg8dO1Lu0sIH4TZpU0Mchmzsd2nxyLqyw
4gX7DdB20NDEB3qFTUZNvgcAmr34PvExRdSxywmTodcY2ku9Qv6a98xqy60P+p02
5NlMXqxS8us/lgcmUACNb1L3ge6rs6UV9kPf4mlyf4dWiCN/2MH+ToRlpPsyAg3n
P23GzGUeSe4Br/FoaVV9KYmpZ/pZotjtLeZpo9JLMO4o6GlbxxdqVKhDBXYkUI/L
kvoHaFTNjiuo8UUJpLum1wbR7bfieViEhEO3FpP3PuBQAUrOsFa1q1oIk91zw3lA
YetNC7QUWWaLWu2+XFLLci+T0C9F5R6lxlgg3Zrmu+vciT0tNbgHzDVb4cpDjFw3
1CqZgCCB53HPuGV+hd20K/pANhjWd8c39eA+q5uq0oRyMABUd+FAjboqD9/tHYmX
ex8DVqY5Y8/bZ7rL1uYTuANEaTKD8Yi5J2LmL7dao32TEINoTxX/C946dkZEeY83
wP3LLUgNPc1KqH5gIyPHsnKp0Z6Wr7jbpmhJJTD3b73LaAKdfZXthO4NJGZojtrJ
ENY12byrnDrVZQeHKwQUC6m0ImD0IFUWkZM6NuhXf1BkObgX6wQ8zX8nSTFLapo9
AoeRHerWMB8C4wnOOL8k6gZTeWi6P5lQ5QV/KeiEXpqTv8qjW995RTNUfcnrJjno
mWhkr+xb5RHcqQVEO+zidNMCck2OeM3GsasyOeZaI/rrE3+7/YLXlUdei2BW96NA
UGHmAzxoY+6bF+k/4kTCK/MaiBD8MPKfUqoRaZeJDz3FoWs6MDMKZCKjJHimO25I
cnqL4YIC/gnxDoms8yP1GnnVf4GNCnSmIV13I4llW1Oz5PF5XWR99V16tAzQ0Abv
KV6kClVhLpLy9HjdiwDuN7L/RkqFQZR8YyiPJRBhOf3BoDH8KIkcQ08wGqmiCt+I
cpIt0v1RM/J+Tn/GdbzaXrgSsU+r8H1qu85EO+5JK5OFzIU8KDOp63+LjGDKlqkQ
h/8xl437nr9bvrGZp7lBXtnyNgudfxIPelCvoq879ae+SSKyrA3fzuZg7mJoKsFs
YbcxHIi4guO2onP1Ryl/Yt3Av8vr1BdTmnJQchqE+8FsLpMPoUUNEVGuiVruJXPW
LazPGWlTAhLKlgIuqhqQcuSdP3zKdryPRMwPwkIOjnS5DXCTU6sNaWUa+2lCjQAD
eivAw6nXm1igLKjM4nh+eYNb0KvqxfpnWd6QyVZq4aPOLmgvz/BvfGXp9bcwqUG8
X+mFmXekgN71AWIovt1wLLZXNWNzqCmCO2c4wj0Xv5/HpDrwG9hB+HmKnKurDA0a
iek1v7Smtthyomxfg41dvkOMbGx5Ss6uT/i94MLtLzMcfc2A9+Q3dI028gOLHdiy
UhfhTAFtEsab0wo0dbnb6OM05b8oQBjBllhhDrH5i91/8ZehUOexQFCgRt+SfNZh
DELvLSS0BF7lnn7roAF44YqmmGlYkJTqrKZC9ntwi/OcTU6jSjxa6Z6ZU3RnRqnT
5iK5SDjFA/Toew7TmshzfjenASMpv2Y+ZxG6zt/UXIaukYwOp4QOFJeq8wxiwmac
I38E7I/D0Ova6o3dEkhBhXg0uq++c1y2U08ynTt0kfmvqYJO6o3hfAFRMtDhu2u5
w81s9CGd1o3RbtlKeF+AZxDg2I/peQxNOz6kEyxzPCav3Fow2okOIvsuS6QLQIS0
rjKroMTOsqubl1QNX+yE6pVsA1cRPjuiWRXKllSpm1P36dHNi6/AZKkTgXONFmEx
2waFaqU3ornDryLySiecaNma2QwQKlK0e3xfp7LWGF0ajqvp9GesUInFPreRn8BB
muzYgXYT5z2OpY9kHUD4Iz5CpgD5DkZCSJS4osScpaQH9jPd/X3JPt+p+3sJX5W3
DwFbXFhMDLkXO1VUdM57lZmZKRFIHi4oPaRVGydlAR9q7hN2jgAiPCJGcFLaFMRb
W/JlSOXNHJP8E/gIZ/Vz52e2Ey9YiOxv39TLeLZkSPriM96LRs3WPDuDLub9I3au
842cCNZ2v9T3AyEOt57HgdModKbMw0RSxYKeqw6sjmCatXDaCoKathwdnj8eecH9
TRMmlRAIc4iQRPOWkhirNZteEkzKNUAzRZgXFThOWUTOe8lh1iP90Q6yCc9KQFPk
4zYjKqoh54gsufEHQkCliaHZwOGUzrQCWFdGotZK2+0u1kAqTiyIMtUANu6wIVWC
3EnGfgpd0W+KBa4ciDjGsqm2FkS4iwDPC0GWVbuAKXtd4KQ2L9FQ2SWupbse+17C
6NFH1EnhOveu3eC6+psqDM0Vvb/1uHyGZHGDY4hg56/Nq7VZlZbkrPMOl8m7f5K3
T5EyBb/I+xSKAb6M5JJY36QkY9ppyX0pfRtmzgVVlMxseKTm2rwyGQ/Bp3gxv4KY
MqLRq/9WoZ91VALFkVFItfXaXairmOOP0o2yQuzSsffqgr4UdS2/iAR7RkvQjHE5
nvPOkLRzCEe4yW6Bu5Q4yhNRxmGb45/zaP2rOr/jIveUHT6lHh1BjquphxzH2yPS
gXVPJAPaJsLIqgW2YwbkHQgxCp+TCzAMUuIfgkHcY9HNCdX+sN22qcVJs4HiiyNq
xqz/FKscK4122Nij7CdskactzKLM9VMtndjdYN7L8Inx7ZS2YknHGilkZ9mb2TVf
mgGYUZdzFOqqM7bgVK2b2n//j8y7Ad7/QToBNkPJyYLcOjvJnZkHFJWxWTIxoaFb
OXqZkB/iro35Il4cJytXX3CMk7Hv0vW8Tey/kILnC3apMExt8yRgesX29KA28qtl
URBB0YZAD658JmxNDUTJgnG8bP/IpGTtHj9CXeAfMKKUdkzriScdcEX4P9J6FyLS
y/vfQYNaa34BPsQMlNvnB2Sv6euvVI/w5bK+JOACLiz1yRBlPvdF+GgfJWYK24Mu
g2ysZBNkmeSvJZH4IKXBd35rksJFhNn04m2/ak10vqegZUrVN6YicC/N48FTQNX3
i0zHpHVxGmPHSlVlzgYRiaFYz8cIgpdsz1X4jYNHhaR8VIXDZ/khyuZeJmydYNUe
IqUpMbgCNbeu2VGuqhiw6J/7r3xV3gZzhXK94v/CjO6HdHGrybTwXPCLpRI1Q7Kv
ABkzmOwi3EWs/TRzutTM+/QLfTHI68DdJqxr6YXNhPzArFa/9ihuijcdlBPP4Ora
gu8v65FLWI+rK2oHkgvgOTpLTYceoWiK5S8jj5IxAVKQ62LsVcBwZ6V4TpsUV2B3
n4Bgmic7EtbepugTs+msGiyFrxaeGH/Rj62b1KgRSnY9hH6ByYh4GrlRbcXE3dHU
RP6V4RqU8picmWZIY8JTAV22d7kVmi5VVTMlAdzzhSccpLYEgwSMOPYzvePwu3DK
bAJE+zZ2d7fQKVHGNm9fRxN7DyH1Fp16sqm5zTXFU3LGHpce3EBYsKuNbZOGf3L+
rLzYVlk7vnmn+4L51+APhe8fxe856wIfvDHKKXhE2nR8WxpNmhcE5zTpu2GFQZo8
HGy9sr3VOxPirhJv1Nv2bUrWWzb+dWXM6WQo33Fb8Zi0vf2azJ94wJMjekwRr5VG
H1MVurZieV4uZriTceQ1Opx4Hv6Q4JrAuEwfFVpDbH7iI8tTVPXsTU6G/yfO6naV
XdtAwsHXvX9vF1Na6Y7P4TGHZ1418gVmG3a6FxRuUoClcEP1VfWWA22bsWZQ5BKS
xkWTMP8dQFR/STNCnRsrJyLjoJ+rqjWV9pTG3IJndUAKThYgXv07Hl9gg1zR8Ath
YjbyfABfCBQiF4qdsREjjUWioMLL9RJWa8kAmo8N0pc0TLi0kD6WjeL63tP2tUvT
eDDrNKPww/6B074BNInyBMZbEtqkWHEQ8dMyEBIztbYdE9Z/Qiks8KPzpsw+HE6C
Wfk1FjdpXSBUDeJAtveZGMF/nAYomlOBmTmzvESz3eV0SJWsysQkjOwkI8uVAgIt
t57i54MznPXFj95Jnt0X86El52/d+8ccr0bZZd+uZKzonBqn5PaVe14LpJr1aaF8
nzmRntAPjnRRz3x4Z0zWJyPXve5t5nbuuLyR3vIQmO7FKuX8qWVdPfhZEbeasznw
Yqqr/TC32+MrA7KQ60sKI4Ge8fWbDsA5h+LdDAKwpYCqmeXlmN2qwMK6tjR1I4fi
0RLhHSYSJeLVnmyktpoJAvD4xFwJ95UOgPOeQ+y+t15B5V48A3jzf1lApjd/qaKS
59/bmCYOhsP0WkOzkjKjvdPAVX1FiTEwRc3ZMH3w22uZueoah0gs36mjPXWGwlFE
kjSgpp4iCDF0yEw/qPwVkCBMx3wfkaoE+uiIBVL6U0aGgRv3pIh+ntMaeBYRSDPZ
lYer4idYLaxf+PIu7rLwkm/IgTeAkr+gRKHbzz282NZwUycUUXaeCF1daMsBYgh9
YVtTvSzc46M3zpc9WekL2I09sk54pJpDH96R2w015LigTk49D+uSL4UlI/dyEr7E
DEFLZSXhD7JDCVoE36KnWzrnt5RuqqSkvpPTa3N7JBs0QwGdKUpn0H4HXuUABHtO
4hLj6EXPgdt57WqO9P0SL7Q0d9QgZ/TIZe6Bi65P/LnCgFHBWD7aU8nkBhaazqp8
HtSpLeAVYGVTANeRoADLMACHmV+pRK2cbWL1HSPZkihkpSguqTZ6tk9siI0adjg7
edK8SxjUd1FAsBxBVmgvGfYSJ6EhpD+WkqB0WVitfNiWE1fAbUT87i9WdSDPHau7
3b+sr383znxTirkXkbZ+gE/poqYaO6SAAr8JRYvkFCZG9Bms1pvA5DRVEVNH4xF3
akyoZEcPlO/P1rjCkq0bAs3e5PGAJ3rglnEzqyuJZEDUSYt1KFXp9vWLWXAWpc1/
5HmYUrJAfdDbeaBGpIpdtYPIl6x1FNhnecRwzkELyAga5eb+F3TMosJQ+Q85YOH2
2G5Gfr60zuMdaKMhmf1j9ENQrh36Ru/ZGKqr28I+4zERS2HsR/If5GmgJrFB/dPC
nSxNp7r0DQmnYd0vuzh1yc5/tniuE57Zo6vIf/klVtWzreAh/y9qDZJfDdUkFd4a
nI+2v55vU2SfazG6w5HHRRxoUXzVu1w8AOePlOpoXSfLChZoxjjlv4GhIjMPHbq+
pRugFAUx6p4egetKxSQ1DLG1FzFb/BTucvbxnxYaIzbWcoU+7/TWg60S51Y/9+Sz
GmwnCGZKKsecs2e6NkmS/NBmJySHCZTuhpwd5wWMCYUJYNpZ0frTQGXMLSHFA99+
HT1HCRQpRptf5PSlrmL69dnDrSPjLauCrLdSb8Bu629X9NRIRs9ImJ5oiW5fd43R
G9KMiX/aLGL1qVy56gBqU+AWDKF2ZjW6+/Z4mNixDVg9yBWbJf1msEN2zhVYAsKr
SvangI0zGJACJ2xudvCgJMytGNCZl2c+r1kURdP4wphr5Op+3Nn4b5rEHPlET41T
wJnG7vfj2ZLDWNcYT3q3K3co+EdX4Wc3+y/8fWdDs1ROa0po96guL9A+l75KirFe
UaIC4jisvsxM7o0bw7Vd9qC9qfDSgvfVTgnihxf33ZHjzxKo8JmKmjOkZViqOhvP
BYCssNOcYP3XrqtKQ8uAN5SJr7EoAr+Hb1NwhMmdZSR+9f1ogIZj6gQIcypYrY4N
IAdeAG/QAzcKdCOYOsjkfvYrp+c0Q9GNxkB5FATrk6ruat2jQbRVrdfKlLJd6Adr
hBWq18Nxy/5M+anwQGcodXpV3ZON3/Ymz1qRGIwaLI391SkIILoLbwDtcvD+hpC1
TD+TsNJJkO5ZgiQmBpXmbqFlJyObdvjYa/pdQs7kyzEpO0Ilp/Pg5KcamA6lAtg6
QtIHDwl8SrcjO7yEfcSgTD57xqEBNRDxHY/yV7lC0Dm3fvS/WLlAUxg84IXrXnwa
trRWR4uVEODYURntYoOm0aAnT2m92VEmUGzBEJtM6JKzdOBYQT3979RDUMllT7A9
+a/++w/vixRIsOJI58edhZ9dMUra4x/KZC9cM9IoKE+7gkmbn9G7d4HPkohVGzHi
+vOdqF3ZSAuqn8quEQEyTQNbr4dVZLuFTrA8/vWsD4Lh4vpiKapFJBTBeAsfDDJ/
3igWAn1EE0w75GM8pVxBCvVK6T/mA1k1kmlvCvMkN5JoUMbuGP7JlrbaDzD1VuGn
OdJLO15sHNYIYK2rOXfjp2iF6TqibCEb65gCLIw+q+mukNFI21brVWQXBWYUBpkS
AM86OgG6mcnKhHIQ2MKZEV4pO3cqn/xvi3GjuLCJnYrqBMzuHEXfa6LhZ+P1043u
aNr7uY4SGXacIb4fxEkEgOjESMP3c0zEM92dYi9lzrkwKeFVSxLrp7ULr1tCXUN2
/u8hjlh/qqY09ytC25JLMCb9npcTWpewzQqt1oqnmtbcxFykM0Px3yKqXjkvfRQI
5BIOTY0lI/jXcghvg+nnt6TO385uoLQiFf41G6rnXxO0rFwaVISzHySN2dGqJ4sZ
TBuxuv9LDa74AkPZtOvwFhdTLmHKEb/vWSCVSgT9lJJOrY2PoJqgW2MbvrAyv+6P
ZAATLuSrmetO1Q177bySq6UY8pG8iLpuDq3jV2FVmJNRmIrmUBDgnxzDuuxde/Dx
2B8VnPS9q25aw1gv4djOE3J/eLKgVApgZMAnhr+u7Tq8BaJy8hrUIklW7irTILc1
mDVERG/FTRgQK4YFL2gRlTM9+th9rKXloLljVQDa7LaRGf5ngWTSSfViIrCHvBp8
dg17+5poclLjA6EeN0yHKGoj58xKXONB4nFllqq5V94CrFa3VdL8BOklUFlO/VVk
hR5dyvFXqlQO6G0KhVCj0dyMgujQhaEn/zZxticNOfQSboH1zXOh8W5jDH/VDhmx
lqw3MkNi6GF1RE4lPm8kZtC0CjYt56NbqiXi4ycD20y+RFtPg6BoY0r83JgHwTFv
z9COIZa54hYW9S/gboaTanQXyt/trDgJVx9+5I199K9yWXoEHDovtBXCXsJBok3N
jVX+G1c2sadOmkO0x3yTcXO3w03luSUArn8kex08aTNnjDEUGBfNXEQP1pzTN4Tq
Rry7BC6mvFNV7PUsD4UfBT5P6tUj5MNjoT5VzyCqPFwsaLy/2C3H7lAN/mYdY2V5
cVrcXi6v4njGEZq1AJM0CoDZ2vf59kWjiwBOogas/XYBAnhC5v8S0sWHfDHEJf8H
HDubWBAF6hnkyio4qRPaQNooVJE6TC1KQNqRG+cqN4nmSMXlDjSsU3zQG84C6smZ
GL7WZ7laLsKIsWXF4NyLqqrxRAC5gSLxTmNte85yhIuiFwYSGQZ9VHZ/p0eGnDUg
4X/U9CabVXgMWSdkoOxaD/eWv7Wo982+HTou+LnnoxWfPqZ+/CMd5MBIiwcJDXxs
r3NhB2JsOaPtKb8pNNEDvxI6cy3YHasNPEkPSh2mSyUJxek6grwHBmLSMDV70k6Y
lOe8oUubU3EN5SzEs213nUzxrUhghZys4UKuoU43XF+SbE9owqGaVZaAc4VT6Hl2
soTyMAYYzAK19r4yXhhDQA4jJsESCupP7YxEryDceK5qaW2fM/bBtbLlgPZ+KJZr
BSgwzibSi8XZgSf17/kJDZy+9qr00YjltLYsVWFQWJqMThJc4qYpihvm3D1fJ0Xa
ENZfAh+/QaOZV1cskjSTUpHyXZB7b92LmVW39vWp8YAvwNsGW8xwDi+s2hfWMcLv
fmd97GavmjpBjXCXCTEqS3r+v/hwzud39CGKnwUs6wEU0BESfDUTLYGOig9huS3M
TrIziTlROObDtpBFZaaaCknDMR/fxWwniXYkjrPfTkGauAxezMrcEFehRXD+lcl2
RYfsRnzVM+FMkOSmexutnRsUWchA2v9SePIOe3WnLzXSeZ1ujfQC/0RgF50/TX50
4gbWk+zgT12T/rophhXcMYyEa1N6ee0WOTWPHYf5m7wMvpTZO6L3G9cJ1H0xcmq4
MI6xigDaHQ2K/D80IodxJkpG5VdqsOmV7iifxIof7J2ROvMz7A9LvKhJvBZe6WeR
gZEETZ3jWdEvh+OCoK9N9cx3UN5f1t8ByXosxwXzzA1p7YYXAjtsnd+wp3TX6Ypp
dIBxSSMJg7PvU52/ZpUXHz49tSUHsTIMkgDS+LzqfQ+GR6Ho8XhFJcZJmF115fsc
kRUG7m2qI8pf8gy6Grj/OfhlAX2CQU29bqSGGURnlDm3q9v9lhTAMFDUQ0owrwEr
dF1OX+E8iNnpF+d8K5W9F860b1UUe9V7ww/Qkqqmz+AHWXl5cjU2KnJf4Xd6S6xf
cTZUhCbGB1y9U7DPlbyPi20LRfiouJG34ylvLuJkPkQLvkSrohURG0K1R91KgxZG
Op+Ct+UgVimhjvJB/D89TBFo6J0cHsITl06O+NaDNCOWrwFnIa+TohoC24ughE/1
/cMaMkv8WwjZh34jNvX4gQXPuQdmDKDDJJ/t7koacfkggfwmddIkhfYGJv2IXYSN
+MOdfIGTYeGCxKlW01mRJsGdrIrm0er19VRLYwgQ3WXagcjaxpI+8mDBLfyhQAOJ
e75mnAtL8uLKMlseKx0mw+j2n9vEVfeuKQesO5Ek6cof6xsrQjQdA6t4mEPAQUE+
CylAtIlD7Udb5LKIn1oeUdSP5R+vWED+UvHcznYFKb0z8RVakB9F6Ey2GoV9J7Ew
uJHd9Y5bWeFTlX0r42Zkj1QZUhxZyS9dXgVr5xoAw19y9HKuwdL18qNccZb8z3MO
E4F3FCo/l8q+NCrBfnlq0F2X05NcJ3BhCuMIcHrHGbfjjEIPk/zkwiPglhivuM6B
tTTN3HjKYzkmm9YUbxaeGg0rQPrun5zr3J4pp/gBpjSE4jFdljGHtjf7XEi9ON/Z
OUrzw/T5yobE0CXl5op/NfMaHq0VMRr3BdXA6acKttSZrC3wdTTNbd5YglDxd90R
t8nQ0hF3cSsXg5P+2yD1t3lrigU26fAI2dA8Kw5zVVPCwNPR5td2/he0CTHAKQFy
vcj1IZyMJTlp2BCPa69hdKn5SQl3Bb5fG78HlEr0+90e+36hiAR5xEMlGI5LJRuU
I1eS5YPMdo+BTdkIFEixfLU1Pn4rm7JRZ/Ux4BW5K7yuJuCKocg2Q16NUZlG9co+
qVAsnHKD/HqBKq1KvOZmmrk6yyKgl2YsiIIF69Y1M/aPc/vPSw2BV6vrr1DJMg06
/l1zChTBEEWDo9INRcyOKBUYEmPf3OVMrJpd9x/qog4oFGsoy+taOueL5cQ02wrr
SINS55tAFBKU6+hhpbFRyrwGd7wOKN7NZM2H6JQZw4OpfkJWw8EcfXkZkqHt9uBa
TbE+8ZxW9vA5lqj2Iu3GS+0srEH+R8LyvHM8FqDVub9N2/UOJAb+IpaIXzB4oJIh
n2EhLB4TbBxx8SgFw8HNg6TLwNzDmPrDYvx7Y7tN2f4HDiJvTn7rS1TmHshdfOnG
rkMUH2BxL4Z7yMXpPCgICM1nVOkbrmTh0n9BMuqsivwyWZMXmFT/nb5/9dIvT9HP
gSBY9qT00Qhd2vTO37Lz7xlaJKjfAt77HMxQFHaGqLoJL9rhFYFGG39L1F8lCAud
9Ja6Vi4tbFHOmGLPO4Nc+Pc/6Hd7KPnm2ZnibiOgFnUqXHGPpB70PbKPToVtXulw
HVESza54tscJ3vU9PXsajFt90NcO+R0WwmMHVlxipNUMpNuUWz590OVDI465ZgIW
EMKWrYrQ4pRHLLUXd6jhBikO6/VBUog9EJrIFlLqPlk+n6YuURAYy0mOktjo2UgV
lKvyBKZgzxhT9mN2ymA0XbzMRY9zKUeDA7zRuIEPNjixsR6NcifT36kzUaikW4Dz
xVuTQNkBtFiim7rBfv7uMf4de6jDN+xcLBvQxFnj88CaYYYvKj/4SCFGxF297Chk
WpLN7M854ICdFsIrXBKDuwcOeGqtcbExOfFnCx0vpZz+rfkEGtO+trOPkV+9Brb6
BnzZ1g9JymjPyVov/vcyg+E0TloT4K/7Lv5BPquUbUrRHtfSeGyqUHibmxVTeWdL
fW8q4/sDc1WZezx4PWrqIWbALMAyBO+MfXxr9yrjcr3C7lKKmnwzgcOVsaJKT3D1
C56RRO9O2JNZliTcZ8NT+vLR3U4j2Wl6c+GiSOkXnLgZrFw/dpN1i5qD8k8kYwiG
5jw5iRlh24ssYSq2fIMiqoWp9oWEFN6rNjh/JvApRskqTpHsgYwfvU2ycdnw5Mwk
6ZdiDRaWazScsMRv33PCrh81obSZ3BuCjFo5eyU81wCgvxhLTddvSLkksycpWdJa
m89Df3AnSfNUHs+1KaBxN1cDGgiPCdC+Urf20G7Lt1QRO2B1nEo2kTr4pQhgFtZT
uEDd25k5MX9Dp5BdM5FjCBkqczIeGv1XTRwKFOAs+QfUrjGLX9KBDdd2IoEJVQq2
CbxaU7pmwY/Ax+BEiMbLSKz3mAJz9+dtLbI4DXu+S3aREWzYVG6+6MI56HWXH8Tg
adfwPkqDeKw7/x5IPS1lm0tXCjTtiJGcR/RBPGUjZJK59uGYtI0uj8H5CGw0sx6F
4oEW29/PLYjmBlLaRfI/6WqmpUAz/CQawbJsnEPtYIpoIrwZ/aWZMpn19Lxa3+1K
AqVAwlUu47q/iXgXP+BAbY4DtUHOY18HtkCr8c4erzKsHah+VBGSPITnc2VPQhz4
x6Kz5ykTJroS8d/dpxa3PdSl/19+GqpN8/JSI+9zWL7kklUmrVERwYAKswc8/mJ8
DL66CBudlYl5xUXFujn/XnsjVc5UEulnrDj+HjTTz5wyhjOL4l61Ps2J34dt0lFk
8w6ltrO7+iho5e5uXHWb7JQzf7Vt8OCaWbViCfbIE7n7MKlrQtJpzFuNgnZkv2wf
uuufJgaMwjvEn9/HWhm+bekEmAyfJtvzbYUp8mqk/NZeZxImF+VZBWi/SPSNAeiX
b/wGJjYJh+U9tQOrk3y4sA1xkwToZtpT6WA+fVXs36zROEIbHEOl9jNCzykr0EKX
GwCS/B+vsuG5X3SkJ1ys8p8HsUAGD4jF87qAybDHPUXI81MWZ6cao5GNjMAhzjze
KKasa+EEJsfQ4ShXRC8tcjeGcS+tdmu6Nx+F+a6ARkaKxqJM7xdp+L3Lqo8zOhYD
Fy5m41elailunVo62jZp6mXiNoBrI9bDDgs/XyZ0ikWMlhlNmw6AU550I/4HPaCU
IxnokvGZD0xovggxle1y4Uf7WCRCw5xSVnO9+dlSff8kXcblnyj7NksnbKCdYY9G
QB+pQCcLsdXk+g11uaJDxoRpSMU7yjH9uTD4RaYrmv+bLL4wI7om+Npfsukqr1Zx
jsMWp9n9/sPKXR8gVEvT309Y+III7gNWnzsntf77qZXEImC8RSSgG+Wdw2XcAdoe
EsPaeMpYdXgAhMQXg/9vDCCVEIWAA8XWUx7FY6Mub34d9HX61ELI1qjK81IMfbaR
Aenp3yW01uBDbqGuXp4/Og3JSfErDIFLLFAzLA80K8pzErZYH1YSghlfL0zxAC1X
YyAJ7IpovPycPLSXGGuLGiwFCCi+9/7i+0020JpHEQWuI7GFH6rQI4k+zryPJps0
YUfPDgf/upqL1nUBTBJ2PR7UN/p6BdYq0oJOB7/1cIiOvcdfQ0bpZUZE5xoCMKQC
jr1u7TkJ1KkaanJ9Zyw6opYUB3z7Yq6/sfdJtGJumB/KmKqFxO250DjE/f3b4Dnu
ZyhM9wYYsmP2YJL9J8eaSMZBdjQnTDLReTsIOggdfKktyOd5KesQx6GEEjwFCJGG
V2MwECALAV5hE6DYVWKVu5S30gwv+7+GI5XN/5f0JN9p9BW9KPLAUpTm3F7koheX
KwdH3N/ri/sKM026CYejfN9/BQ7HbMy6PtcgkFWMqDhrDNpULVl2RX0cQ0qd60yQ
lUAKLomqFNEcM3OCk1KrRWi6c+S0dK0JdehBiC2DeJp/QOlS6a/u1DAIYrnkqa8t
btx/H7kNHtKy75GnzYaxjPiLyS5l3AGiNLjVra+vAoa/dvXeqjrECTdMVIMrC0Ri
sGvu9QXZ6wuv4aMf8SeKW2JWRLWgtS1QDqzQtHbePBe6V6ED4S6kA4D9mR5TZne+
zxK1qHL3CKP+pM/JmiVB4QIGPQ8O+J+sDfdnbAY53dyZ5ClTGW8qtQpZGbscZ6bt
BWg0vAPiMdfBWVUJSXO3n7uF486Rt8gHeZTjCDIWsjRXlFqTREeVFXsfcLZKh/zX
iB1Lc4+QNWC/UMQYs/AQJ2gCVivVJRCg+Z3VW/q6ffX8qZl9EfMVpNRsmhA6ttBk
or2wSSqZJDxnBq8a9t3fC3Bbmf9N/zOcV+HfEH2dk5s2fXewKISA+UjTOW8LgKEh
sD2d894rmPqmm6I9m1sZGU0yz9hPIQmw1kpMALqdfnBKt4kX0Ze4/SCI55Iy+j+c
H5lQhkbcW58k8mFdkU2t8cWDnVWJuhws6GRqmmUdNSsdC4Fe9m6kVQPj8+5yYAtf
H3vJ3ils03S0RQpEGWWXBx87Gln54Zt2E9SZBXBrP9VRz0eXUCuWF/+F6WvJlHlD
Q7RZLvKSB7eGB/Xvtw4ghgHeBSevtaq55MYrJFQ+o1RdWxVg+zBhzKvg2grqowLq
d6LAutoC3I44LY6AuiYqYMY0OwZfq7H0AhNX/2WWe0rhO4/OHT1EyIj9/S2ZUudo
zP/lu5UJcjMPOOkFt6QMV2BYlgm7Yx+k0VX7RmaY2DAU4OHuoJHtrWkVU7zbTtl1
yK3XnPlmrvzzKF3CQiugeI7QrSSZx292polMx8ZM57dLzPuc8H/sV3QKVoQJc7Zf
zY0OUkin6y6Ywb0FfLCmIO2VnPqpTyp7WAHDXKhB9+RRkpheHB42bBgI/KRY2wpz
9dj7IwwPcLLH2jO1juvnVIv23ctoQn6dnxx/Z7MlGqE40de0IiW+wXF1pUVE3GNO
OANI9J8VJRByg0SgpaZ01YT/9kvHoiuxBruIvFIHcoRxFBo9V9Ub8IL7SjjqsV7v
H9lRTfQns6XSamLV6znoujwn9KaFBNQKYKr6ajtvuzIwMwGk2n/uhzcQjkdJ3t6H
azevUNjinvDIO/8VaE4eUeQbU7H5fCZR4K9vIQPPFUgcASoBjQjTRS+1DO8TqaVs
jbChnnuLqKYyFu7/U9l2JgSURZ7D6p/1GjqFw1zMaiu09eJfCvBdLEQhtagruKnc
YNLgOmlR/1ZdPPCY4J1tkUDjnqBcoygoARFvsPk1cw827qDlI7tg3VSFSw0UwFXI
BlBVp7j8B3TyhwVQJM/SfxcdXzbNkwuYlhzUnLUGPwVnJbaOWHjZVgMzmobKVTTk
9R3PVs4S+wcolRbRggtkpSzgFuliCj/DdRDANi66W8jKVxG6vmZIyMe9njNWHUWE
i0WdNCBIblFyOpJprr7Ii1IlcsIK0tqvVlvxhbzomkph0t+3MGGN0vuGf5natV/W
BENB3utb302R4xV/P+WI92dvWgTozHVFeM5M0F3YCUXEcr08/zlWNwrBmR58Z/LB
1Y3tlW6Q+fyF33491L5glks8m5xSq9tDzD0FisPUUq3ZPJF/fRjT6HYOzs8Lj2P4
WwjW8xTH+L54AsCPWcE6bvLtvpU8gXBMcGcD4KDZHfFm7wbFXGydyp8hLAtrgIGZ
63OqziqOMrDnQ/aB7WMTN5uXxKuj0TlorjQ0/IFVGrEKfot+sU1GgJ+1D+MJs01q
q/Yv3strw1xTyktf4wERYyNt702+7O4c1i6KZxvtOX/n2FqBrrxK0A0zeENwaEQk
hA9knC3B1rT/jOJQ+AoW3Vv5tPHRi7rm32QjulSn3Knx+KjpMv2TLQx8+o5xZ3ov
AD241PguYTcHtP6ws6KZGb4hZbWLgZwzb26WLkRX9uv6aj1I7e03h+TfKnzv42mK
oY4hOlhh5XPuVb3Mrgg7A/SzOiTv6adGJbzXpLb2e251tkP60EjZv/v/Bzqo0NQQ
E7yLOr/rtoRjqfzZvRM8tUNfbKxtX22so/WsWvglPrMcaMRsuVD5BVFomjmuHsFT
Ht8EJw+kClKRn8GuCyqOCbjzRPEgezTvM3DgSCxEspZvQ83EA/XJ5YbuwjE0WWow
cGOzjA5YCfWgGxEZI9X8kGos5QyBHFUA5iZPg/dbo69v1+F4FoqNI7Cm48denb6S
tuwmHW/2noO5RBwgqQaWdwONsZQiDj8/Y5ftHoeNuTNO3tuekRxhrk41UiX7/Z/9
2ec9yUnImSnXQL8wRBl1euFm+NN6Yh7H2aXD9BVfMsI/JoiDTkpTRDVsG1IMXDoD
i1gURlE63bnWP/MCC0rnRBZJSh1LVkDPgZgcPAgZWeKP7wCHYNENv+CH/W8G1/q+
I6qvdBtVgWOsys5BRGd39oB5g8bufQZPyS3fEmndTU7LZs6Vz1/6PDaJVWbNOHkl
OsPq7eZkmnZtdTr+iD8tGZPYABioJwtyQOi8nm+pwSoeECiHu8GB9a2E+PkiGl5B
XPySmVHg5zy+6OWjpU2vqFBs1GXGwMRNVzqNLzQfDZ+ABCPRJxXUaN0H4Q4T2l+q
ZlDDPOyawHgippYaCNRMiIIIDDBdDi8ApEgW80zQYEXTKWpcXqaWTtsqHuV7NPY9
juJPJ6m4pmPsXn9Xczwi/Y8SxHMAIqOgc02jFNGnw2AglWhJ9iRRXUJxHNtXwaWy
H0kfhtjNqwy0dZaVebEK7OddLaoGDy2dqavRZWvegqcRdj+PU2jpYSWpcryH7hlW
4oB1N3YgYz+hKwBVrKKrNdaCb1mFCnTEL5uoHD1szOrdxqnnvSRJhff8lD9qqo6S
N+jL2S8yOmK8eZSta3cpxY/cZyQrHCLzgQYCdmNdbXdguuP2ZxWpluoEDo962TGv
gx8L/GR5vwGd3ICJWY3DrnjnaukNNtNMgeee4seNstdwAU7OhvDtpwrmlh/KFX9Z
1Aey4hzjOmDCdkAoqlwHx4+K1pXE//lo1q1Pwvyr8JR0h3cE972kI+Hz965ZiXQA
ztUvlQR28p8RZxEgpIfOA9og5Md0+JGQN9ylPOzj3NOLE2Vf4y5JsdGAQkX317aX
2RUBDOlDCvN/SBEfegux20IoBmtL4I1YT1+6TfJn26sXE3CY5d6uRKqmGVETyjEY
3nOUyhJeD7kqabo4EjhUrlOySM3X6n597gA14trw2XsDOP38Bik3lqZel7aQTdm1
fhNgdBWtejqBsTf7Bv1W3rGlmCdtRkdi9sKkSsfJb+8aUAxSoI8pcazcVSj/R3Zm
bZjO3nC45qNcSvCCbttdWa5EEMU7OIVHUqLbyHWczJ8OGiE2Pl3kYDLmv5l1FLjb
hgVYLEoaJ2Z7IWkJPBwdek+DKAB/gf26vsKRQrjh2y1mo05kpdHO1hLV8FsnTNlX
lBViPdtto8aD1ywrdLCfEoG6fXU+CPjjWJJ0PrKx4qFJFvKCBdmywL6H0AGvp6jT
OOJhHPu/X6fcdlBCAcavaDC4TC8Acs3rVUj4mjoIcNvX1g3Iaj3SLeu0QlhTJFd9
FO2ZzMVKuUL11/UszEZ6WztoX9mNyNywG7zPLJ1JtGqRgklYSbyAenQcJaFrrUV5
v66XmnlAlQ9R+t92Nfs5IiyQVLjVsPiR8ithpDDVn33+dIxetre9wOR9cQOsQaqi
apaQITLRZuhB5R2rE+COPn0/U3qCZYXYRGVhIcM+vr5H/C95vx16wwoe/5dSBe/1
lqghOGRUaNvuhybLtgBKu9e6IQMbFS2Cyra8R+3uNMGU5EQJ/qF8PdmxWjuQOIpf
Nea/ld89Jdn1orK03fj5ypUpCINMSbXEqDpr45WtJ4cZ9YA7ndraBqxEyTrC3lQ4
R+S1l3NsqjCNOHUPwjCWLw+0tHOr7PxbazZ7c2BAHx8UuOq7aDt5Le6rZi4xfAgZ
bJ99jaDX6qJHoA78OWusUvWwLHfpGh3oPGSxlmUW2Vwh5KKoPqGuc92mmCfVhoy/
3IcDjUnH34qh+Y5WHBFsy7p89eSL5uGPpeKU7WwIfMif6+1uvDty/gWUr+6yrpkd
aL1SA9FyQbTsOpXVsVWwGUtA46bcHqs17rWEkHZJxVPt3veZj4EON+cnWn7L1bba
+0fYndodrnCkRtyvip65YUXVTwSMaT/uwQpOb+NPzEllZekRBQNNhjoWzLSqs+8q
v012kglmbDkPsccQinEeSmtmaSPb6S2TpHdLJhtBI8W+uRb06Em6/nBmkiY94Gai
O7JYP+DWOH+YEMpOD5WqpbqMqYTi1AikTR/m4vf6Lnu70HDDpzxG3EQBqAur+egp
4Obyc3dQltr+u6GZWbRUyYC7E2QjxT5eeTpeFE/sfDARnS+GFplvse3F7twH3riJ
aBxUkweYE4X/+XxT9t6czV+g2JwAF9fD/lGRWUbJu0ab4uOA60Qqz7S/JdIragHw
9nvtgUer6BPe+V+vNMOao9er69KN4pNFgJDR1PuehNz36BDQToT1lMxbRLd6vTyY
uKU/TuZTHdyLfGBg9Rwjh4KhLhN1YwpBe44DgnjW52rKgwcyOcBFCMZ8sclKhbPG
YBnkOrF/zKo06A0KUlCf6BnnkvExIfU0YjER7wnxVM/6HEq11ZYBYAbESK+TAq/q
5xz+K44DlgyEVNZ4FivrcChv501COlbnRze3DRTborB8he7W2Haj1TJuAZZY3Lg3
KA/8sqsLOApkVYz+rLicuGrOIsJtqhJsyHyfOH0xCfkJ614jKkOu42tzBAsG1knY
9f7I0iyIdSwKSucLRuvr+jxUMOr+UsqKzNnq5oQFtFn9xmFLqijqQ9Ur/56Ix279
o3d2SKQODNHF3bHb0h/brn1m1FgOoS61wo0ZcQGTvh6ipeKRxnHiCpcJ82nUwSJT
KaGc8CG4NROh6FxI9R/tkaxSnk5kLMomfJVHcWrJT4ZHUhsWORdVcjbLH1rV5uGt
WONQrAWDz1gAPmJYrpkkWa24M646+2OUiEyeGmjE6Pb2Y8p269LjAHmrqE9e99HQ
qRrFjikIhWboLDWpV3WRO9cmNsavnPX2tAIdOM/C1d2kQRnsQSUTL2h6GR5lbt8I
gWY7WFJpO9drESvcsJNZFAkdGN+3SN/W0ETlFGe9gcjlubdoEubjVX6cJUvgHLnx
NEsJ4TEeJDvq6ZlcRBO3+nYkzgkGQSaUuZx6PjrvDUksxVfkLAUQxfs1Fzx3+7ow
6vLk8XVqTKlawP8s45T/p2+t1eDa90q6J/rrUWWvzDGnFXI7hKi8FwBm9tDNMO1I
OVnys4afrforC+xPsULZeS2G0gIgNmyXzLUSP/tzTQt7TRm6Ylj07pM8NuPioEqD
V81h3CrKt3FH4V/x8Yxe/TBbvzUR3H5TKJeu6+V+/DsLyMR8NyhpGoFfEOEH7Qib
j4RPMaAVjaZVtob0mJmXe6uB/cfJlmEdb2wh/1jAnqGYen6EqywyYCIShJIUjwzl
WXtncK4+DnJMzC1Lcxpx1dt0WtECnYDsDEajEV8Qslba2SbJrRHddYog19jmoq7I
8gcYW2ibI88x745nGIZbH/WLCFHqjUXMuSTBQDInOZs24S0QO058ooWyaAN0gXu9
IrshVDrtpKG9p3HLrtFL/c7pLEqpi/fAbV5jkb5pFutLjGRIeR6gEEHapCpTMUEg
gvBelvI2CIAsVI/rCQKKiwQ6VvisTJBCjqv3X9JIGc2sMM2viMJXQGlx3X4wi9Qu
ILYGwZMWZ9CVF3bXikvzD+0yEK0sm0eFSNVCmNzPY2VppbtB0vLpHivDdDrkgH1N
QstSam+rcVwtSfcL8nB+ZJTPP5FLL387pTvxQMchvB+kBHuujhharY1pNVNTMFGV
liGP0Le52/Q9bFu4JKQYNtnths4TeDH9d5HwMMW992h8Pho9yYyB6INz6oV8YT10
haXJr4yWhBqTNHw820mQQmRqI0EFoy77pk2pqW+DApVIRoNKB4PiNV1lsar6rtmj
Ok7ZcvJtDxWDe5LdeYJt7MYCPYmHhbBG09Q/ZbJ898onM0QQ82lA3zdcd5+qaLPE
BuAb6Img/5VdRTo+IoX/eeiF21+ikKj5eCBmr4cpji5YWo4nNIpht8BKb7pBtzjv
GDFS3q+oPajnSu5PUdC+a8nUKjsLRKLRRU7njzZIqUGXgLK/fwqX7KNYDsXpN2bf
Q+LlJmqZ8836cEoA55qM9Wik/wmMvG5fMskR3lzZpUvLaK4KU5t+kYK7zdLnB3+L
shVN3p3EZWi657cv3WpNcjdvQoKRCvb47D37COANago3HwLnF7iPevDpbzU/+oxK
9tLRdP8jaM/4zNf83D0FSRFI/YrqFFvSXdYNjKN+HPdQ/Fw8fbkw58oObuACepIv
K5n7j/6w/s+Lciwt4l5RKrsrbyyCakfjvBRJejvv60gXimbwaDzfrh5za8cRRZ4N
85hn3dNjC575SC4BAQvK+GlljGtOYwtkMphV+5WuibAjVS6VjnnoMFYk907Wwc73
tEPdbtCWzb4xRE9bWiN0yBfE35OHCEY+7s3Oa8LNJ+6t3NpZowLcXnxaiF32Towi
NFHECYJ8msihpBj43gRLSANN8DhZ06tZ7O0k5iu6qBdjJBv9+G1gYk+vTGPR/yl5
uTiI9GZZkpn4b6zF5AQSi1x8NXAGqV3tEAK4Su8J4u5rHvUMQtGP0f9EMZ2iNRmR
Fo/zVu9Wkzzq7sog/D9rqqUkPqp122VIthcaMJDiHhaT5M7cSUdHXNkn77grEznx
XSYjGsBVFHUMB7Pc7Z1YZJ73SNQTEgTtovvZ85aZmuv/MFFcqLqFzn0qEDoH9Nph
oZ9cZQUqUu8Ok0Bbfj/F7FYkvP32o5agrh7PTFd33kMvkYkzWJN1JVEMgkM7ZggZ
4qUvYN+6VGQFw3Kw9YdQWug+nWzCkvd1Ndenp00FPgbWVssJ2Z4zIHThrvxC2CQh
/UD7uJL0AcWAJwwLAkEX2yN3xaGH1t4A4eDpBCXA5VSnPwbrsEm/+FCJFYIsuApi
iKvZz6+Ki6nzsFLRD9q5sqRlVZ9vc3Rt6gWljVIcfFAACFBL7Uuvnhthg8OxifMb
Zc1hv24sCHBpXz2NfYlBHpiuONlwkpl4sMf497203zIBYNzTkCvAZSlRseaHeNeG
VkteWyAvnbYorjREGfhMZNnhb+LtLORgIyMF15KE75rsbngjMQkf9FHCcK85y102
UdFn40sCfd6A9c+Pzgh+Yv3f7wZCiNt5+xA7avD+bfMaWLQZ3F+Ax80N5ehsriiP
hk2OYqLqUlpjrFTuLD8Ossm6Mv7RTcU9iUn1aYPS/TGC5lbzWYHUIPNGN0QeC/zx
2BtHzo8GF6eDbX2kRxbJi99EdylouyUZH88n8xugLiXoJXLD16IgqPgNpaZryxaS
gZOjSZUpkCrGlCIChfe1k39pS904cMgqaEHWjPum96JsXg3+yHjP4ZeQSBVPdkBE
bn4IlUKtAO7tGTwGlMDfD6fpmksW4Nqw42h+lbHYziL38nyHv0zdwksPfEmcybZw
cc5O2waUBcm444MrbrQGSEyxTv1Qk+gMCatte/cONj9aLTA9YcdD7jrkoV2+JBD/
sn0XYnTvEcCmDOzXSwLJO7Ikcq2YhttY+DWfsXmzxCfnHQk3kw6DdW2/NAk5fA+0
aYRWXjhjlhhXHZnVwIFOZJLRvRqZQZvrQdNJljlm4HdFefXM+bA/ZPQKpkxLutKF
h0iMqTWl3A7/qI8MaJf8c/Ted/BWYcts2Wfj58QDm0oNtdETfxQvOL1TGmo7f0dJ
GplqKeG1jEIWHuOqg3lv4yPZXwH5QR0pt9CVoJuxbskEI8uAgxK5qVP1ux++SPQ0
dlquZoSPEc4oWYO2HMyQLEWQ+av/xM/eyrw9VlPMDTyoHydOYptfRvVXa28qVhf7
cFb7A5LD8hJU+nGjDfSgvUmPlAiiym3KSrTXnbKCvLliirpiI4LDL1K+tqlREDQy
xCf+TgzluxRCtT1crrtQTsZY5Xl9WLH2z7hrghNmbbmTwPNBYbRrrxJjwiNgHHPi
eHyY7vhH3XMIL/dJ9A/jm2GxmTv/h9U35Q+wuxONagWLWQ/k2ozq4fy3YgoJA7cn
oUNz2FBkc25dJOqgxHA1N1kK5euLV1S0AQuJ1KwD/U8Ety4PQUWGJEvCcSsKg634
VrWhRfzLHJ3rqdXVNSSXm8ZIJR0TmmuRcQ3NHcTrNBNG+eYQPhwQfi5/Zf8RMHCQ
3jAhQrgxEMwrllFBX7MwiUu7IBqH/F4bIbAqcle1UAzvU6D0fLuFwq2INljDZH5B
MhlQONMo288P1d8JIw8oPN/hPdHSGeHPrmgTr8jUH5A7SVDXptJjURulwaKCEMKc
AJgnHFdU/oOA2/mlLBOOM1tVvq59HFHy3KMYuO6qMSY1WAwIhVFeqIFWkXRZqPQi
62WZvYePB1S3cFObegFMMZ1cs3R+5EQS9LldVeOh6K7mD7XVFscJE01B8Sz08tiU
svRZu1AzvUmfMwBbr+LObahSsFVLgR4MbuCTLOOv8VXG2UV7QWIvZcixgtq9hIfR
f52vtL8uPkfe7J9OEEfkz31PLBXj64pryNGhEJZmuxZ5m8Sy0PTaSDjz/GeIwadG
xp+8pig4D+rlAku6HFmvvhCKoBAMLnXiocQrdGJ9d57wMo67BJwSmPPV/cv0cDpT
xjgM1+ZcuhYuS408sJeGNx4d3/YoQpSU/PFEGCjFiAiYMs4axEn+tpl89TDzIzKM
lTk+vQy2I5f7T5z84j1HyP6nVc7+TWXZXgwNFhCOyl5lXnmEDNPWFEuZnToQ2Rhj
ddF41giQaq2vieWzmayobnvfC/51GUtWAtlEJi1LghOlc+CAluetKgNfIDibKvn1
H2Ok6m+LTD+jmumfLnzZxnBE2EQc8Moi9SS45dnIWGTSp5aT5PqTWP/noW6j8E9y
DK7XB2FCMGOa+KaY6HrsP+CYSEhu0oIZMKQauCHVnzXxt40e6s9UnsAa4DTEFIj1
WcdAiHUkTspCSSG6nyyB+w+QdtAHtkIu5SxjzFVeQFb3O+LiTMmzTiG8iYuBW107
RoT+p4z7SbYqDvycUWJQdQVjcvhemT3Et3oDmz5wVYCVQjEwgbG7L1yVd9b0I/It
bGlJWYe13fvGPJzRohlCRTSe3+JxjQRRb513HM5qYzNh+cDbmUOFZr3oJgSyYvu9
0PBrcZXceT7aPOkeDyvttG8ZmuIRPgy2BXsslwNa/qcaLENhIy8qyGaO79LhaHlJ
ze1jLFWM3h+tP+Ytb1hwBqxGrp29+Kz+CP94Zu58ZCf0UbXJ2UmGfddVh9zHd0zB
dM9ASmFUAXQs+PJ3AxniZP9KXNQsbPwjMJnzbnY9rMFkxIimaTjEnccpZHb2YjKT
J90uXeEKSDipkRTaLhiDZO/jEzt9JD6uQsrTY+QpMjr+leL3DVCaE/bi1wVrf0CZ
WSHd7ZmlQJpUUg/vYbUNftGswllQMFq89DBTPXylK/x0Cpxm38VyYZJHRrHAOB60
m4DVw2VL9pUGW0ftPJoaEgePXN/JtEe4KTFDMVSci7XLLpHvjUjLmbXKQuIrXc9J
wEBugfinB8547rTAMmefWkhO74vO+Q1gzNF/tu965aVDltjmDs0D37+4zFaymYIh
fJk/+xeVN06BIOyXloqoVWEDhDkJjQPcV0ozhkxurB8bafvg+kC0DBR+5G7N619Z
UUetOxsvzdsvWJzcILm5t8qKv+zrRLNco7HzCOk9MbjtozvAdo6DEo7FIXlzZV8j
3l9m79h1degAmnNWUC65UaX7/dfOegMqp8Dqh86dvk65AVrz1ANJ5Clp5GeUIJOx
8iuK8BjxzzOPZb9dBpJUi4jAFE5UOQdSHbJG2H54B9L4+QzKB0jGJO1g+ucMi1p9
ncPF2aUpCw4+cynConNzJ1S/J7ruswIOIjEhHCOxXFNkaXPOCNYaz3TGDIUGqkTS
w4OyaANuLOaWRoYSR2yFjJqQuhrW8Gh9HKG293Ct3WFHeN0t2FovgX9q9ms6BWab
45wk5Fgzp7/zKU5UPlar+9MxCgV7E/MYd/QkVJ350Qkx9GTYqBcYuR7iQp/jPliK
BchRaMYUB9tfNQxLg5lanFluNtKAGYIktnDgVbUiObODGMrkLWmyI4nVHeF6KD2z
602n2fPftqxDzGaSJ+R7MnfrWMTUAQujUax3O29jyfSBVqZogGcUCPV80ekKdE7q
BL+/9PzO1l/H5jKYtgmbJQUJNvphuIBiBNuBe2mkjfVmTCfDLrSUFTZll3EhWD3S
nEXNtVWnPqUvaio0jI66lL07UA4Mijndf17KCFKaqk4WPgYPcwNbpgp6YvN6p1FA
SxO2OXb6xhGVcvYM+aXJW5XLRomgVziyxRJEApGgQdRyW2RyZnXYGaIeFRVow0rM
eMhqGnwRyfR/PCciRQDoW+5Sh8KpBR+vvKgYbxdthLvZbnfb8q4qwr6f8sv3c/g4
8UMO6Eyf526JZPVc84N3xZq4RdqK7KHhD4ETMoTs6BgPFFg8H27t01mob/Xme3iB
3JSzsKIr4+OjTas7grBWTmvqKUjxNsZko+z2N6eAcnU2tBJD3FZ8+dHabBQzNK/j
grpoOeu9rLGqO3pbHaoQRZQmL20tgOxFMwlclvyXgxntnEpFHL4G1wlUxCxJv/OP
KtO7dIu1BQaYpKt2tRG8w8KcFXD3KNUgO6/Hk9Sp5OVTrrs53YkLIoFzofaTj4in
AqUK9o+zNR442/mI8fuCcYpBV2Fy59DjTLP0uKOGkH6bhLHCqHfeaMcq/fPjPtyA
YU5WSJWz+W+EGUa+zyXodZXe9XOvET/0oqy77LtYGHhogmIN7wM7gtyso+r6PDgT
KX3XtcqFItx5SkVzl8Ob5NHltnHY2wZnSTCqJv/1VenvFrxB14h54kWZUqj1HjbI
QFMT5+eeolPZrOvl8FwRHqT2oC8YmzivRiTSIEt2uZV/JmsoEa46mYTPjJTzX7+O
DAfent65V1tUy10CLPu5uSgqbwbl8E2MAawLz5OJTWCuYSp6kEqwzcV6VZ7QrxSH
hD9RFj84/CxQsLnBIQ/QQviPkHky2L6qsGs/LQo+nbhgAGunM4+rAO/vHRDDBfLa
vDmNFBL97v9NSsg21R4hti5w1wYMGg/aM0kUmOPN0vqT1MZPG2bdU2wXWU7bhp+3
UCGpCDT//saElgANMZLIZLWsXNIzxlf90Gab1Jzw2imWgAjql81eh2SaqNOwMqNq
5xY6XvO8ndD1d+f8te6B3YLGRf4c1Z0G5WpelPP4YQusPpiN1U9qhic65h+wgzt6
+NcPT8ShkqwX/+muMdgpZzuFu1bYLY/bS6r9d6SLsKBOeggy8BTLzU9U6rjAMT2O
dJ0BhOwP0ZnRdKOsOoseGNFFzhvvlPuGVqMAe/VG8AQzf2jVtYZMYg864UM5X93c
BmHNV45OK/j8RXLGVervmksUdMCr+3idLQ63kAVnd239PttHL3lACXd39znfo2KD
+FIvyq26E7sV3aYNmSxy3AXaqjFKkcPnup7oMrJBoo0T7OmoGn7IVZA/qmGz9NjX
26bdw/+bVSw7TojSIxggIERVNqZGMgzMneUIEjUHoevqRVzeWMnPuDdybRfmSWaN
8LUxf/R5Q2rJcl8WXZg25DR6QjiL/OkCmR7JFZstkVogfljmltHA7GOkg7HrAfxT
0NHCV6LtzgC8n1cBJaDcnfbUbK8aJl1pZNb/SJ1EiOkDZkL+S2ueeQ0QC9E0Eq30
CuorW0WlpEBxMrTMgesHbpEwa6JKN3MlaPVEhEOEGgLuYJm9IHcOWHfkRuSKRA15
4YgA/JkT2fdq7QlHNJCIjwHLwPk/1sJkN/d8+4ZKcNC8qd+FKrXJ6CRWvg2DpCyK
TDX09iVRB1XATRAUfbX+eQTz60qPcdwCRMimRGloA/eNv4CvPolnlwqJZP45kF4Y
os9Gp0tFBCbrWsfFJz5Mij5RxuKKS7srd1DFbz2ciq5gZ10Nj48YN8wSUfinGbFl
wyqmUmAN+5RG26/8YDb0U4lrurTmHI2NHHYEofi3u33ilY7Vu8UPDjRm7ZkFf3zO
SOoH60qM0lgmw7yZwyhHqb94O9xOE5/wtPcClZUHHV4oygrTG6REchk1jw9ETSM2
j9bBQTIrCj7D1bTqEDBbiGxiOY03dq/3W4RhIKTpDo4xVSnyGAbRzcbfQxhlldm8
oAQsCWci+j6XrU6za6or1ASHCOy3nzX1EXIaXFEtB9GaQ8JOcqhXCjZELFvvkdId
Mj16TLYIvxk/qz0Mk6Se0anzoDz6idVMVzoXtN4Y5rhjU11ACCkl+LxDIEXB9etJ
skBAR5rnm0CW0xfrE+GSdYR7adFIVk4k/OxRg/2ohXvllxWna97BwKRxwI15gaHi
bbO265lZ82dB6jFlsdj6qkSOUVQc9RK2LXeGx/1ZMWYxJuZ52lzsH4UfWgNlSFxm
V75T99kdtpl0F0Sj9gEa64eQ9BluoRfzy83+0+5/GIbUTDrYV6rz9Lm2kLDUirkS
mrJdSi+gRF1eE9NoCVxIZOiKiHBNWNVrtZFto7OhDCUafrZKdJu3nA6JTcgYpIvE
YiMbGJCu0JeyOGZd8G9ubeZo/U8phS9OFk2Mv8vHdwCMmj8ixg36F3Ott6WJ4zv7
JwEHlz6INIHQJd4QFcIXf97mWh5Rt9wQTGNv52EYGV53d85jlD5qOob+HxabUdUB
hdawlEOSyq4dF75s06F93V6HXf0o3a+jMiVE7svC1ra6CJpnuLD0welhf4o/eSkx
he4OoxZhh9iTozcqwa7jtUgPnRafdZHsE4jw17fdFx3NyvulDJcRji6PeKfgrdos
/vKtSCUT7ECsWnPD8i6qfToq4E96N6N55TGVUtl1w1bN/JkA0ncZRq8knNDi9FKz
JaHika1jviU0Db+5QcJ52lhIWxWGxwJGQeIoYU4qavdDk6bZa2Qm0avIIceypNI6
mdArZpa9u2RA0Dy+NgEOSMR9f/Fj60jEAUXzQ8Scaf0KEaoOExpW94/1sfERNM9t
sa7u/ZBF7bfWFum0fp3/3SGb6IMDvxQ04oBd/xWf1+5xL7YHvyKDYTEej2OH6Z7y
Drkazy74MzOyjUafViW5/IlHGDNP8CHcAmI9NrZdQfv5L8r5pb5QQS3jQPLnOUQs
rvmklsLvbh/4PnNCH27/LdtbRJ8+Vv9Tu/XuIWLiVmSsjxK/dVVRzutuwJl3H+ih
53LNSux41KIZnVfpXGdQz9ACZDjFhWf0+rt3AmAKEWPhsgwmUWS5iGRA+c0qKcmq
+enpq3VSvAD0YG8ceLsU2rQYlMnMPhARzM6iyMtBVKXP0oxz2fAcZOBoij/yv7DK
yotpnfwyjimwTT+Bpog6v+SShacFVF0soPpX4uDBgiCVIzvncItK/ZVILvHyIqO7
HTd+z7NjhthEnHxIjJlRoZsZXbHBOn0rs2bcsIS/hsNPGfNG98baOmXN+cDgxbVB
aaEaGzXY0p1/SPZQKRsQLLgojB7XEBLLpD1uZ12CJMPLB9G/4WyzynZWnKYxjFZH
E+ojTPs1eWJR/2RNmX8RpiSd55T5J3Boo+9QchWLJ+nf9ShlvWogDuy7gi1JKuPU
VHkEO14Sgn655XVpHykDHMD/tcTXPz6WdvxDaFULzzY1bj5+yDzx2jN8bNBY9Ecz
YWnSigtkoK+PkSy4GO0fRfm09lsmIlBtX0W7Q/NIlLrbGCFSXKTRtbSKCofELTXW
AizOTLAi2sbVl4voFJew6MEM2I7OP/larnvsK4eSRxRhqv5+SLKGwXoJGbFnEu97
P3r0GrhT1IpLOCICqc/3Qqhjv9h8Ip15UH1ZOmTnWNEIGhO4ztaExiCAYg4OIdNS
zXKpxwxkEpFusLY+o7qvCUE0hPCfXu/38qKPFOVS+FNQEQh0KwGmHsYIW/nq6agM
1YU1oXonJHkHo/FfG+lS12dejK2qAy3hS8Uw/GrUaCbU7nmjVM7KcgPtXM/3Kjjz
CjoX+wP1i0ytqqKeFUYvopBT88MdqNriVOPsyN+J/mBTViNzu5e6KFKLSVJF6c0f
+K02honZUIBRwCuu6FhqQUKDMcc55AWUdLC+JIPRLarIlDj/65glnnUVcybGUxAi
sjRa6ST7vsoMm6pXdeLUmCVO3u2nacZ4UYASH6DrgwJXhj6d47j3UjZ0xMeQYW7b
YVSviht0vFWY8AzG6+kzh+si2QYeFFWSwD0YwZ3OMUnXESPzQHMfFx5fedUp2nlB
TGl0NI2sa1/o55t/R7HE8QcvvG19Nxw1ADSUe0HvD/v3YgkKRWADjteZ6WxIDNax
kou4cv1B0ygSstVCksRRDcv7nKjhFWheUnZily0qrf1EjKdyqeata6lm3qt08nsJ
dewRxOdQASDSqr6EUY7p2RkqUvIqBI6ROB4+G9OyAkI=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXEtG7WUpLf0dc4OCDAwUZdXPPiuNcwDwsUx+8ZjG4QYsBRsEPjffwrg1v/4yfMU
vKrS4TWSfamVsGIJ4XOB4zaV4EZdPnW2WjJeiHbzsFlTfgFlzthnJPSXIAq4EHkQ
zeXiZ/0y9zecRXb0HibgmokTAArxIFkCIXFoRWciU9gz2ET1BuYUoLkeJpjU8i2x
uOl4xt78sdj+BihCTWJ/RC3tvkWMedBbdwuUnIhQg8LYVwaIJDw4/BCoM4Ta8GaA
rFNcnsFtf/2GBaSvKMFHj9TBhjoAdnZhEtlWOSdRMc3FB3jNIY9EFHS0gJ6q6mF6
Qn1KxGaYqTYAyRMh6NdiXr5GTKBlVZzkZNL2O2l+kDSfres1slxONXSPFAbqEoWU
A4soTF7WPoQ1mDDMLfs1AxwqsLmG/AWgoiHW5FEqAA/SV6qzq3uMhXdNu/JFsMAs
P97fXvEGh0OVjnn2cBQUJfSd2gnaUuHDtN2BtqNq+bYoEsY3dpf8Q4D7+PmM/uuc
Xic3JU6tUve3VuV/IRpU1n1chykbcVOuufzPL0SQ9Y1tBgWRSYDkFM/v7CoQiKxM
5GLZ0rNQK8Ba2aLF1I9rvG6WsiSdozzltCN9UrTqbhuES7wyDUAik21EMhzL/YK3
JfUba7bnvjVcAwdRMNFrXfbbXBiF5m/xsIEgOoBBiXD+MTk+R2XaSCO8BuWi7tI1
4vXMiAyfcxcT1NdhENJkXadn4CqJ7L23qh2Rd6W75I5Ht2A4jEDDSa/4U8/5sZR9
YUy8lnV8sbF9eXFTBMVqHiX0EUNI3jpPaUxYvZz6dU6gp1nEX2URg6Zv94mv0Qmb
6sevmPTVRd/xPiHl0Bhom1QY7U8p+Byo6p+Ett/pryGfAp8FVmqvBTCZ/Ixci1O+
ua2YSOkrqFroi1edkYDojXLQ/Da/R8WiizL7oSvoeznAn8F63iOpJz3sdq9IrTks
q8VjPhPdP/regjj/lymzTaKSmyI5T9A/CEVPAya0dj3t7gMK0/cDENjPqbyufYXF
N++43ATISW6cXzmKv8cHkxaU5/i5iY6cHVZE/m5/DGk7mMT3ib/aLbW5HV5IpdJs
nnS7m73IVsRsdRulyuaFUEBX0p6o4bbbf8NdlAzaSy5hg/LWzgntw2MsV892r3IV
F6JquCM4+ViUzrpkLq/101VyVforyppBwd6ERtRFceUINKxkcc0sldsS8NjWR3ao
d3QHxqpA5RxQJmPve1gO3R7O3RykVQfh0vM+nLqtST9kguGTiBewLkapgzuyFxne
+KIIgz3YGC7fYSRmv2yqh8Zv9wkN51ca6OqVRSOJ2/xnPFnRuHnanOR55Yb4fd11
kzyV5/h9iAQDeE93dyWSoSVhtSJ75W+A8YaHonfRSNOtirToaV2gbH53f8yUpfpt
qrAHbY1WEfgRv2flaYA++JL23QwXo5ht62ufOKo7Q/C/EG6U/Pwp6enx84k38Y8Y
pwSUil34sL2tVUMfeWWIrwxqYwMb4wJ94BRHB2m3IL7FGS6jziG7DCZcANTJPvXK
fE9WDThbUha36XlVePDYLqpDwcm8bhZwXwTSJFaRaPVFsF4HTIo6l//X70BhhomB
XuZs4xH5b4L67s35LbrwuTeawsUq41MAsJRGeDSlu3vo1CNdwZAdimHPHt6Uozkv
b0WOLa8xjwlcT4UYpCytwoL6jxG9SNiaTuESw6zFO4KMyyl4qdm73QJm2/ywsl+J
fxY6ym8rzvBEwJO8V9jFV1kUl17eVxqOt9auNksNp/RAaPf+rGoQC2aQhz6G4YfE
d1itOEsejEh17zk8K22oLWsUysvzfJmzwRwv7ZCiqKpBG/xjfHAaqMrgRh1l6UTo
EE6koAArMg2qNJEW/RC8jmEUGgcgJLwxMX28jk67OUJKp/5QaPGqH08LdavJi985
IiV7I70GUlh8ndn3XdOp41IZSlaNHv90At7Xz1bk4mtxCOIXgQgVUar0Aqig+QIm
H0YMsQfGSAfzerDIN8xToHWdaKMUaqI7nbBc+hfbx/BjxwXkIBy50HpN8WKMnYVZ
2g+l/JCoNeZ8VjgUzVP2qwYm43Wnp9N9w0TNJBU+0htRHCyUTWo8fOVmLdWiIszJ
3TlLcs/456C1/iKJnVIgrKVxxl0cClwC+ojAoq5c2HO3B9FD0Pxzn2SyeAqEppAs
QLJgrPEUDsZt95+zhwQ7NvOabyuxKL7KtZuz2bMMXUdZw2iifgvuBkEMeJOek7Dv
eiGj1RvnVKFW2jBOG2MTfREb7BoEPTTa+PLS3bEzqxxO8EYpCYSRQSJhlZpl0URL
9EgdFRMrzVR6bzF4ySiGKGTvYFabK8X8WsYrAit9wF4vnqfwN+hYi2iTTCyCofiS
JXRhnALtM5ZXVzlGVjtoSIub18RasTJ79YbBUItV+nVv5gW/yT/IgmMnyrOISutB
muAOoj0eqJf3KtqVIYAaFbgrx5ERwkWuWPfxTsYAAkPjXFj5qFno4S/WspilAcpJ
3aXIF/PHkhOaSER8JwwNwYwjiBOuJkuWNoeB/KaurBjEUmV7y5NShD+HIlyyTrg4
BdTOcpIEfas44ElKCZBRmXLVLWkZZCZgSJhUWPOB2f8eisG7KDw7G5GHoSb4TWMS
0egDz0cWt7kd2AC1amrtDtuF0avC8mq5LIcPOgsriB8/XWKzhAcUC1+5z1bVMb3o
rbXyJEHNQwTLlw52NK5Kke2UQy+SdkB2cjrYdOSVfH53s6O0neV/NuBKkvUyf/Fx
FxRiyWyFm/38aWnTvJziCmtv+OdlGlR8nKH6LekTQfOH5n28v1ArKw0188aIEQGS
rNhP+cpgdld3ctx7S88kpWWvv/qSU1XVijtvyYo9XUB27qIJduxKPW+cYmtkEZ80
WRyl5tbU8hrsePmKfmmNqqu0BvUdzRygrP0eRAgaWloS6RzaOyFvtMWqYkCOfwtT
wmWzDrt6WPfO9oScGyKXYMW0rJhaLPdkMrnNW2PIMSvqlwqCZLvkOkHPFVZN8X/a
6W8v5/fmyxGU5Ppod6Q3Z0KtDRt4ubQSPot45lRxfNcc1JZ2/qVeBrWiuyAugGpl
3clcdrApwJDKzGaoZNQwivA3qYTnSmp6XztuQeaGHc3Eu31bOaLSMTKiTJlTy5Mt
cthPt7yp7XLc2g2dl0Yh01OTR55VAGAyYhD+s8oO3JAOxR8+6hVgD+fMWkK/4XbL
eHHPR5EaRJT3gPRHSaxJk41lrdte4JOfedptdweiTkjn8sIIqy1sYnOcK0bdSOyp
cfB4z7iXeskFeXSMr1mlTk6gRw2SjIy2OwyrbPdIXlrX6X6kpTDJ4fOwHyTj7RQ8
eakO1mj5TYDf7pRbQeIhEijGCtnEsf1kpLtEuSOI7/PM8bZONebQ7b6lTYN4Qq2V
4Ek1f/vpCohx6Q1gTORVEZqAsbvk5v5+wAescPHOEQmgKojkJ8vDmS9/g14qqg4S
plkmsR3HhqcDr78cEw8ZICjT7yKy4OnpAGo+5rN4ZMEkid8ISbjjq/jki/VtZj8y
rwxzCva+6ZllNWK5u7BgQ+rJ0iWqFjbfYLLGg3e27q/KsC/VJFImirGPUKO/mtKh
WlYnpmAzj6RQBjjnQlLUngzIy322qdsttUMEg8zJsW00AHTxn4cdLTdxwKHMVm3T
lHzJgh/y+qAVx/Q6BK6jB8pTBi0vC42eRe3qX/Daf7ES0a5DjwMoMrqpXA+ik/5M
QIqEQi8WyGUQd/vldUpmrtgXCUQtmSCABC7vLM4Bi9i3g6ZqWd5afb2Tfivz8oYI
0G4UcvcD2KoY9xC58n6wgbbGOJUsJDIymr4hKAl1Z5CSma83optN0wWpKUwIoPkE
rJuA4ZTBhKyYG1G4SOdnoXwaETAhzql5GPDsdM5w7+H0WehxHDGdnEe7SmFIfZ3b
GO/1USODcMpQodJAtZ8L4Ud7DGmtGq0O13X7WyIKaFRlu5fCppL2P2GRZX4xjKrY
DxvG0V3XtD0Ke7vSWlbXsGt2uo9gHrj0qAUvjcf+Qu0rhLsA2HIGYE2+3cVL3fNh
cZYcaL/yX2whcoPHcgohacUjBH+y808ET0RZQxcg2JPBNy36Mxlj4gk2na3R3LZd
Wl/YRDkFJHR969CAlwZ7oGBEBAAv9iDRjwqHkJTZqT5m20A6p8k6VRmHxkfJmQbK
1psdVwX8bwmvvSqWRNSZQ2mbgfRZGI0HycAdwwXTCZCtnptgngETVIZIIS17oWU5
7RAS9pL0YI4hieGQAtrcUCxPVuKXc7dRODbdcUjBdzjyaHTPBz97CVFO/vrW8Hak
Qepv4GBbDDC7+mnH1O+bzSk28/Q8+DNCgTfyNslKw/aUcXDANdOU3aMHu3V1UZvR
RhkmKLRzDPAkncLv/XoDPEt1K6650n6E1BBSc0Wa72GnyYZgGr7uSq0BX6Md6MHX
rfeLY855+5R3HKjIJNZPcH0/Y/HhnW2T/Z4puywX+8tykS5XVu6+tK4n3B48KWRM
45WrKVkZt62bVlolHJE2dqesjnNHh9RlQehsD5dixpie/7FPy5X4SCfqcNn9RUFN
cpwdo3fa93QkFe7IfkqYkBrzMG2dz70NPoRDzL3RWlIJCvy+ok5Jsyzy+DstCkca
8csI3dhVnWIWv2QaDaJDpv18LYXifPr6vBOYOk7uAxqbYTtnmQo71jyxNYTPMhN1
UfUTAA9spFDpP3H3bmSbfZkQMQpKpvtomYWE3zCcLnsiKalNnJjoIbwUdRnI5NQ6
6TzUTtTiFNXxk3qRW0TA7eqGgDSG4mzplVPa3ATXRve8ZT7Lkpk/Q7JSI49HuVPK
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvLX0rS/OENLjOTJaOMKtLcOkW2Hnj/D6FE3g4ICZUB7WzzmqXCix6HpD3NG2QDc
0syFN2svMFY201XZB2Ch77NcvaT/mTnWX6bwhD5+OwnnyqDkBWDL/FWvmYE5IFoO
8M4ywP1pHwC8yU27V5ZnjI4A07GSo4adoLDPVjAtwI0L6tTAGpEqSeDmsdvAYYS0
joi8Els4sNoZFVTP5zrAlySP5jlKNWSmIIcfgvWCEV/0Xg9bv5SiyeUOUAznvVXK
2i8hYwUY8nJG7wUbgHthVXr0xtik0oHhZr/ZIouHVCK+XmFOX2UtH2QpF1ZaRmtP
iFdHYMxzoG6qXstE5uLlz80g42I7wToYndu3BqNSabGcoT15VQoF2042rPLh9Ih6
uoTQxK1pI/5CFXpFOw7kvg==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aPrlrmJmr2O1Dj+A5HgIqnjwin3oJYbrEfJNph2gbljo8RFpDrJxm8c56/GimnpR
DSa5hT2devEYVVFETipHsxTvpEWjcEw2aWnzWT6uid5S4V4XjdMb3kcPJmPq6jgd
wiUJfeln00XB9xIhid04EH+7LVFwq253FqUIgE2Gk7CJiqa1YMekDGgGu5rJplXT
F3WqcwhNEdpyct73ep7CTTaUAQt0GTQG7j+xLkVgHPamvUbg5raBtgmqpP02IG9Z
T6c8kby6LVWIn3Z8N1WIpjFbmZzZX/8xYj/cJGTo+M3X9HHBbDaTDVUpXvTHXMuh
t3zgT5GobnP0sFFH/TiGrCQddQqcSxFW4GzcF8BuhP0bbgFoY81SADu/hb50qQW8
6UX2vwCYQ+/XAxTO/wWJWYlOTU5Vy8FWYp1mpqYeH2OYfK2X8XA+Ymu+33T/2R4J
2jlQii8eK++hen3yN73B90MUNdil3NDR88CWpyaOL9rHt+3d7ERy6+WrF6sKR017
O/eXWhAISz/TXbtpw7EWHEvXxIIycFlDXBs2OJkvdmnBt/Z06N+bSk6oofMy/IVo
vInbMPrD90ox/tmRbMCDEnnHVumcTysY7aMV97a8tMnJGonVowGyccXQTG5ihm4v
YGr2/GM36OA1a9VsbpChvPoRbKQQKCdDeoaE+lPJ6+eoxbo9btwBloF1zhEzypdh
0rsythG4pTAeB1Ra6gZfRpW652eIwFupisVkf9qP1oHti38x8DevD0ySXdZ7puPK
14il9usvvHvowLKc6mYytrh/AwpjP9r9XXJOH28OaCBfxZUKUqC0Hy6NUBDaegYG
ujBmvbeHb2UFqa2vAOq60hMmNJU9LYh3Q005OKHko+IvvRlE6LxB5+c2XSOI80b9
umFmN23gvX4PGy++Q/XiyEZbtUZwSIZWkXX9A8geieS3WXvbFqaR3V0+1HHZuapE
v4Y9GC/rsehGyPi74kLSQDdFxgVEuHYj++WTSjbTguEX7DiAfNTWfnf5i2S9+Hkq
fMm0oCL7kb0JznN/F7b75r7ISOp//uzjse2TcIKEXgpGZuqh/LHyve6rgfL8h6G1
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mDYls5wTeAZ07aF4d/BNfXpFBRa9T5Jtffw9B2RTSsnvJXiAKh5EtDdyh5A+ZKg
Uyux6Eclbwz/j5ZQpuNGwtYNSSupcxmL2eaGSUWW64zjGUwr/rxSh367oEu5Lgq4
MJksiaJmf5uCCOE4OdHaXJDH4Cn6m+MjlCnthhzBw8w2Y0pysV8Pabq4Y4fYI8Ea
oHdL+34VY6PDDwGthfCWuLyZnWIqYyo3HeDLJSkZJiY6thRzMG8+rSNW+z3VR3qY
KsDczNOK5SZHDPVeT6JNgaRYgLf4lvwJQPDO1c7fxibFMoQqXiP/nrm4w3hou1F+
RXjeXNZPsVxJ12FovU3nxjri/BM+OqHcG4ubO+ZkaQG4Szk93/sUnzfFW2oXiEWm
6MWLrfAWQV+EwS9y8FACVfdvBvZsOZP1ZQb0FJuu34JkR9zSKJ/irdWcrZnmZ72i
HOJgcuorGO7KCIkQynhxj3jxbnXKcDQ5ZRRXwczACEeCOkAzuXXU3mKJWBTVjYuL
UbLWnLMVKqynwzsiJzHE3f2fMHDHXYVtNGZspJOhwrUESsWZVbNELBw8eVeEWyI6
VQJxwQTZbJzFG0Q0DHszf9wIrpJOaJlwiSUTV1LHrHxkVxINv3x5nC2z5qvN+wo6
NRwMRMXvIsU+jEzxMVFbCgY9q/7pWv31B4NMXLGXWLxyeLc7sehGjrlU/tM10FgR
Aka0XyAGG9U/q7OU4/XtTIfHmHtFqS1naaUMcZ9npQuQxOhGhhQwv7kidBrY17bA
3iD1qhBsybD137E2MFpfbfm8DT4QdsuzdutZEQnBGbdMIPlbIepxLpq6JkWM139r
Y/yvR06iq86szUaIEqwhoVzKQeym4PiM7VCQX6jYAjDK5d9Y2RZCtEjVS1Wg8poE
kPnyNfoPc1jL0gILuv1Kvwm6zGl209B0pbF6eZ+RTdMlgYQKRzYuMfCFvwS3hELK
`protect END_PROTECTED

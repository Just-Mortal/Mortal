`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6yQw8rk8Pal+xmzjcEqdmFlqupiyS5u3W96Le5NeiCsdOkCQq7v/fDfNIM2/97gx
7hHYgLH5zkGX8bcJVo0xoOxUXjSH070Dzih4MzgcCwoe+BKJf/T7Vic6Azo6/P03
cA/WkIm2m+cJEddwH+haTMYzqbbNEvQsGzchj2L1xqTD6VQ0esDOCzGCBWMjpfma
vaXA11w6i7OZgqXXBcVZsMh5i6W1j+yZqLsGgSlqunngri+IKPg2V4JxedY+PzRH
D3iOlj0RdzXGyZKbbTrJJhs59vPRKtz/i+Gcq0HFyRFuyJwXDLV7wmcAWjgysYy7
9P8m6lL+cvsqZpsG1BbhlqP5me05mwjF/HILon4VNL9NQnIreJDWBWI3LSVgD4IW
f/8zI30xc/vIBjMCddK5UW3kVhJyRsnhJVt8qSnT9kIUsReCBwpdprumYIWFZUXM
MF/gvR4DynMFXUauF7pBUtgizgR13icsD+i49fkq1roswg7SGI/8aTL5JBY2wGtI
Nd5C4PHL4v58TzkAReuMz7XR2DLsSwD9uIwsKFIw/1yeIY47EEMDkiH4zr3CzJe1
LggHPHKKtherRUznMNI1249GN8Qtv7eMs/PgOAGJO1N22T2GTyYMzwdah3//lLk8
2ktDf3GCT2LMvivDQ3yMPyBf+qRZswMjzdu93RMM2dHL8EyGx3HaZh/qut1GUAhG
sHQAeQ03e8+UMQsE+ztXwTHDAFqUzEMgXA5K6A/eSYnRGmHJOJgOh92vuSTa3Px/
qbul1Wo5HNPwKTxwz88W/mHNxhRWfEBWeNLWsPjkXxBcRlv2K5pMjQW/BDqodZ67
wyuQP3Rwi1Z+/afMz3Vi0odfOvikrYq4+5AcqSpaGT8QD0c878Jc7eYlC9kWCVbe
ufASnb83s5nGWKniWDZvqFkXbdOtBx2C+pVJsu4GzoDowoqB0Gk11jbx+R/VIMAl
qrNDpz1Gxk3Vq/zn+iQPMuPspcF4zR9EZ1K7fNjz8hyMq7bPopLI1zcw1qph6Wbq
yKghQ9TYlYeBd5PQOCNjNbnfSfkAAiDtZ3bwdQGHXPBLkyqy8oRWWHHS5dtNfyAF
HtQyDWPEA4EqTt8ba05D1DUYf0u0XAcSmIBSISNAwukrfjolF8qWefSiwu69LHDG
rDF5A4/ux3CLRKiKStoJ1I0JtBvYra27+0WwuZU92WREwGpmcb5IOfMKWNFirE7C
N0RVj3FctV41AW90Z7LJgLWEehNvrTqbYIZAH1+BGMa86tsHp+3Ro2FrfpmF+qex
qmH6PIelXTUotiDjPgaXi7imcu8DnRkAtP85pvvbcsTlR80T7yJ4vhb5mhQitYML
kWzWyOdGcRN4JSDKFECNLhtN2R0k9rOoKvndDswR4a9B5MuFAwPXwk9fPTDhOIhX
mIWWh3ly9JpNSHCrv1hdVmhYr4Pc9Co7+zN5ssMyMo2CPchhm2LhqekLPjBrcCn6
z6lwmS1VhRnb4EJDeEpjg2FXepVb3m4ckozf7S68gsy/0Ed3Ub3oBKlbhBtMy65T
g8oCYhrAA8UTg9KJCM7vGBJFfRAs98W9Zngs7rb16w136pCPWMQQC/ZxzBkWTKGn
NLp+PuKEuzQJGVGIyiie5IxdBQp5Bqi2p5TezI8jhTFNZJotvkv98gKnaaTb6uaf
64RXOg56UtyuwNfdSQ2AknhLbwwZs2UN3CbPZwPr4NT2To5gqtP3UE/WhITetkls
TW/P1uv07p4XKWhQ5mq4yummwUzrCvbfBmFq9VaDkDsyTJLe+GB38NHGORvRWGR4
QAZ/LqsFquf7pjvuqGEOtGXw/V8k6ex1c1nMOJkJhbzV4wyApAPJEarSzjeFt159
xS57AN7NVrB1MultS3bkgiH8pMRHTuKDGVTsxmtfDKbqExpv4OAHrrFSaj+Gce1J
oX7sM98tYbW7YK7w8shbllUQPTnun02b5SWEa6b99uL1/O9sIxaYNp4RU/dns9El
eN8YrWq+WdTFFiNuZM9AlHYrG/o7TlF0T1EXDVwk+QbwzvVS8h2OT3Qp+i5pVEif
ucoWMZKeCVOi9mHwvP9Y5BZxoC+EZ9dEZKG/7ET1gNlEt2RVLo45QX541EuC2S4b
AX1j/ZdxFBWNNFfymu6onaEIjH1FH4IZncnwC25W9frv4FRfr4f918EQl7cEPjng
zqK93z/x1Y+6oLfOKi+X4+K3ZqdqSbuJi/X9MJdHePg4rVADJnnkAbI7ZbE3R9Q+
a2MzsjbWHQpYNbyvLjshdbwh6RifGwtkRtvOtMyz3IKl3q3CelPgWgUOC1rdV1OE
NxtT+p55u40fPpjjWJb1DdiFmfWPdV/Ypgw8+Vi/Grqd+JbKaYbxy6Gp+1hnHO4B
qc9rOm/CiwnusSOhT6KHFCtjqETsxcA6bD7QvBQEzLxmD8gsOQKh4yuiBpWeouIk
WC9I9xyK5qwA+Ebyb18azchTqqnHpoIFdMrgGS4qp5X2QAOblqLXLc0oXu/GsKqj
o++Zuxh40LO77CAYZYiO88LQUg9qYT4Y+awqvWjmMYXDuO/B0UAgXkIQ+L9V09SY
dCea58CW42uVWPkw0mvOTvdRH2WKE0gxR6vQW/1bkkCIueQ7W9ue/iC/izfyNIvv
ZuRfqUKM1QrDKf3+CjibAVqekMInL1gzNg3f7OFfV4X6XWjoOjLc0KKlQw4Z3m6U
AhKI9JLdBmEX5UaiQoXB9iLCOaLhleMxlZlQDIIPxbUTnu/rB6cBY+/vmP9CMzxs
OwF/DczDTCZV6+Or2c7bAsPZoYu4D6nAN78+8hhrMacgfgNneQZ/ZIEMMFdP66mh
RdgNUmQz4VpoyyfRQbr68I1sOO2e25h1Tw7fHpvvM8TTp2pre3YAtbAacOdC/4OI
JOL61qtH3iMfxlrMEGpJPOPAStCEEIZ10b3vsqUfHB1HqYdVsI4wUhvZ8t9z7WCw
MY0O6Mas5YWwXcx5xRqZ4n9TZ5KRiWShs/C9fuFpdOo+g0urBwJTglVeJQns4K/j
zFmsHrf8tWoKUU1LB5nHetj8fQGBm6Rnc6MlX8EnEj0Ik1JstfBE5PepKYQaJ4F9
UnnOntKauR5iO8xKDWuhk6Ltqo8YW4hANFu1pmy0vZTc+5g4BZZCAuoWFjbFu3UK
gvVtQt4k3D4CAoQU5OpKvh9Uvc+P73SOA8M/1NnwcPIockaAuV0hAASw2wirgKr7
HhRkGOENV2z/iigY/MNrrKJGqLQ0Gfp9nU1/bGDZ82+8inYMVujvV2A3Nukdwmg/
1mWB0fgJOONWlwncexGPCjhHolCcrEJNJYpNT59XyzQJh3ppsN8dNPRY6nKUoah6
a/vqJ5/YS/OqDyDENWKp6IdXMOU8o2FHGF75PxY8kLvq4OwCpcIwKbG7eCeWXbk5
ZoRufBnqBeZGPafCPVJNep6GQQu7iOMgLvb2JjDQJtnqyON+xTq0PXbTALvuo0Fe
d0OL0324CugLP5Ytd6ELRzh/KQr/rDLnClGz8LM9cbjJEjjIL0eTWatHybWxnXB/
6kXSr4QlNPBrtGZtxq9IA5g6uczYRuOeEG9mmuzQETxyok9AE6/an+uhZi7XuBUj
PchfLrptlT6Ktac397ig3lmoyNpnFSA3uqEr3ljV0/yk3UaVcEm8Ka6VXifR6ftp
NJ4OEZHXR+665nlClVLYkU8leC28ejCFhsDawNu7uz5bbkI5mIdgl615gsWLs3F+
XVHruDOTCtVRxQCtnUMur54CvAHHE5NMs1JwuXj2UDzK2Q4DQop1uzgsb4Y7Phxe
C6QoBYa2RchBCvPDgDp2VC2Lhbt/WjXaCHnQfUdKXA1no4xgbc5V8tQe2/aUSVwS
ABmzW/yOS8KcDniW9YjyQQl7Kdm2N3MYQ3jhMxK/DP2hoccaAycl6O2KlAMq6boX
EZJSNIhPljgSHRwnPFq7MZLbd3OiHGeSB4cji3eqNeI1Rx4QUMcFfTuJq0NZ7oeP
ii3KIV8uHzXQMKlRdjwKg4MDlzsIsFI+MOxcBCQdhf3hvAEsSDhPnxOdDaGti74w
mR00WSbXpxZrpeTC9gwR/qo2AcRAIVJg2LoEbJ2altQWVBFu6GFVvFh25JSjhbOl
39u/SAdG/FfCVt+6h137JzlBBOGAIGi9S5Fn8855MvQSGqB6Q7nf03rn6fwxB6VF
g2m+UnaCJoesmvWhQtH7Ws5EAzHhuGUafGbJINbQJijlaetXUTGis2ET64wgzkxQ
pb/c9ciKJuXYaYvp3k654ydBZ0glY5u3yTsc+tQFb/051Dc1fmlu2+ltFJYvdzrZ
C2O9Vno/BwfFaUDPeP3/d1ApMewJdj4M7TcFEnl9qO4YLgdLOp7Me+g3nmx3XmaG
ZLGoTDVvGCCR56/3PtDJ1sLt3cLhpjwQTtFGE1t0ra/QcrWJfTuwU+0oD6iqm/tf
reTb2ijoKNP71ApJjhIuHzlW5XBPAJpu0Rm5ASGFY0qX5NPOTLbCMb5jD7feZBhz
V6WUYub641IpaBj5bBHs+SRT0gNwZ4UKQk3LVcEuOLiZwVutqgof6ZfGD31ohOjI
H2eDi40jsA+TnUYKoLrQdo5rLj9Xumkdso8UJJZLMGYBl9WOJ3IXnyLMQXWj0cIG
xltsLy07zhFfK5UtEFVmMEAWmQO7saKs89Dl1VLyqa0HmkylHiWiPFwXMhOWhKDf
WsC+rF/ASwm9tJjIrFcPSuB3yf46fuc+6Rfk4TBa6+iaeRVMF6wUsBpKfTGBTzO7
Mvuy3avrsUOtGigofDx/OF7wdG78d+imjdEWRJs8APEW6oRih92XyC4lt0MNgMP6
hUtj5uQLBrvVBMDb7wdMp0nIstF7um++C11K8IEHjxYsTaLjGnUYYLAKOYTOykNY
s6BjECDEXQ47rOlUa4SDaGhk0FAU9i66rJJagBA+tyO9tEx7c9jAq2dYmefIfinj
9YIw4CMuftw1wYO2gtbknQj4L5lv7hayA1VDSz118MbKgGcmqFdvRsAYbyCvKVzz
R0ypWR05Ds2djdJxcyylA0q0jQTbKHnbUcwpgxrXrz/qcLHoWujYwhzoABR+qZI5
zP+1weE6RgGkhiPY/5W8/+dTiiV0O8UIMkhk0Eg2m1J5MTM9R8SnrPMDAhjBJE3+
Qj6/0FDfp9SFqtRoBFwM4ldEstB1H9+kon+dQS1kKDuFsPpkIKGnoU+IrGfhcJkw
XxwTVFF38hQrCV9NzHVvkeSqpuIe42WLAmk0JokZRCsilDtOgpmDZMwI3SASJ9fk
f9nbZ2mbuxY6YiQvtt++x9SGSgfJHH/0GGTiC3eNZJ9DwMoPrZK7A+a34qxtC+Q1
yw2mXukXR2pwBR72UMG0bmtbI0Yr8AHtr/UR72vUlSL1Undhgrev6V7E/yvRkJp4
a6kHhfm5wpLgLo81GZVJuyxn/S/PwC4X5W3gjjjCPD3XlXlCpJGPh+vAjPBaurHq
y5WtYT15VPwaHcIsCqnOb3qpqYNziYdn/cN2TOcuKSw/PDTh9fGBYVhLquqOaaXx
y7HLG4PKy2rw/NmivzO0bNx2vVKn3cc7v/1pOpZSJVRoQbEH/ISVeo/FJ9MOhgkM
LlFPKnBKRqyTbDaybL++HMbZOwLAU697K1/sl8QDwlBmppV1DHMvZveALdrucw4d
tIgZzEwA+2xcAuHENv9z/tv9WwZ9ThImR6K5XvzrsR/orp2U87zsrvywURn2oUVE
kumvADZ1hBNGjgG0kgfFyEPjW01CZo7TRoYG2JA65122Hlzp9OLCNXhLYmUUcUOA
T71c3+1Jm1TBrzVfozNDZhANvAikw9gbXs2g3uinasgUQLiZQXmXYagsjhPs23kQ
UpwMW1U9XqGZQO5/jaG2pq+EpnLyPiLTr7E5tjQPXJuiDHuDh3K0ZAjBw1/J/hrS
Qrw2V6t28j0FdJpqN+Oc3Pid41wRRKs7EEyS3p9KqNLr4bTyjaq0tMjN4g/s9lox
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYtS23HdCGTka5iHExZzPd53t2p1qgu3grfGXPXZja5Vv1PMRfMtp+5wSN8Pvie2
Oz1PE03wgH8cnCNXuJ267Rf/ZBUT+Oj6F4UDfsupocKFp2KDbS1p6pWJOZiy1Wah
Hau1shvTBe3JupHdg4839pmLSxuwxfwy12wKCGy4/5rFYdSH7ioRzCqhlJt8MwF4
R40HFicPrXW58e8tx3LlEX0et6nQq3j7yl2elwQi8cyaWi72LtVQ0RzDUdbJvTDF
lucQxiwUWTtzHO0pV1Ly3kQnn3z/7VoCz+7oPbHseJWC12SqBULu/AJmC0crIxSI
2FwRMy/FTPNDMr2OPZK0AHo1E1ttKR85Jpr/lRtJEOsPy0I09bpKT2gnReEX5730
kWIZVbEtL2DXTzRRVSX7Lm5Tuf3+hHZSg/WI0e7Pu9XFaHGQMx5jr2WE46AVdaPD
cVDa+LkeCTndhgch+/fNArfz5w25U/KWHjAWetMbdfUf3mfvYiEuiu3jdIL+SoQQ
4/LXBQW045Vm8KomFUHhbPnA7Zucf0wHJIOyjwTDiuaPT6BsQkOxxwT6UHXoVuPE
qh7Zx9mIHfVyi+n/7kwUo1QsUmyDFHver/JgpV8Zejs/8wgXguSJZoVZ2Xxb85zY
NBvaG++YmJzMyvqU/cczD61u53D3uKwzlEvfbwmO1OuTYLY/mOcSKowGckYd0P3A
3ISJ0+ADmHVSvzdBH6nNBJq35UIazbufc5BQD9I9boOoR9W7cFMBAzhmX99T29oW
AFi51Wo4L1Y73H0bDRLf4EN+8a8NBRXjgYWOQMMfFbwwZEkJgehLCYZ4eo5K679P
dgTzP/sCP5axzFjDwYD/I5SXl3bPt/hujHvLHUUbY/0Upg6J/v0WKXUpCn2PzpYf
wSK48HV4KfkYmdNReBy/j/AFk/SzNzOVCWWVR5Qt+NI9qQqwEVQ4MZpbmy9b48Rn
LJTz0FiANceMgC2U5mD+sNrYL7BxeOMQRj7wYr+EdXfA4+5NJZ2mHUCyGhP+yK3m
1PeHTI197JhlhfqFE1su0C0DkUQX+e8BiCzTYXq6OLUhYLFrfT3R9sROstrALAQ/
JMWcKyhMjYO4tfXx4greDc4LgeTmub6OdqPO8BdIiVxnaAW0fBHyXvoMY4uujkdU
sSEe4ZJeDhqy+OEPS9zgiOuX/gfIb/mlfxMAWwFRpKvH06/u0aiCr/0dXQQULqIL
i4nLBKn0iBx0MgbT03aNuzYBBVVDCjlhcOexudIJNQueIJWvpb8CmcnfFID3frXM
1R423YFUP3BOKwmkXy+4yHPQUWFfyxgS81l0qzhInAehCndv+uXv9RPfq6eqv6Lf
mjxsGuWZ6Pex6i5IhD/Xf6WWHrF1s/aUlf129kUPUejYlMAqQ46hmLImQwirf2mW
ZmW2GrDAAAuE2D4E4L1Iq6hhr/6bTh8uN0Ny9vyshDiPSgIWNByjuY1FaQm6mYEn
P9F4UrBaEwG93n+Ktmp/xXoIzKsqxqduYvLZ+gms9kD6buE8P7gOIv8Wl685pg3d
HEj/6VqwKyrq7W0e3H/RgpxAAUAiFoprwIUmRcEQvqRnoxLYPSEO/5JHuhy/e914
sn5TncktX83vrJaua9M30CrbOzt6fPQmg5xwa3c4+hzcL6XTGmzuMreiyNCJNhQL
FxFPHqlCF6nxhVMQvZ+zccin33/QYPAFNdD37bs7mGMWkih12OcOJafwBUaCkeDM
FLRXU1rwVBVFVxWHK0lCwfud2vB57QkfU70Zu+92uTMXhanLSlp9+8hy7vYqTQ90
s3zul1nlKe8Mh87uPtOljABy/LfxSJLW+NqINnA64k5KzN2SFNhHWyIpJhRj/4j0
b5KNSzcUROWbEJ9hPxb7HJxqHi3sceDJnSYXBeU6+MRc05gO/npmv8+7hjOsNXNx
NQRQglhayMtNeBFalttvCp0Kjjc+eZkds1c4Hgr9nQwpXoeRga4aKbH25xaCRUKm
ubPtd1LACPzM1qLu+ftQcChq5ZvXkX47PyY93lq2BMjKntmynNGUzHrv2+dgWp8f
hD1qfP3Hx5dmpr65ktYk6QA55dFFyODTzlSjbyEcBYDi/zrRv/Gq12CtcDNzrMRz
ju2S/MP616rhTqYWZnDCYwhc27Jk1Nw78zqrBc9JZ4Y1Cs25IooXTC3CmbMbJKtu
l8bqWZFc/xYqA3AdFsgbx62cLJ+vMonfMQmi9wOXPmpWXRjNkWEZ4hXE25hojpka
a6YSlS5lJpmN6zYASqU2OW3WXrZtFqzCIwn4k8sDyTq/xSyYT/Db7fU9z7fohVB6
g2t4T6ryLY46/zQ2d7ZYT9nFjVZ0lKnHfIrIyxSWv7uo0t9XNRoxWTQVRuHfC0Zq
mmkOYaFmmHDH2nzmMNOSlwL4mN12eT1Ivs6ELW5GLVkmwkik5QI270qBZEe4f/zC
JnXbfMs8D8SfmeeRaNCQpuCzmSCVQSD5vL1akq09MM/goKyfDg4XeV9v+26O3f1j
sEw7x2xN5IgcK0CPu4iLnvunJ1jVH9sOfygzLmLVkdg7KkDNmcVby7lxjjG+emwf
/oQFCVXweq4ch9JiP3vGMFZZpmeWXsnB4y0XaFlbI05SDfXpvhktkwLgvg+GZavZ
rXjXdczw/0ColgXdBCe9SsLKYr2dNsQOQfusg4ND8bLc9fFYlNd3J1tWYFXzHQP0
6UcgFYZ3GDep0z3f90p1Sd+lzf4/aV/gZK7ehY1voMOCZdSr7/vhBk2K4eLT/Kja
5R4JEk1d+DEooKSUoSiqO4076ntr//ESewQWrKTrwXzt22/QX+fbvSj0YYEZfSdO
oiEIBfbjW8bKQoOCemNpbMU2B3np44fGmpCpx59TmUxbvJrXwbZieNsihtv0NtNA
i0OazgpktvA4n3UGKqlNGXc4oj3StHhtDQGOLml1asEbtAvynMfl8iPzMAp/Y40R
3fOB27fplcyCGPHTd/x1nce6bI7fVHwaM29p6CQOu/mbf5W4iEK0bmNGFfk7OGOT
rEK4vwg4bnOl0OmAQsusNlfTRuMUIYOvEsD3rX2G4p8Ksd9cfh3vo01IP2NIOyLS
kL2Ok1pQlWOhqWcE8k8N4ug9Uxi9TKAamws5JsyvijwnIdjyLK4nviTwEbQKh+z4
icnMzQaVI0x9BqcFBq0Rc3Z00E11oecSDgW81pgkd463//10Q47RTYs9ZpDk3YJs
CxdQRPBL4qEkTfIxtPUgLMfxEeVPNEO1CpLeqYSQTDDW9A0Csx5LGc/QeMC8ogUa
NrUoWNrWg7z/1zRDvTBWrBylpqKJqfTJ92hNAPiugcfSPcPP2CkPpWVkBaXmPxHf
9ehaXxZUI4WyhJeLn/i7eGVDsP1P5bZzn1Q+UFkn9CPAM3Z3a0frMCeJRM1rqf/U
W/jGkofXU16TDsUjvzJ4YOOMvUlYU4UjEh63ugw24MRDqvXSqzZulKZU2gcQAc0x
WF/OgxJCKXWNF4Zi7Zgi/SWEBKT0MuSaUuSz0MMZtyW66L0sABwjQTqf41WBiwkX
BpWNu3vbtr0loEdXXlqWGEjsc7JNx7tAKa+JGZUMIh359eVnF4/VmazlG03pUaGv
11KiSdm4u+eji7vQpHN51cb8lhpm1QZC33tWdcLYajtwIP1nWSEc8A7WYQNMGZXk
fSeKcpaIx9c2sw6HNzl9UfsAlc1BwPaCbjWZukIGGDBpE2kLqS3CX9cDd98VQF41
H9Nln201ESd6AVss2kZ2bkT/gNZPTk3mRz1rVtB/clrLTFlWYVvCeLK1ftwx7+1U
WbPYaYTzVEYwpzzXIJ5AUw==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rf7odKJ6ScRb4Gk1IUFXq3PfUkNgSkzXFx1UhJkIScD/jHvsVBJSGV06W9PBIWv
xbjKhoXXbMXtZQFCOjAZE7Y45Kan+4NXKkUS1OAMR0iVTQJq+xTwQDf5kEjZPsVV
eRxEPqPVJudRYD2KBLcVzIvGc1HejgqSRLYT1Uz6zwYGxQtjuHRX7zYTwhLKTIhv
EchpiNw2YZapnyp2rDgBKaeSQBq2BsMkThXxa5kju1ZvbOnxU8mmIuGZ4rCbiyeA
oCEOXHCBCSCquq9JiaECurHRM3d+8JbSF9cBIvxbQTVQs/Al3FynRCuU3tNI+mVc
I3n29QNPgCuYUVgAWn11uW1gAAxO5TfLD1iVWXkMUOXGCM9WH6ASzxXmQEYst5hW
+ZAw67JUyIbgmy1tf30xhyo247bWWZQcXVEI591z9nHN6BxWm30gJ+fjGolW7eHv
IsVn2ZGP8WzdyBDXyl1P50eng89CYZiPYTy8yTDv0lQ6C/TJrGnYAEYQGTIdF9BS
lyly1+7HaqqdPGVJcikl4OHD3P7jMwrqrY4SlNFv9KhcAwpcvaEbsVv/JB2aWPJ/
3RaKYF+g3gS+Re0/S6RUDUiWVDS5f0KeHEGEHTcqDUjAY7y6d8OWacC0ctv55/5x
2MIMobQi0Fy8Vk+20GSYdMFbP31m8Mcp4CNQGi5j81ovVrVgcp1+7tzNtAj3x5ZM
BD0MCubEPCcRM51TXw28lFcnXUnsirsuFqw3c+2BpZSBWb14WCUpaWplXbcbTOx4
BBYKgEva2yOFITnM65k9Pqxd8avkUbx0K6GAeKUonytP4rDN+x5NdEeruG57jBH/
no4ShGccWwnVR4NySGQeYsTRjL76KCZopAbqpssxI47bihJqoKoZ4orjXB70EMCy
8LzyQ6dnyU7hiw3hMtZ4XvYpvH9S9J/0w8TvGvfcMaJ9L4BynQPsFWwG8UMDwPLB
GCgeVn9Bge4YUtqTBvSCt/U/0PdvN+GFanVWPpdTv0vYS3bEOs5FU8MBilt8lNB4
zZtLDjiEGysIxI1jiYrkMoJI1xXzLK1dsiEo/NW2u1fhDpn16AsHci7zyMGQoWzQ
2M+7KTnbr437cJGH/jFZXRYTA2KDKO/AP/hqWbHHt1pWB9C+JTDgs671oR4dF9eH
ZEPsa1s6QqHTHeKTSzN1IQiXuUclyyscWEskTyG+TJHoV7GRoYCeowKKAjSZavbg
MA7HBoAgE98XiIDFPuqFRQ2DSJ/p9G5jRaNNoCpbDgBIZ5vCFkIbK0ejJUu7TMbd
Rg2df4wSQ1WvrkbIumTzHqd0bOj8mGdf8scdrsJMy7EvHC5vvUdH15X/PEwoTgkH
tuBZTuDmgxc5ax8QTeJWk0WCtU7cD43v+rF/vdCsXEtFiKpG1qNSkQ9QC8ps+ui/
i3ddow+rebyvS3c90802Ejzb8JjLgu7CY8RpCNYdJFh9ZXT4DQmmgcKdJ3P9smqs
ehSR92AP4h64nWpbsNBf+uOOSVyfzkeNQsAxWdY/V1nDCwWrM6TFIISQFFonbcct
Uglr5ex5jvO3rhnQuA3wzdY9VhyI3fZmxv38KvpuWbA9m9o1GgkmNS36y5jNrm9t
I39vocLIbw4yJMWsWzQGXQgdIzgzMMSGUEMvm/Wk5B4vq3WWCIJanf67IZx5bYh8
ay2+JKX0vAiatROjTEPH96fFH/aueuYEPgNV38yu1IKwFvgLtR9K4sq4h+bQCCRq
7Skw0tkPVIugJW/FzSR/DK/Yks6H1job5OsAYJgWh+Gq/B1cw+/NT6sh0BjXwG5H
Gh44qfv2jPTdLPlnloBBCxZhuKFsgeUZzs2XvHb14bOZC5R8w5FKop9dF4Ob28O4
9DA9uYhstxarQgpCtlD4r9g8VuBh8MwwelXzT32Axw4cu5QLADisb7e1IwPW5vks
bvMF3jDCQrDAhzEE5M+Uj8Xi1+Bp3mC0cIY8kFCrrrpmz91B8RD7PNOoJCAZT2WP
gCNFQBgtshXc/sr46x9ttHuz/vvPUyHheaCF+MX/qUfWh9ViIQ9dHMtCDk5bVyNb
5NmmCuEFvHJop66Jb9WQ6CQBr8aQC4KBs8f8OlBk80CTyw1ih3z13y0J7G1Jqz26
apAgM2ik5EYwzWNednjZ/BqVb2+QCyqIO5ZlRRhsyofzZY98CmMhGGfohAaNLGz/
jWiZXQs8wSS821St6AVO5YnR9KaUZ7YHBbotOpwjQrXH0lL0goMPAeDCc+KsNa9J
J812QopnpjGGs62tvZLXD9CYOdCd4MLNV2EoLMtQMiRK5jrvo1QQsMOcvuEoHpWM
Q48SD6W3Re7ZsQQkZueGOhQQ/+MwxoQ+wkP1lHRv1/lHzO7c8taYAbTVpYhPEpTj
YyCfvwaWfwnzTHiYT/+celioEtG0SeelhhWYmKUcnHtDOTg83Hzg3NBIEP1UBt8v
tPbqXUrmVcWTkZ2W5PybJ5aai9BjOKxo4VDTdL+gZBIgLJXWr9FtQosp8NVDGDSD
IyC1qk3A4SWR6iZ+GLIflbfJwHFk4Ik4YWSYcEcXSSLXM4IkEFYYn92z+vIsuaW/
SAzTcFDONMs9zntKZADEVvATxYTpMDmWdQmWaO0bFTT/TqG4wkZoDVFuQuMxO54s
y1vtS7Cp3PJjsB/bEBQ5MtdqPwi7VitmtbgaxIC9czDcPTklNpb3m7GfXVd4dXMK
vmOh4pEKqu2UKscyIHRUea1mt4vvp4TzaXBKstGn1HV6WplthhQcaZK/eWQMNXGU
efXrS33HNyj2HfRWMbezoCQ9sOSVlgFSSLeGQdTR0Z0THrzU+5YOHst0A6BsUuDM
hpy0ErKRbygrAOtBWFmpLQs8sExHNoZrg3tbEj8F5UX0gVHpQ00ppwsU4jz9SRtV
fH7aDaEaw/wtMiW3LqXiSitcUPuYvcKEbINaI+6+zFrAojwLsGqkiv4wv1qnXXWN
iUrkzY0UmqYhdgupO/WiUg2XhHfOIu/Qw6qIpvFjWoCjlglzWTicU4F7UZ8hf2lN
pFrVaFvZWFNvwZiG1vEkwtvjxsIF9SHJeTOL5MLASHPl2ty69ZlNOjrtHWMUBKB4
H0kB5k8kVWkrbJc7QGaUjl5yck/rfD4b6TcDqM6b66F8UD/Q6nFwAmAkeDmnmxhG
+Lk4J2MjKtvxE/yQ67fK17WlcNBHzzBdw3g8DupyUZelPCU26H7NkOJiHWWFzbcw
i4JV4CrT2BDCJJLyHAjySuUSqvjEN0n1xHR+jfG/VmMoGrG/uZPO0TYCO7rvSdIl
8oOISOz8CCzXjzyT5Qu+dpAunwG4m4sEkcPvtsPax2HeqGGgkup5/mDLUQ4n/Fp5
BHy0NHH94ge2MertVvb6TOeKWzW18+9bHCbt1en/uuPYdjvl0jdJFDllqrNloorL
tTrU+CguqF+cobhwz5nxV9edpWGvjNaYBe2+f13e1EbRQIDRSAzMc8qzS8AkDN2h
7m+TC2YXSjogCYP51PX3zTOL6aDODhBuu9wmeGoNgS5/jHMuhs5XSrD/YT4Vd0/y
2AAvd0FvvAMXMAhpxwjzP5f/23jfO1rIzygxxBV50sgmHEy6su4KeUttxlhRWs7f
cTc6wsnkcGtjrzuXTHs6A/jbmBkBiKwnc/p2gjuetCwPysUiDVgG0A1cD27k0N6v
etBIn5KTFGcACB4+PUMbZWaOIx0LMLk703W/uHwHqQXKYf2c20D4/aHVWEwlt+/P
uQPIAaT+VFUEb5TfNP8gvqgT6z6DYZrmSGiUwtbJ4BA8Fb4CoKi2hLTZ1zyxMlHS
OT3eQaIMpiglrYgaOHweb5Q3DGLdAaTkezShUz6JkvkJNc4a8bfuznoo/tGZzJAm
buskvMoHnqen8jU1aLOW02BZ5UArIyGTjc+uLq6KtddOoGbahFzuYz7GSh9O4TgM
pISPZY0fqVB1Tg3kQM5GGncAMKfDMOqFHb7I291pJLwQihxMctsGbpMeIfORhsn7
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nngkB5ZiwazTxIF6dIFEwlzhbVemPEi+ZWb3SzEdS0ncmnzG7SSwOU8SlWDmuOwh
6ruOCNhTXTSBx5Z2J98+EoIwSN/Q4FTfhK9AO4d2LBGZSAlI9xMaA3lk3k7WBWzh
Rf9MU/wXxCK8ZSrFy1tLFJHkaADsICtF+uzaCBOVn5P49weL3qdNMUh9l2TObH3C
zS5fRec9DEJBf8njTX2hn5RU7ZBM1jSetjuHSht17mrFtbI4m97ivzS8SaakarBb
lmca2XyQrIcKhpu5TtWUfiUDIiBY84UlSfDIse1+VtlaM/WXiGlwt/fO2j1+nfKs
7G3hySOLcnA4sQxFGfhIK543oPrG78Zets7TmHgxj7VQAS6k2W+K5abj+FhVnPP6
OVSdKRlBLrg5220mW/iJPMODQ3eorpsgcJN6/kB94IWzKlnslEV5Hbn6Zd/glF+Y
CqJgdlz3KpW3N2kfZiF14hYJN6GQeR7nWRmnYspFxYtbNINeZB6TBv55PlWd0ycp
MBNKIYJhk8qfXxu2UloU21wSKp28uRNsuKfpltNvL3oAMhZM0ph7WTEsDNCzzaeR
uLNARTnvyUd+kNNExqYd4Ism1z/7ygSRX/NzEl0WBIZJKiAREJWd7Egh5uQK9UTx
Q2XFYRGNHr1JzIq68pj2FukRM2zGcAU8ftmmgbM/cWbnRVUmsyKPENMDDB3oZVcX
1HYzfiRNrRoJtzjYgzTDFRT+c0y8rLkbTQTxFiEbGmoF+Wz6Gs+Cwe2zWgWOYlJi
zyikXNzOzPcoXNjOi5D21PKpUfKkazDa50OUJY2RazGhh7bliT6pM6m8hKG1nduA
DUM3MjKRFpwOaJtQGEvb7DfAEyN8kqFW+odhweHOX7Bta5WuYnvQkgrrK77dSbsR
8NXhikcmc7xbMJpV4T7f1cxphNhQb/cal6cvqNQep299oPxHBoFd6VeMZDBVfWCg
8HzOystQZx+yH9YtOckVZLG3AD2tYDzdoGfMdbIkznIkQhR+M759zBO1GrYg80+E
O9aMJHAZSAsZJINaWNItgEGW66hGuPRfGNbFwUxjSAWgpoV826ocMi/O5LoCrWB9
n153+/uRYvRzZ5Lr1m2cB0MjA5/FUaiRfrF5E38dyPdWnNIy9tkOww53enUF9DCX
X49jdye2vgbClZCcLJZ98GjlxZEI7KG/LyXRnViFWSmfaIeUwkl3vBVy7cWtQWY4
qOG1wzdTIVLV8SY1ygN9AP9o8lXmqE/EvjvoYRnhu1VZHieEWVk4sPRKPsu4RW7P
hTytWlXjr6THEXbo2pIQdiZug1HeHec/bAeZMRvRxvP3FXiBWa1jICQoYjFCxU8m
wKhRQQiNGIt4K/1Hdy5uxUmvdFIuzxrEgjGwCdY7Gfs=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yE349CDR9QigTZSA7T/DDzfBnQtCOlG+qNbR2RrF2pjiLu5BBM9/I4PBCT94IKRe
1Or4wtnGVSCyYI+DPb4Igq4zy23iWJYt80DZ2OiAOexcLW5XnrLsEALV53Ug2hBC
X5N7nGnFA/WCDwLmeetS3+1R5S833VIEHsKwzHd+LkEE9hLsnF+qTbRMEe6cD7Wu
C0u6eiuO9XOq/2bVk2JxI9M4M3MVMVwaQFopCfPssclC+myIsvIGLQTUMNDr5stf
rYcwIomrPPsPYQMXRIH+YKWNnr6lwHrxadCRw07TGckQx9m209kkgX7HZadE1Y0z
R/UjpNH2dGPGDOORWJY4xPkdPwezrslgoE7pLzDca0g5RuieVI59/AwiNEOolyM1
ryYLJbxyWX4UyADE/PHZBFqvS8XbXDu4BDYRLcDiSfZ40lxQ0y5fWinerCmCfcFf
ZXu3+v0DZKy4YDqET6JWbeX+8LDoH9tXjAnRDAFlLTnuacCIAWVMMI9Rou6IPj4z
yQQN+MygSG5VnKxoLWy6jp3xbad5/agVhaei3tpf0Ul4vAY9JT8/BDZ22gUtdFqf
pNIHzP18UEUgHsEwDdBZl33EoxeimZ/5zzuxYX56zQzMr4uzvFpzV78JSn0QZMUA
+Gscbwht5peZLqb6HZleOwfPMECtikn680LJ24vSPN12tNzogr2dOEXMhDKh4G6D
oJLL99hkKEfvPv4a3oFC46F8bXHM/UdFSGxPNxac2t3glGqszzjq15C3pnnA0RDc
EAwZub/pFhNESqLTAxddz3HKj+tP8yGi7GgyoKZev3Ac41YbAj9YakUUcMucHnUp
xVTVcQ7qqnVKPDP5sgmXciSNuO438ZQuTahvjbzDqCnKzvn/uAPHDDTgHZVCcsNb
4QvowUmr7QKUIjQaLSoys29F7mB/FqH5mYGcH//JOEp9Yo3Q5YlhhVZwH6xH0SgW
HTMdNdnC9bL3KgGYkNOC7Ngu0skTrl/mZcjh3yZyWqqcbZSBfup6wtU6RdPPztz9
DYsI/G5tCh7+Naba8RlnrhVhYQ5GnkKam2oS4lZwIs6udIqp4w6gNlUaylbdX2v7
XLOZuAhuujumZH3w5nMdPNwxRCbN3K5skc4GSs+v7EyrFvD+UMceMz3fIepcaoJO
MEQHuSq+sHWIw0zqWiEIkgfY5TKJcEsM1a/AdjUWjlMxQ36CuS5E5Kuq2vLsndtQ
i5lHFU6X1zUw1cI83aKQ7vRG7uJDyIXt/9dQWGh9ODbqnsKoDWj8OLvBFLxvAyWf
GBh1E1/lOfE3WtmZHXCEsxHNFAKdlrsDIdgsa8xhga3vk7OtznxUVaL90NxQBLPx
R134yccPk0uI8Tt3MxXaozJy6lk1sqypJdocx0729n0RgOaU9wQkcGvL4SM3qQSi
2qg/2BOdD1Kz1lYFhKsOCMsW/LpcmeLDxhZ1A3sh1Z8QXQuJ5p6onBlPuJL/OIpX
`protect END_PROTECTED

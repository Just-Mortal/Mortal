`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvtgF0s1YbTAu2s78ELw3HEcH1In1dkWIirYdVIIqI+t+DeJ3XJeWUW1CHpaPhB0
JlSth0JrxARNtKf3QpJwekLYkCSD1thTh7amkgfDCFbW0HzVuZfdEYDH2wX36pEm
1CqdVnfhxCoegOEZtGs96kv4BhjOMTC4X8FNsrBRZ8kaa4h7zy1jt+K6Lou8DIQQ
bYsLec2xa38mJ9jZvVtJI+XSWorsyCgii+md6MNwsrjGjVd6xoLNBTj4j/B2NN/r
egsLPtZd/orePhBlSRz0Zzf8c5+YBb+i9RpkruzuafFo1d46Yes5vaYe+mkO0JLr
IX7lKM8KoU2dLTrgml3O4hXeylZikvLgEl92/OHZNapNzu+GkDKNTeo0dgV7k8RW
PzBUxtY4xDnXvksy18vil8GMJkzHUZt3c8iRzqspLW1JMMtsd/3D+pSkM7QLT1Kw
7ZD8Tk7xaup8LaX5uUZRrep4J2eMuDRIwIxgoCX8e/CcnbdH+Jt7Vv7MhGBMtLDY
1q5cnoobArHbUHW4iBFpvkdpjdm5wmFSOgcTrSJ9al9/Xtf2111F4V/jJLa5X99I
9P5Y3IkIHbof1GXBTE6va3xNbcaXkYQWoIlBKzUI0hngwNgbTVEQQHfxMsW1qmPr
j+nE41pxepUeGxwnhL7Q8I5JFpCJZHkUlhYDciVsFZ52okxiD00K5iVrGGN4NATk
jEt5Ub6FAei1O1oqVOQoBXfUD1H+0u+PWczTIt4LQvtn4h5z3TpIy6tRT44vbLIu
93rFH9WAMP3fsoSG9V1D5EUjz2x+FEkVlJ7IdYUWj80eOfvoQiroRKqyAlBJaUvg
WYPxpTUI+fl8HKk7iKPCtwHomM4I1Ui2gYA6UZtD38y9jx6D+1dvBOi6cDwAGIDi
CqqqmO6PXAjO/3ZxxUkb70NrpxXupTj8Bx+Xj94IaFeImb7HzxzrgW1te5CdTmxW
0Lg+DbRiQHBvAQ9Apw5del9xj77DZAUCElzUP+MsWeQ09BjhwuFu6PQIYlUIAztg
hKs7llu2kD5PMiVRLYhSpdw54jEEijXhcN0aJTyT69E5yjF+iA4xCmZNl7zE88nL
C4BtbAmAoppdszFJMQJcmaeZ6iSqgjNG0hQHaYn/ASvqXvZeBGGh5Q/X4gomTKOI
dByMCNJD/5XXZd7/dwu1R58FJB2/q91DdPpUUNhjvto38INzh2iDu/FlH/Ar25u0
VTpPOL+M9zlKdXPsjY4MTKnF21EeoK415/+luXC4qXMSDNdLhY6XA/lyG3onTMR0
rp9FpoLd7BSa/ACh1GMNkYOMNUHc2We99ppdEYZTtYbR+3IYYKAAuq5cMkMoHQaz
rmCqo3Tv/m+TY0yRN6fx8x3LSRH3rQ0HcxEwW2kNwbDolkZOs2RtC+57Qd93p7gq
4o/obz33f90QC/++PTJ22ofn0U86oFvKWxr6vdRptjlQmupCD49T3MLuy/cYgF6q
EreOJ5fQhBGy9DExrAyZNC9I7kenCV1Mt9a0o+Irba/UBPE6HPrgsvkK+LwNda/N
/5lK/9cJQ52upudFtbuGV5uTjBEBChAzI1C9/vFcA9w63ZBRDXDf2Bqe+5uCRF4q
pWH+qkSQU/exoir35TO6Q4ZqKJViF5samZxQoXedzH86DFeb2yfF/B89fZ5shysF
0cWbggrxKXVP5jgiLb2w0FFi8AZy0l1vpAHpe+cPVh1rF6zIdIQ2Zneq6G/EvXgU
F2vhWOtJ1Eaq0TAiqJ/G1lQ68xy1FiHOeB1Cowrea11TyiCNCFhy4eE9RxD8uKAH
E21U9JP/PUUJpyZTZekAw8VYe+/UCijQN23+0PWY5s8wo9k3wF4n3qbUgw24WLNz
bSTA069QU3H9C8TQCuN8Jgbo0kr45hLzM6JeLwOR/vGruxSM4jlkkG24/OBhKQl+
aqfYwjm7M8KK9KDNt1WFXJ62btsokkCVDQW5SoJ0Irg=
`protect END_PROTECTED

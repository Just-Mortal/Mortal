`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FKKaW90QdgRyPy0+QrxlKuxchGeXgTSmtGy9CVB5smV4lAMjGWXoKTdjsWDEWFTK
6dV7voIXEKSL/oyEu4BJVSz76GwyE57PDZKChAKi9ON1ILsZQk0LbdWE6QIDTOTk
gmpNycHPqoRPm8Eod9DQLFF+woNTgIp8vDcC4g7c5i9DoEv0ReKAG8iC5U/rV2CL
NI10b9wBA3l93VYh5QjVEV0hBZcew28ZEuU4igw+j4PJAxlySKGyr5jSVfNxbQbH
j5YraK/GLZWbrMgkWJbbMqcSu+QrEJZMub1C8mKjv/g1TclvN3ZkiZPhHaQpsmGL
Wbxep2JeD0h45zCIlDMYXNZw1GiJEVo0r11MEnvCbuerPxH0kiDkTm8cwM/d2IqM
YG+x0bgUh2llHAtTw98iJhndCsSVX3mlBQ+w7Qf+/iNHLGdMam8X04G5scDCyt4X
XKW8jzP3eeysx4NXRakQyGRzU4jhjOHgpN1HonSbRclDdEXT9EH6ortndoIY8s42
OasdFhaS55DWQ0tAqiIqWFsJSkfpO46s7v1Or486OoX85OoPxk7whdTCE+zRa+gf
/8UbwJlUDrI4RQq9sLW+yeb0X+A/14pZHPCM5ugLpOCmaXs+M7EZgfZaysfQ8ZJH
tb87eO/AcXwuc1SvD7RrdPlFSn/YEeN4qeFe69eTQ5WmTGu5un71bcQ1L3uviPDD
roH7UBl78M+mVtvMIOHogVVqCWZDBmfSW5n+9altryiczWAnHrCci0dn3e32f+WQ
8tlJKnnffuuDONbHIUriGF6RoUuwfG1ybbt35yFzMYYhg6fg1xoI36nVoXkwPEtP
lZyqOq+IQPlTrKkbFdZRThM4DrRhKLCTy29POBifwKlk/6A6JY/niaLef6B0B2+H
KVC2h0W6zlEEXrlQpw724PMWNLg2AeqadgkEXHrrnty0peiFnzKiKvgDKcbbNtgC
PNThNehxvL60ffz0JriJsdg61a2SSGK1DJAbjC6y0MSZ8/uxFLSIQLWqYZMBzSfQ
Y7DvLu5W26TMIxZloh7juWTXLpabKUh75ok0BsAzeCbqqfSIa+24nij8HUPWKQ6U
lG0IIQsf4u8FVAV15iI9d83sau+Vau8inpWOJ9Orntq0dsrMAhC1tD6pkWk4VbbB
ylo1DQdsffkj3HI3Zly1ewb/IYEXkSi8ZGn9mqA/Tk0zFL0MsmZnn7qq7r8IKYmq
mg7BGBOzGnsVKIqLqH2h+kt6tqZYHU9B1nA8qANbQWLntf8nFD46FlXJ914WbHff
0eSxU4YwLtaprWvszfI35sSMP7wCpgnycYRI+9JQgXUIrKbS2xgR5PDVISl9XofZ
leMSlYptXTwb3kEYZSaueXGC01JNuVHnWj9TRhFNTvCFq6pcEDPGrt48iby9QCdb
8yYM8DgPIrsdTv8e/Qmt13mbFGF1k06UZLJINsfgnpiAWdglJGQShMmEHsmTvsJe
z/Wq1iwoR2zUKdrBLMoUyVI2oVKr72KNttvMHYnd8rU4jYI9XHBv7DNJc8r0hz3r
YagT7+AtXfliQ1u1NAbZwTaV6IgKhdbNljVJAbkytRH3jz6cZ54BuouR9X49kmnA
UAvCYbzyMCaZSSSvVEoY+OFGh0W4sm1LkhUHt5/d7XUFKL3AGELx/f8J/cuJWRZR
NMLcL7Z7DGZjuLQE8sGBctsiS+VDNMQeUyS4iIma3sr/g/SmdXp9JXREQiV//wom
B6Rvo7lBtkN5+R9xadGj+d5AmjknEFEZ9suGK2/hsie/XGZ0qjpfjokF2RekCrSg
8ja8OwLnMOmbbmGEVr3jqjh6rof7golQXr4QV1qxFNQbPCzRkAe+pdjUgqG48ZOK
P7d6XJ7Zowbg33K9CGVi8fwPIK/6llL+zndQHfCOxI1JJtbPo5Skz4Q0/yqu8Mly
ElANIHvZCUCHKGuGfQb3PPI5m9WlsDRIC1xy7F8OwbzvVkUi+nvTNyBdgDVVW2Gz
IIxs+3V6tMtOnyL9pLMh+TWy6bEHPj384wTMeBQOIAoeTtQJHQCj4G0NVflbpUKX
1CFhY0ynrARmwXGBlzrL8hFrEAmycVij9NMf/Ojanum6w73RjUpjGYGtCD/DfhWH
Hz9XD9SsKHs7O2YTSu0CYhfhQPDyw1NWbcAhCAwS0SlgmOE4GiVN/n4JahklokWr
yolsJrnqzLnhWwAxaI5OsNVefEGF+M2BKnaA7x9STsjvh3DKOlZG16wnIHNSNqoz
K8cMiesYm/JXjNOlC8rqsWpNkdptXBvWrPpcm1oI3LEbXEx0T8TycB1y/zFZ7xMM
n3hTmTYWQHfCj82JwWiiGj9hH/5ZJ6P71f1Op39pxwwCkeE1efSRGqLLGbMU4o4M
MqCpjzpPMfHCcdTPkyfF63svFlzxN6JzBPejueLItXbEGABUfZ2G8/an09bWiW1O
7+W9untWdvo3WKlSvFFiwxIF449dQ7SZ1orO9HJWNSGP81BvxHnnnPestLUxwc+B
J9akeEDBnN806GKQKXAwx9IvBM99RE7seyhBiTOkPzrkXxJaZ3hzewsZzZtwqVxL
a4DN9cOjaZObSdKiG6romte9bRmu5UNpj61zyhWOiIVyDpkFGTQA9R/vWBXZwuiK
fDnZzQLAoAvKBauP5f9emOoMJ87UgU9aq0q+Q1FwUMsscOy2UvzwYDMJcEdjXgAC
yWO7ClPO9z/EV3SaG2rdLQjb3VrYwhrCGUDREVSYDDG2HfFG+UTEmdwakx2qEDb/
FOgi602EMNNP/9hr37AK297iQhMrjT/37xCax7xPTwQ419uH2tthIj1FcH1LWZd9
7SqP7D3sRwEiX8SNGwDc6/xFCqgtIDZJB5xEEhIe4Usa6swf5EGm9pROeembIVG0
goIOHJJDPOCrioR5HB79N1ram6oywV5AltQIzr5zDVSIJjMjR46xRrM/fnpQISex
j91cCCdZ9ISFSqANQ5GaBBp6T9c1G1DRC3NMdRRrLfkSeJVdJ1PVUhiXC7X0R6db
jk87KBrFfWClryKBVsNCnOm98pfUcVYaFbLeS/g+xf07ag0lu4wl8hTdZoRVtFGr
4hbYsW16JLMFqs9t9eGHVOKhOrU2/qDwx8+x1TwrUnTSpphOuEaonNkitcGUNBHp
PCOK31zKgBvaePjpfm39Nlna+EvFVNOEafVHFTJsyhXqCuYwvtznZwlVpOc56pu3
jewQZ1LqMu9RjDJ4IsJ0/RiBfwtoNG+TALJ+9KZjw2eH9tqVlQXyIbmTQHwpgK3M
gpZzYWlwCkBlOfjsAV3oWLQH+jVrb/uOZMvw1OVxGW2n/GU/xAodZXAeMrFLG5IM
lHWg4iQdWLIe5wqFu0tiBYtxk/PUcXJ9LvgjwWn/7XF4x0aO9eBXk5DOgwyR0HUe
A9qDrYcjIeO6AYuNc1oE1xFGjZyjekcli1NeKhinroYpasDR03JtOCxjfKjM4NXZ
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GDvSYFqiLJw/9XASptqktIrkOmuneoPowIUbuzEDf5vwmaqpWbBZEGBA2AeG15FX
P/e0Dc6+NZjIyzdpjx/qziyuj9wA6GgbxP4qWGbExR+QhaDKlBYpNRSYPqyBZw1Z
PUejwI+9MVq6vvbyJiXudFhchJwDUNVe3A8z0PUBFCrTpdEaEqqEZzl3gSbHlYFH
9a1GPjcLMhRawJ3cUVU83eHZInaRjfDhBHz5sr3c48AWMQBD7+BWqquXtKkzQ33Y
DZsP1xIbRExq0SJ12SKZe8hsjSU96R2LtgBUS4NmhEfMvA4C3acMuOhQ/UdEbyIz
FKFPo9a0OS9oTdoaL4I8k/NnhixsCKWEVqaiyGx5zu6UOPiYtthmZZvBRvPDIg7T
VSZdG9Yn6rB1yqCUdbl1bQjaTKVchHY7P8Zv9lo9+ud7zBujbVVB+e7YD/n1JAx4
GByN+KdPApoKtffEaUO1mv/AEAt4R+f1QNWVqw4wqrq7Ez+HrDHIEOdECd0/Q4+l
GGhY8ye1Ec1UsoBBV8GUpcgkO1faHhroCdDKV2r4mcyNwOT3dvlhO9Vd7cFUIAH3
2vphvptQWVEnpmDlcp446TES4Qd6pwL1MdZ1oe1u90wnsOAmE0c+SDJtx0jmwcjn
jK3NRkEjPNR8FFAmqvEi01hbkKQHtDrCqTrFTA7Lsdpv+OfOHtLsZlwgwu3tLl3D
wLv0+d54APzNRljmlo0scQ9KrGfDQQymCKUPRTXZd4O0g3dG4dfsXHu9P7X2APk8
F/5DoWQ0eUh7RVHdav4Juc+GqcgPWUqX48f7e6wB/zMlo5CPBAm5hN4MEfwIk0ei
mjlkAy1ab5Bjsq6+VYdeMrdM0HUAe6jubIDIrZLZwX9Nz9GmSmee7MgMehJEUr+A
WY7at/vdJCOFY+P5/WdEDPz/1frX8cYR8498SWIbyZrxF7cA9SNFDENr0cut9ckl
Jd5XXr8oxLGO0e9hdBbhyvFbW+eNshKyqTLivjsISW/yMfxQPrWX35hMqbHP65jy
gktQPhTEOT00eAil20xcyplYdTnEfaoA+wXp2Wtp7Xjinmul95ZJq/IU6a/idiHF
tTGWSWmtFfPiP1wnuAXQD1kXfuOnarecsUHwdnTTYWOEtrj+lTa6z9DP3Qsa1PGn
dDVMTlpx41dvsOkRpduIuRwOzWDCpbC91QY68tw37jObBOJ6jWV4pep2LNcw1LVR
oQM9sQYNkt4fHN3ptxF0iDECGbddWC4Pc/iaNBwfQRHU/Q1uNkkD4ZdFXqUEQBao
nqPD3LiFXmXBz9iqaJOgBKlgfVkwyxcHdId5tqj34RItUPg/BqRRgYvuhD1gsj3G
LWcTdzxjUJeKR74bHA9ODXFWmAlxewaHzDT1GfV7R43WzjY0n43hFixi/LvbrPQi
MHAnhGq2QO+dCb58VXUCcBUFJrSjXG7YObM45fAL/iY=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDErApr8t7RZhRiUe9r40NF9UW5A0GIIMrxkGy7qIO5NqJgWxI+8MH6+/kI/gKS+
NZyoskQymiEZvBFC5UGbVjyIc/lIsGxqpZvbQzQsRQGB9eJ+SYqCNddKbfwohqhT
QrOevrxmGZ10FCl3boVPzQ1ogSFpy1XW/osKKX5887furbQNpKeIVA6V+/orke0j
uoHoFD0ZVmm16Im1t4yxUYhfKEHM4uPwDABV9tJUOCvx6XummoW0aEr1QOMfvky8
kRX0VV5gaBOCqx29IXUdtyw/WBYC1/I5jQBnzG4HC3RlCXf1B6NMuCZ83HkRpf6a
PiayPnBTM0HWai3SkqY+X8NVBCEYWF0G3DhxkX7Rq1SYBxXXDrfrU5yTbPkAvW1u
+MucLwO6i9xBFCHoC6wshjUGdjjAAvjdG4uPOqzlN9i9T1czwhDSUfllE3Kg4VUI
GpTNotX3GNkWn3PXbG6xvyw16bxiJRpx83h0MnOhKLz0Zco3aIA27lVwX0DPDzJZ
YhKRa1p0W2mqXg+35HiDOfr++YCxSxpK7IJPfbc5O7C1B1lBPNIan9ClNe++yy5O
kM55Ev7Zp8e9HT8VQ7MJkwgI7Da2HOg9tDG+VOma9Jfz5jxbgu16gfoD4RZa1SUH
z0OtkDMp+y9iYxoYUH/2XTAInAsOmoI8Xs7JK6P0E45mZ+f95hnuNhx/qfun4GZm
3KVBLLF5gKksPi7uDf9aJg8zSmhXFKeKBuBWYTyhqm4=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GaC7zJPQQOueQG2XtFp/jbkRRJefbtwHHQW8BARqA7rf5j3tngBRksUqVp32fxJ5
ZLiJC9vFzY96so+3aN7uClCrZ7JhmwaeiMtZTMOKJJovdemOW2hpeYmmty1L1oYz
igXH1uK7uT+K7L1FAJdHgot2ZZB/R9cdAgvz2wEye5yPhW6I293KSWpoMy0D1WLX
Z5sxiTzy/vUrOKgZp6+xZwfLLDxT+VZmfop6jz7y2rfF02qLb3n3LafVXtsBqz9W
6ZRAC81Jo04/Pppq3iTdG7QGmcIVhjsLHwosYwniRrxfuVTWFMDRiiXwQEUL3lr/
iJa2ekTfGCUrz6R6AfbpnbuS3ZjD39nySQCx0flZ6uROyntbFkjiS+nwbfyS9L1o
/BX2ysoAzcy+7ywnaxQ98ODBlZoHbwX4bjTJ84gek0wID9P1GiXiriDcrCuOQHNa
QrRn+Xw6H0d5xN/1G4UWunmvye5MqttkciNDr1W0P5/jxHy3TnFGBdlddAALP+c5
az6q4LpUbOMyAM5O59mDn3lW8FEwgVV7nF9V4p4giBEhkYdKaZXKtxo/yRZ6nA/g
WrB0m5UgCMUDnpIFfGFJ4EyIWjQyeVow3MSxGZuw9i/qLuAz/GBvtPWGlasVmYU/
CxeRijtb5QPCQegU2gXzhjJ+MD7hJQZ8/KghbYaI/kCAl8vm2Fb2IMtw5KwOsCuF
WVppDBCwM/3PtG1iMquKOG+R6FXFx/+Lt7ULJPdWAZy21OBTLQYlQ9S93LKe0gkW
xQOE0/DiUix95Ad2HffeGcbrcZiKosr97S+BYAhef/Xme+bpDANbg+Wj6LHqHVOn
yiqyJMiUIHu/BiavyWxmsbx2el1sRrycAvsYq5AEvg17Xa/6pp8ZugcpXiiTO4BD
QjFJMoZOCYgF01auJC1Ua41CyBr6YnZA0JlMqUfz1tiiSbJxw5oNuccdk/LkXS3/
1FsvhH4BAs3VH3v1LPjaj/mOGTln6WgFhwbYXJD9+xdLX9qMROWKWJyOMOoasCXm
G9wn57TehV2OwKRDz31ZxdywAFJEkmCdNrUettOqvvO1KddmPNzG8hQJVvY6PjCH
sXw6x5whVhiQ77DSroHCEgB4XJmq96uzVR4tdVS7stujH5YlokY8HUUGBX+tE1SQ
SaIjHtadTYkSaXmdAcSAk+ZakRscTX6r2HMMJDJ3wfKXTorYdWH8aCJIoC6Vz/rK
r+iKTDgW5GLsPwFRThTmzE1iq64MmLq7aaaV7UcnNZbZHYYBEj5UOLFGGu6xGREx
jy352NJiSyo20skgI8cr1VOhkDYqfedbuXvfGZNT8ZHcBrzbYrwYjAPO4Zafj0Q2
fZkCRXf9RboLntkad0q8NI9YxsZYCUEYA5Ak5Yd4ZEf20zHq2xECCrCghl+ezY6f
JaK/hXlynuiy7zvcBMlCSvkbopVU6Cr4/7NNvdVE8lNdXnDjPRxx+IFmGbw43oZ1
2ZUGGDuNiWrTI2gYR6vPg8rbbL62QPE2tauvoG7gNWocwsN/cBZ0iFuZbkF/D11r
HNXURU734AglgRhI0Q4WZYo/NFNZspX0W7vwbS2Hn7dfEwtoYm/lUdqmWN0ixXmA
6u5cadOkv+WgXsFHst3jNVRWG2VB1ejirMlWWsYC33QMX6bcLmZPS2XA3BUpUF5R
cpp3GlfMznUVSmbq4ykvejUPEaV/RH0Gh+txUhK+Fpn+LK2s2Bk+z/+AgCFTJ+2r
G2LLl3J1/mqI3KXeRdJBHdqisr7DdCa94AhF0mc44H2rTfMU7VVZ+QmahqYKJhNR
KaHH08FWuY4c5YLTH5ZrJgo7C1bOSlAqYQMEBY6yxseL3fPqNrd7o1njD3vlRnTy
ZxayG96ME+gCABCwLmiIxrWzc8qs9HXY5Qk1yyoedD1jKb+ffBgWM1+rQ+9Kn7k6
GFS+gVePd1+DgadYIGZ7huOVQkLk0ZQHzD/BG0l7o4MvquwvSNcXgll8Lm23RMk4
rCtBfmS/mfc5Y700THeQt4GaergAVbSRFapmOrQApz+3Yn+SA9csFIix7u/NlgWA
xZ7lJRduLYzukefxBtZFzTfAMRpy0CkWf+LAS/iTHGeI8m/lf7W2ccNKWrdSM3Sr
MvnERBf8jxg5tPXOa5STMxaWdT5mKQ/ygostNvcIkjWIneLbwNuph2FfAq3sLISc
6p+RaZ6TNSpKSwu+O/8EqAVu9ASSYorejC7kx6uOoGAJvFsVigGHrxMKsafU9QZ6
mzY94ykB+TqDhrF291tB2PacUjn6qvAXrrKsMILSLHilj3qIYm9LZTmQaHZKnmpD
44DxoKbTwOqbqoS6wD7knQl3ekPz7jyUGX2KzuomqJaClGIhZffr0EYzD2dO0fXZ
WkqFP2OT3KLkJsSA+kHiE0StTFOhgbykkcefX1I4y8CQxRkbYnhiuJbwEfN0G4UN
CLKLzurCnrXXpKAcKKM9tQxfS0ROCn/nx71r3TpDwzFQBfrnDH80x7csvkbD+TX7
gZ4aFv8tBkZkM4lzBoYX25R3vN13fDvEsIbE35wWTroL/Uk/cgG3uu/SjCTCavhH
OIyRY0fCMTEtqbFZ+9X1pDfbSASUhc1EGZXL6yiLZfMkyOlBQTQ995xJqXuNI1oM
to20EmJL3sJUB0kuVmR3L2S61gbovgQS5HjzjlHqwvCZZnl00JKZu5w3/4JIv9Dm
CwwHoqHd6Eqh+KfmAvODmj11oO4VQC++FugluMON1VJ8j8Pl0zPttOzwfgoE6Hcl
4Q3cDMJ4MyK7F2AJmjDTE5AflTf7splASDQP6R1N3WX20YT2HrJ5zjXt6XZxKqth
5ZrlMApfdvTI/P73pLFji6q6igwRwjr8ZQN2/y+Wrd8xgAytAEUgSUxn9gaAvfYS
TEFxSMuNAaNPArUv55UV6FkuWEi9CtWNoFlHTcplZsjZj3x4ikpAzQWD+l04GXVg
KOGUWHp7PjBVd5BAT/zPaOqx7r3MQi1K1YtBahxjpPV6FYJcTOhgCRFfr0EFAKRe
bPox09SVAVdZieVSyBtKbsMDtfWtNRxRryIcZEIyp3dyhisS7foL8wSjZB07Blfs
P9jslATdYrS4WXou10nomoSmclGecf8AK20j+oZGNF9w+Qm23umibwY7zJsSuivp
Nrm3b2CH7GHI6FpRC3hKsYBl5xEdHZZGLyPDwBcu3qyAa6SlLe99UavUBzSw/Vd1
fVfJUqQ1V327ZOmuRphzUgE/tGvF8S5fiG8VuvbVQtYYUQwdgRyDXVj5U4/Ep2yB
gn0czYEwMu1yI+r0eYaXrDraZkIIGyphN4n/aPysxdYEXaHEaciza8oF+Q7PMacC
lAsDt608oQ93vvWDfES0Ek6EnTk6t8g3CtSSBqwHenrZEHIDh6wWam6l3QIq/Nyd
HGOE64eKdA5D/I+OMaWcrJcCIRnVGHX7Yn5mI0ewbrvWQkthWAQjev5dC7kRhybT
cKkosXZ8EuEPJfZK8Htr1y+BFDlKeXFvSVYoslpdCRjaxJ5dSx4gAykwKiQLYj4F
i3IkL7sQ8uBdDT7xk+OKwAVpeD9NtC4xgeTSWDm3gcpUE5bDbsnDQMfaqsJwToPZ
imBTQXANVvl5MqkZvevmEo4KXi51hfJMwI44gB4xOyBdWZYj9r/EKfMuAEr+gBLc
SmgKlDHOCfzOTo3c1ihqG3BMEj+rYgCzEpsaHkPI0tWPQeZMq7+WN1dx9EHRwgaz
Co6hXIPF93mHkCJLq7Cajwj7Q3URs5PjnDt/y9LqeQYgeOnYs4npFC1Khe0ZgaOZ
9HAx6Bvl2pPtrra8rXDCjfK271gGOQSUGEslZLk20t2aVNjs8afHt0Sbuy1JoMwq
qs7KaGZ142grwXmPRkSIu2DLhHrVrZ2rbC4eHOC44Y60MaQ8oaHbkGwZhRzgnUrN
m0xya3ezg2f5mPn8TuHwN7qMnyn0/oBi28M/6+iF5VNR8jWhykwZlzyCvnTDPGUJ
FiZREIbNspzixKJvyAfnKWKR9Up+27iCZ4gMwCc6/S/rD3qzc0fC/H5DtL/zlMbG
yeF0/GIkBpG1UcmW9EXkaAtvt/AT47aFN3nA08btmJvfQLkz3LO9EVhyQUQzodGN
7hKPMjXS2Od3/Bs7vsZoRpE4wzAaiZH2T3l4aUn2HpdkG3zT9I+W8gZoFGz0SltW
+Ci8WS+AYdhvWBWLyITMhtf3N8VNUBGqdymmAa++38VWrhQ+QHUcNmpyo04LlBmW
HGua/YwFqnxM1crvs9nkoMic81UTvzxYGei9HopDooU93gKyL/stO+0rdL2speYd
9hM75NxnqEf/+2EUuBQzpIwmaK2r81qWG/TtnYU+fTsMfHZB5OA3sweXgxDlYAnl
Rbv+8zwmIl/PqC08Qvgjf2Z5wWTEjoMVL4EQCbliPs+40Op0gZwfz87sz7KP0575
g6uABxX1iGqCAKYMh8dtt9ofV53KvVEs8JS9dt0fQE77/o3DzC/E7YkC65A05hDh
KyAq5TEOfKlnOHcoFTUo056fInOtyjj2ICstKEFWdAi7Uwv+o/idTIzEOKzuD332
PpCT896QwA/3r/sT9Iz0eGYfOcYLJ8bS9sa2rHNaPXm0u11aiZyQjSIhNrZV/uc/
6y8k+VdHwc5Uua7jJPE9dIc0aOU7gImXnMknK0Zx179sfgWKvb3V0NA+lMx499sz
WAQbGiddPPGI09qrU2ZjKfyPLHxqaAj/K1nsrlOy8NauuXCAKe3v3yHUmAb7LPX+
54albSAGO4EJv/60HLoIuyJYAhfDJUJsT+JTTRnzff6Mdr7zsi7jFda8xHhERbCR
k/x8JRN/zlC7USorQeJtZrzDHCqlukl7wTb1cnlE+PCAISPdq/xLL5MoDSEb/UFV
GiY8fpyzxHsbs6lm5ua6AdrlGYMjXfbhb7yJojrcw9yC9qbD7+f4eGW5j5xIwwVf
y9sSMVW9txBD7IJwzpdVVSPvemq79H89tYt6VQBNyfYEfUyIWivqbfd6nHg+l2rC
NfWbZ9g4gT+ovW3puomkRI54BWMBzxHSgaOCoU7oncrD8jABHYo6rWmT9hgVMKfF
279z50s7VjwYl5LzNzGztsSojL7/4Rh96ZnHIJSStboyPuaLw0EWVQ1QT0Jci8ns
8IaQ9rKOoNDXywQ8SaIFRaAs27dO+VTcywLQsusUmn6uLyPK0lUOVQBFhbRlrJip
BJfVyCIABMJ+1rGLq2ja4KpdhdeAjI6c5RwT6B7uAC+34LhNaGm+K7ou3lsS+PAt
ou+dT1TgwoXJ22hBFSNYgnEFMTcgfgPisqIXf3vljl27lSDCnqAEHewzmn/4K5KE
Y1oCh7Ppu5F/qsyWuMpdvpa9O8Ru14rWlSDqm78zwmJofhHCLJmA7ykyTp+DScoc
5vjDmozQ5xazPqZLX0Hwp4Of6pSbtO3ap7sNa3XBrxqWAgrHaR2zrVNTYwwW6TYZ
GS6I0stBB1zD0i11XKsKwzzXuezpm1nTyt8/xXz+2vc3hD7DgQCYEhgty7Ts9T01
mkbSJ+huasv16LbycQ1H/aMm5yWa6/JG4g+v464XJSKcMsr4erG5Eb5Vtw5ddZ7u
z+oH3dldGlZ9gKfpaXJxln5pV0l4niCqGSB/dhF/A7g5B1yNWpEG3rT/9xIPR+UT
0t5PLxSHvGkF3nIFvGF+FSfGX3n7XtIxzVvIyqsuX2yi7/uY1dHhXPCaWXfA0Qrw
jHJIMQNkGeULP+y1LWipVhH7kvOmsxGMuz7iUAOaAmp9UopEp0Jk56Cy0OPaNKD0
TFZzzjPMFzc2DJDnD6RJszgs1QM1hcatZ9n6pG4kZmkKkCPZUvzPZwDTH0fzDM+Y
QIspFmpoNISWP61bTvJWmL9eNNlBT0aB+7M7HhUNZ4B1N1wD4jLeSOrJHpFube36
E8OFTLhZAG6V8jgqNgu0ZbI14gqlNg6Qi0jVDBP7V3JVWi8KnP25Fuw6UKP3YoQj
Qy/ZSN8cqTQSFHtQyLoz4aqUM5F+25qt3FXT/AlU6kzRL2C9gdCIByn78Dv9i8Zv
oqACP68niCSXvFKiSvgKfeH7/NlGOPXtQBzo9WWwfKn+s4nU/hbiYa0GAgovd3nb
bzeewMbxVElfNBNubzY/o4Jikth7iEU8wWyL7X+FA75NztWXThgDB9o+bHKt9yhR
etd+YRIe7eiGeDWSg1sZ7sRbxsug5DZWiYkq/peJXvPUNA49cHtGM9/Lo3nlnsHo
vW+jbyNiu9NrcA/EDQ5UI3D03B8uyl4ipYLBXLXK8DkYTZjxfGu5mlakyYepq68Q
gcBlrUC8fuuWvk7yZoFO3rm6o7JBU3fD7b1BnPd4Tk1nWGB+4Nbem9LWjl4SwWPL
Mp0AeYe3IqqcWHqmcJQkzcNxLg0QNlGIiHfoOU0dWDok5KceIHTOektv8MzqX4MS
HZWD9jbbHvPLd5ZF55OLi1d9Ne1HAIlduNO43gq2aTnrLI61lkKtosTDp+Qsar2t
7GwxfxTHfa9+En6x9z8RZRK9rHXznqJGtgmTO46zy9GYzYcsZVY4fWQvaUT6U0kO
cpnE3KsNpK+TPj7Z2y1vu+pvrj6jRMaxhvSRgO33vQLa48DEp/vvzSgLwhrbRLYi
0Ytpz95Wp63dG7tCZ/hfp4ChDEhubmLs8EeClxXesynfiDABkb2o8+wP3v/0ELZf
LIQzQqTBowULyzy+/SukCesTcj3McI8d1v1QizCxNnjN1wDbgC/oIQptjIn5hwqy
tPtvoITHBwPJDl4d7E2P5B796b5p8vNCxwsiVSJ6KwnE11mqZJjypKZ0ZOKQNqDs
5xIIKsPK4uTaoufhPjwtRjo6wmaupgIGDBG+bbHRpQMRHfUhtuheZEYHpYOdpOwH
QBznoqtqsSF8AAsKqBZOdyZZ7hp2W+GIlPnTI1atnIacoOW70LT7v1TSe7sDrpPy
DLldexxouG5ihV8FFPOncceYnU6rQOsXWlmPIGsDSewvE8HZ+fSi00TvRhYCIxEw
nbLSkqTcoDhrpT9+JUM5SSMAGgcuZA48iRnJxiDwHbJ7RzxSfP2M1VwhAbfB3f9r
vOUli4vPHqzr9zLF8QvlkO52c7fL3s9uh3i1YaXSzd+oY6lOREtuazgFEuaZSJRP
NRvqrMZcoYRyhVfjbh0Fx1Z3BcavCFT/yTOqtjLBqBS8CX7haSwCSURdj8o7xotx
HRsM9stdZ5SPGWh2DQUxGY6GiBEipdB/mBRr9xY0KVnqkWPHrm5XU3/nJwpXqe2u
X+nAsWMiy8Bi2WKrmf6JpB/CBPv5kNNGT2kjoXpuNGHYcMFO7ZzIdXiavU+cDI2r
FoByw601UyU2mc0v7H6I+ikbccpungxam86EZA4kQcr2whsuksPv2W3znArW7hZ2
VH7RXsGzUK3CY4zhkm8KG00r5TIYIhP+rblkOaFbottdUIxZPKlIVnIx8Z2W+TDF
vPy2QHZKa3cLrAprN8cGLOsEuaokMC7hFfNvxnhG81Bhp5/l8jzAcygg4KknosCJ
u3w7laKwtX3Jmnnc71UvXF3F9MijBG5/w+bljxyqKKz1YbtNPv+JAUdXIh3/hhQt
ojmpM6ZStHuMJ30ewUEPZaQfwMppOKwszRCrVkzpMIAFk8YzsxVpG38nISaRMxWF
lQXGIt97vJUKrq1z7JKHWChvKD0BDdwc9BKY/PBTM3D9mt/tvnLC9HvtWdGtpjZg
cQXXRPdtxzbvZcRn2QiyP7ChNlTnPuwzBXWdjFsUqImu+Drg70ri2sePPAhjHRsl
ov9bKarfPimGIiwK9ZKQpM0JL2eHgsTOAX45LFq1X8lTWwQlaM7KzW8HAOmS/gWj
Qh0r/Q9PvRsHm7vDjWCFpIfMC491w12APYnDKD4c7CofifdOgi1oe1dUIpxkjE7V
gAGvOVPcl3GBzZqiv5c29idZob1B3emtq2FI+qRKvytAEqu9lLQUjEJbhEBY/G74
nO/3h113/QnNjPsAMrOiwhxyiFsLA5oUEe8XdKTwGp+ns8y7NzqRbdO/wzVFxQMz
qpsQy5SbEPUubIiXL1gP6edXL1GBalvql6jpBFZeYApmjKnBmGbUMMJppcZqXe8B
WVkKLdzBACd7MHsY0uuHQS03SQnUAkN2m+Rs3C8Ka7xuw9zT7+9svkSec50wKXB+
mXxpYwFeUxPW12Efc5RJ0Aw/H/FQuQdrlp0ifr5CFZ0dh6+PRS0Av+/6TT5lUllq
Qfhz4SbyoUat5L69v82LzFpk6at5yxb3Nng9alAEjC83gXlE0Drql5T0VxFJ8taC
3L4Q4pGgYekEN8RdlJA4LimpRHIjvbdU34oJPsgCYVhPwyvfRL4X+abT8Vfxpvjl
tFh8KyTKCGv+CE7Ek/mZMZG1b42vOQegobd3RwRMjAF6QOCB2lndmiRh/RJE2j2x
v1VHSQkrxROdoovrchxAyGk4Log8PNhSLMNaFCsZvKeWmpP5z1pePbPP/abeZ1lz
qRAkcjSMh02mSzsaZBmsGkTJ9Ki44Wd9OdPJF5Z44Jck0Efdnnzuqcd6tZ6VkGjm
OkN2TYjejFH8rh5Mlcxo1Dz3+RcqUeQ2r3gWB9KZn2j4lDuZpxZXtht1HlLHjA/V
tJzgDqol7TsH4SsPNDfhtNuumqVsl0b4Q2ZFbDs/eQpLqnFvFQcmhCUhj3HfLLZu
qXH14rhT4ieZj4cEGAoexpJRWSxCzom4OCwH6wHSEfwJfhIcVB078K8MGQHE1vu0
nbofqEsoSZEM5QOPPPsIGy/raOFdCY9/Ver+E10nDLsqe7tor+sxywcKBeFHKmS0
JVnJNqCFPW+J/2pu5msSyIC4ry8VhjcKG6RA9n69kPlIttYbO3vfxUmoh4rxSKzm
8/F1ZdfizZkBhLbtt4Ug/Vdsl5AfUKtbm88G/n02ShfsFdjpSH9wlLSXKoox2SS5
0cRA55ywYtHw9AOolte7Bdf55/8U/Er6luKBbYFF0r1AffsJmCZsRxEzfNbZaFWB
oDcglifVGqOgLes8fw0yyQiKPDOB36HAhDcaHyh9BFPWIcRH56nd/bAwjbn5WPsQ
8Cdb48SZtMD6NJIrhLZ3WA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6CvvlLHp3xXfq/+d+mjqnPPHukYs/M6lneSO/0o3pwF7xKRH8hdYWvHUbNhPLhv
GqHSu0nzjLwxpqUHFgPP+/jxtRBUpRikd9XyJQJ4rEwXiSFPA8Q72D0xdLui/TXz
iVvIUVXt5G9BDg7wzC3kThoOhR6VGo4QzMjJdCdUHyKtZJgQyFA2V6KE9kRYojQ8
iZ8o+EYc3KNh1qgCavTkI126Bp3YyMyU6Z97isfzIIwaZiBi27tAFQ7psxFlZsro
kYATCn3TSEYNt1nqxuuLM4/x5DMuxiKmRn08UaNtX9Sc0VRyBcBfHMVLpGNTEZWU
so7go8Xqt1lwC8SJmt9Rg8aoA0n+YvuXSChpRsO91eG31iPp/VXZQyuhu3f57ejU
ArsjnoMRmYbZBlXmwJ20ewD1pWrQCsbyHvCi2sFwCPvbBUx3eUsXplhDoBrx10pV
sa/QaYUE4gRN4zNRKcHeFArr7r34V/kLjQsC1gCtZNnKqirpUgRFryGKyklE1Uas
uy57DsoHCgdTRMGJW/ChPe3pcTLutfrSRuvjIu7YXpkfe+FRLV+E9tetmGv12RTA
8XxOEcNngOOIeW4+1SZCwvqIaruBojUGx6jCZ0h5ijGDyGLe4Zew2LIP7ikXPCkG
nQuuMiG9BBQt0X9U68cud1KE454UKbfmZoAEqadGRYZzlXHTD0qgYbYCsnP75Zae
onHK6q+peEwP/aoPR0cv0Lg+kk5a7gUIV4fQsT1Ky447JYMCqHQtpSFTOJSXnEjf
QsDEJG/Jze7JNr7apWAhf9SBtaAsjQNEMlwN5jF9r/2AGE9KnTv8II91yzmKTyBb
ylXJseNAi5SeY9waCHlQ8Aj4PR+0i+nCe3Oilk/vil5k6wZRhed4rIstEpCGRAws
3hZvP7Xetp4HXJI70c/fyPww7XOD9wfLQIp0W+o3XQe+I9v04W4iGi5j1CmSrMFC
HQWHYENh7vuAOLlUUTx+np8bBrnFDJkIdHh6O4zJ6fS4sNtk9Ys1mSDksAnM82Bh
D5+QjTfZ3AInxJC5ahSVClywAOZbaYZMhLE0/CGLP1C1gjpzAYOAbsVgG12qtc16
fJULrzbUCgCJd/1EYtlLJgedA2ztDiZJ77sqgDjY7l/5IM9G4Bcl5gY9Pjp9XQL3
njLghqtkXSyZsvFZI2nUYUJuyshZ2sWzmqv6SbmEhMZiGfzQNsJeYuGut5q3HCsm
B+E+ZlnezO5EVlY0pUk3HqbvCr+NxN86qc9dmFxnwg+w70rVwHCKgI7YkOt4C5UO
RHHrK9hrEVn8JLhFczOJ66sZr71c0cfxbJVSpXjwuYkNMv1klZ/lJN1n29rKFuCY
owdVzqZ0SneRozcEaj7NSxMGXObOmA7GQGcAyDjRfGZrcyC/PiRM1egMplhitD+h
mfS/vwta+KiPJqsS3pqiUt4bU+HP+FjVqeyCu3PK3GdNz6gfMXDxkQLzIFsbE5R0
F4BmtrciZ0o9O4ZMHC6NtAcyi27Y2ih4qh34Gxxg0YbYTIGFr6/5O4BhWOkXzSbT
Wn7JmzZJslFhXbe3Q3aPaPU6wzxpz19e1pNhGoM26sU47LO1cLDROjaD7CtOq0tx
sEw9HaagUdUAJT0WJKds4p2gjDYNfo1UnU33LBErG0AiHULfWABGh1GbUwq8o+Rh
XS5OoVScFaKmtqFjilXOxg9xmDstPJ8RJOBxxq8cbt9P3XlJ/qgO+qqrtef1OrQN
pZbg7kGrqFHUP3daG6mQ2mldfrAp2361r95dWb4vqZgbiqDcHd5Xrq5TFoG7Tecw
v7xeAkSCvuw8untCirq9txsfllwx58vBIQnKo7dDOU+o+0p+L7a/HyYm6TZrHIMy
P/alopUys/3wMjmxwTk+Wb7VtDhVIWwY5ttuYDfNAd5WGhsIRDVw8d44SnT30bOC
dxXXGEuG0WkyytMEBIGE2faKZnH7uWj9m1ciLG1SG4Y7mnuCxHUev2/Czsi2thO1
YcnH6K/AujMGc6Qd+S/qqv8r9NKau+S279hfxHvu7knArZYZNR7ZGER6quf3jZSb
a+fZ0MekjumzBhlHuHIaRRiOP+4d6Ljy0UJkqdcPyC3Iay3s1biHGV75Fh49ExOu
C1p+1WIhyNsN5ow3pdqgcQkb146OuQ09W4Ws3CYIEayG1HbsEAiu6pQ2izs+uwyq
zd2tupbpKSLaPUABUqhQTWaCx8aoJBU97Ufzu1cpjm1hrX57ZNdE6Z1MFIgjPwiA
jV1XQVRSY7kSuY7KywAqpVs3v4D4ultcX20TMP4vv3uoeGgE0vZOvDp2kzzWA14G
Z9L0c4tQn51BgUBFHNY6scky+c42J6XQ1IY+2LBs+sLwhkyOroTPncr75FPoaNd4
ArDBkWFNpvF91pcJ8ZOMgVWMSr/0lofLkGHqudmeysHwAGu9uvUcbAwDW2MB7egE
z3rtouv1P0k7X8i9EaP62tt6O/tPVlahVSb3X5vT8ednM4Umb73xdgi7blXWeoBX
EXqb1hbLfEbSwbU7Ti6WbL+sZDaZAULIIzJHWtu7A9EXnbfS2sAI2epmMfwDjD9I
rL/3cLqV/fRv4ix7RmPq1WPsBpgxnuFs4rZDIto/AsMJYg29vUnTUhq1ehly+rqh
0lnWudzPzFA/PYkQTxGVb+INFAu3FXykbjxvrLf5LC1ixbThE0mSeeWPTSHuimef
nPky5AkOJoOgpHFK2jRf4jd2GsEnlixsUY2tXFo3XLUddnOEUqfIxAiX/uiH+pCy
wJjB7PQK6xi3H1YWABm4ghj8kGxFDp/tu9X81V5H262Ab0LFhysL8sG9PPw8VjUY
w8vpgxjuuGgZkGx6+Dx/TmnsWuJeJPApjSSg9wzqv80nQHdlup5KJA7ay04Agk7k
G7b8CZsMtMMJjUJEjwJfeA/ce+mlJb1T6pRhc/RpZqRVwEeTCYKeq6JzWsmtVQQJ
0SkqkXN1MZmjdAAuTjFMOCHPjzV/eg4TJB+uOzO831himuMACumL6q4gnJrXCsKD
F82ZLFyC/0Fpf6a3VSUoMnfi+2HV2yq8VI1vxNTpJU+uK3dleCwZcgiMH+6NdF4x
Am+JDTe7FDfLzhIYlt8FcQjpmp/iAQa0vTru9Q0UEiHJv1ZwiNJUQRKcTmNcSHuX
MAU7zXXdphaR6j9Tyw1IIHLFGCwYpJg07vFqPcvY8vZYDkvUUl6ZuVLUD9/0f4th
r4lfKvc50DeCiBpsGrBL6qlc18j2jfP0OhGbovvu41VPLY78x5CD46UJB4y7Z+mT
MZP+al9kRiXSjN01zVDg1t5v4U+SeLYcE/s6aIKJIb2BzC5SI01h8n+DOxnS5MVE
mNYYrPOP23rhbzYHQnincSifz4Kv8YCs2J73/w36FXXE/OK/yyh3Sm+DiibTZgXR
1nV0Okoo+rAYyqVtZVptFBIy6pOSkCrpg/rUG+91IjqvTy49HCstH+rUzzXguB+c
qwrD8ynixHPHsKQiD4NwnJTbdpGWVvrDWhtV3sWBBeUczYX9sNsJzgJ0D2WOlYHE
p9fzgIk3s9XRDR1O8keMR6uE06hlr+QxXaeh4lAzPMBkwhTftrOUQCMfJB0S7NGC
9dtj2CCwHHAED1P/mx1aEt9ptqvUCo5POwPhamzPC8M0inggdfU3gNuGazlLZCCg
azXbnXmK3FHabeVEubSxkq0uE0aGleTe8kl62XR6tU7Md5wxQf3ynAYUTN2HFBmN
LiKf/47xQx5aDKaUokUI+52y5Q9wsQcWW+m1aJPnmFxrKdB1ip82kKYsEu8GvoMI
vamL5HNxHo7axAPgM51dg2DwYnFZl/Zq0xrq1htyrK7MliEtPmck1eN+2GlmeYd+
5z7EY/+kvEYWKGiLpukMXA==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kzd76DThRA2LXCyAhjH3OWa1r56aMJYZnFzxAfupmSqb/AI6KaVdHed9X6XGuro
TsJic5Orlc42a9oGL7rDVgHEzUaVFKG73NPkUIZ35zZDDmDUOFErjhMJ30NvnuOc
rksN8YwTOFRAs5TWFnVZFKo+XLWcIl1J4kPjD8h49i9H7G+Vtt96zmI8BEup3ZM4
BJbuZwVpVoR1GaANpdaE+R7kqmbjO5oTVte8M7ZY8XqS5zGWD6rEOo9pTKneXHrx
L6tJrRPtXskqym441s7M0T2U7BHgQufIlWN/ETqYO7wWdH5GCZLAPKzmS+bwuBgi
dbm3JYTN/o30nwWOT2KuoaWtkqglwQeGbo3gzB5VrIl8EIEHbX2kOHwvyc9JbpGB
qx6Ss7gvyXK8Gsp0RLIn9Bvu8+UqW8+oUSJi7mXSYcvntoat0mp6cdFmE/55OmF/
3CEd3dXhHgoXqFWhvxSiB6SGDduakYlqBJ57oV89aZ8is+aZV0Uqb5gwyQv5Q9ZY
bKI1vhSZJJOuTxts3V9744zHCrqHv0Z9qgDJs8iWmuqCDtGz45qQGghcbyASTtgn
Dd1XMBB6C0tqBiEg+Mgh1+iDEU5IDWzxjEg6FkGDunzEWrqUzBHXwnbSfDmwZ1M0
HPwr/NHcTPZaf2PuXu1YsoyiAAHhq+avqPCYjKpRrLo79MpkFN6vNjhjHceYc8Zg
mvLxRADB8l5YjrSpUlZfdLFaz5YCDiH5+B1pgGd1lFPpRwyiZumPsqvI3P8nGjiJ
Bpb8AgoBtv8YRiiQBePIjyc4J/FOBWmsBtr4aeY9vdzlZbrlFB/6R/EOgqn+egLt
2hpwjqxz8ZC7SrMFrrSoMYTyH6lPKugpzvgxFCRIt9JXLo84lghlZyQuJA5w0vj6
0F+lAMVg8BVrpubvHJp1FomHlPw9x/agnNJLhE+plruj1Le2a3LEMi8zvrvmmhnR
6++0w282cXICQBp2j3E9DW7J79RcLwcAwFRMqZ1VVDOMADR9c+nbdWSQIBxQ96ml
U5d8lRlA/LAqRy/Of1korlUP7uZRTHAPz9M+Ax8LAjIvZXIHUr1Cu1anVO8r5bXA
O+4F+Ell2actuoIe4jjybEpsA/x5bBpKe3+KzvsBYNSwqaLtAFiuuctfNFqHP3KD
kVy7+31V0XcSabk/hGGbHfXY9yNvW6o8gyQJddnPQM2ouFb9xsO1pilYXigY32U6
7ZBLm3OwRk7yLhCrNyttOkpFXHUJ37SyWDl7GKAwszX/+qOUYPd0u5DYkn4FHLR/
dO+1eW5a9NcoyhuYEhhHIx/pkY43ihgSeLMWMR7RWDKHU5av80eQAAOdj+S/hAlY
MzSJl4CebLAqip3aUyhYnN4U5XlM3XluzR6Z1vaMIeusFMBWMvUFor9SjV92L+4h
D36bWYyRvwvnVkBhJ4ITZMEaIKbK+89PaPVBd0liR9fSLGnLMfzD5qwTsRwrcjIa
m5YH5bKyBi5i3YkzQBmeuyg5i4ixf6cJJjaphvE25x9hprsKJNjGohSWdRk2eYNn
zVxdHQBAeveLnIe9fOSP6b0WKnI4Y3Wg3w05N27kTtsZhjpFr9OwbzVPLD+Ncj3E
dFO0qK4DbgM3dd+Y5WFOgImxItTg1PkrdK+MtnQOzFF8ZisXDPXLekMJuPMUERJj
VYeZJq0akR9SYkhy3ZNlyAg75P6SdFOSTfIEPl1nHCre/VWlF2gse7l5/hsj/ziU
qsIRaBYhghWhW3ZTkT77bI5hVzkRxLp1VnsbGtEp8fjtDxDGME23UCI1EoFQ3/F/
7NGgeV1U3ShIpPbt0A2zx+rsaViJ6lHIDCkQzdqhPhnyvuYG8CngIO6wu5WoKM2d
Ood8TlGPD2Nxs2uVFDbpt6jqdbkHaFKD0y/CKJ75MThqlx5PaaYBgo29NOQ8a1oi
OYsC4j7/3xULnWGWjBrdc07NQXm4b5fiYvRdEqNly5iPqXp10fS/ot+C99ho1MZx
GxXr4gQsyddFcFcZafoCY+b70d0eKcd2uJrli5c39mfKxjWpO9JlltrxPSb0+oRk
DqC/hNJdOWcKcvLZbaYdsR0Zp4oOQBhalxq7v0sRK2/1iP05W73DXsRod+DbB/vU
BTuQZC0JSZOdL9HltNtGLjnN5IvoRdYe9XNrjsdn1JOKImIgd6x/m6QGv9OlRMb7
ggIlAcwvb8A78tu+v5vuV0wDjC/TRt1KKKBcd1Z1vpazN7JpnJuCFh50zD0L+h28
ypJZj62RiHNzsIIokFZzAEpnWzGNMlj6Y7Q2JF0Kc9lSUFvBN/u4zGsIA/+BgAhC
KoJCd29DoTHwqID2XDELSSfcTtXCeIREAQu23dwPuiAesbV58o0qcG7X+eXl0Ckl
6HZJYq7lBN7Sw9OwXk6qc2GtcDE4cUpeyTaf1xs+RrrSOyMr80tbvLU6fHwymMhm
2dcW8pQHiRl6tznfIE4ycbxsLuabRKLF64VZwK2N3xBPsFWHbH50xkGyEPrFXh/j
JGB2urN5Ah2j06+gHjcVG+UkEoLecFaOwTJ+KR84kkiMxQCWfURo6jZZ0jnYgObZ
fxVuJiZ0aK862jR4azpOmO0YEcczNCAbmFjY0t2r8YwBrvIJP/E/bSWqVta8KWdO
R6vPlpIyIpZI21EtpiuiCAYbjOkIW7rvcR7MYfy6YttId8PClAovjxqZbsHbxUbn
AO07OVtsEGtybQe/JrBzHBnI9UDEHtYfYS5EfZAujv/tjdaOJpXaRlyCrIAyjjwB
1XpFshuy0m7iic6adjMDC6Mw8hcE4PaKjk/a5Et34wKyINElDB+l7sMwbHvWyvV+
mBbbVnQ20oWidfDHyTzTdPd7c4QtYoLn/KqadEybHnDBe/o1r2rdDQIru0yU2Nx2
YA5A0CHv7u44ONDstCDvk0JLDd+ebyAlNc5Yl0xdMsjqnx/QMRsuoGPsgbqdvuym
LI+cqI88UrJYQMZjGhQpBFZ3dVEibegJVZRjPX2weoHgY5SG3kZ+YjNk8HnKc2+i
gCHzgV4hUdRDN/XB8Z4MW74OK151cje18R/EgPlOgxq5/ZqD6d++cNyxOiWizdDg
Ae085iVdKXUQhpiZm4splNjgYtPpuGtRYdMkX99tKAy2IedjKSeNupTHZPbpT4ui
C5PetMa4eEyE5oMUY9sAOLt+0Z6fwtft6tZYH6mljvVAMVMR+4QE03iHy0WxSEKI
/r2fgO/bP2Ao4fhUNoxPxElrdtkr/XmyQkZO/mXIN2PWJqsmFeHwVWreiLVh/lZ1
GzqHi9n9VwJlR9mcx+9foXp8YJtytyeI8UXBlHVP1Hub3omG90qMOqsNL68bSNG6
tipAZYoEMWwk6q+Bdpl5aGmkn0fFvSR5ukj8+XjdtMP8s7ozFe30i7AMBNNmJ9z3
SxBMN8hB+RToO/FZzZkZ7pb0byHp6UW7z5FIKde8KjC7XI1AB5BrqDB2d9UD2V3Z
Fges3UNONgbyHhtG0s3G5UehxazXQP419nIosXvpLuxNKVM1VrwY34+DKyHNQ8mx
3M52+KrjD6wD+r3akmaG6nWS9IfJQSJi7sF/uSop+byMTpEwbnE1iWQSEqKCq2tA
q80kIN1W5DL/5i/uSFa9SQvEMrCA/j66+nQ0ZlkBAebSUQ/XgViOGSkHB9dOTYPQ
GIKSBWzNm8WfxrlF0Sa4UJ+giFc2QBJMLmzFjZGraplQHv9AdD+RCxXmeYIOmXLh
T3tXu/1ikXvQYTazWkc5itFhrfefyBmdDdbaMKvQDvU13bZvSskroT3Edu9Q5Jg/
ZOUbseZsqvGgPjJUv96+S6OLAcS5eKLr8GGYYMgnJEfBV5wUr1Ww4tj+y1cVvglb
AdnetloPA6lhHwswZTHwZvObxAnElWEOwLBv+Li4ZVw7Vu+mP/rC5PrupGIdy7VU
JRyrEJ9QiZdY5xcOLCzeq8gtu+oR737vaB6f9yyW4WAaQWYkOu7TER4T8TNoULt7
V3jgf+tFd4Qq5dVA5bUCM21ao1D8j6dUaFOSk7JdoS99ZijOVlAU9pHUedp7kw7x
1RlWoY2p8jX5tkfUb53bCGWHxCC9dRiirSTLMCOr+C9Mjntc50vlfNHyq/HBrowO
WHWdKQtWoR2onRZJiujC/hkIUCweP7LPmkLYbcsXFAn2NVhLmnboHAe1aZ+zv65J
x5t8obYTQS5UC3BnzYI6D25tkBQupwaFlat7enJ56xPgFr3o8ksAjay6jqtWaST4
qN/GJgN34c6rmqsZbZGlAr4hnrJbPIol5JHSVd2NZjYJk4Ru618RfZRR8dtg/BS3
`protect END_PROTECTED

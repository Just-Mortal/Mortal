`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYfsquCrILWzleBOzTMoR+PxlmJ10Tt/J0e4zSt36erOnESsNK+v2CLwbvlOtQin
2XYfetkjmlDy5aOihAS7yBg59ZYM3/Io9gftbCK8O2mQCfatb+h4rvFkmMIM6+Cz
+/94DhmxplClcLsfPLCpInH32Gh+GDALwM4OH6q/o1r46c/dslrOqwb1021zqAS9
zyoyjMFwTqU5nLCYKwKiEB6DaQ89JXdtEQqxUnAIqWCw5akMAtHjJwICKboqPbfv
Ddu5Axm4S/SFgab79jj2pxaFXazoISEVwtdcWSZRRj6J4Xt+5kFzbLv/5McnnMT3
Sh+Lx9aXCilL9F35ygJ1y0QhT54Rp1dgavCWuToWGSCRUzGo0Kn2+OAFm+UwdjaF
VqTHbXWwOz6UZu/9cFlV7nN1cjkp6xFUe7Orirf16zhZjXouseYFBBSNGWkAHnv+
zD2JUe2NkDzd9+56OtlXzEYUGsVA3rZkr2LIWIX7hqo=
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chzXbJrM7iVIMKz2Rntgk+ux/mGzkIlw4U2Oo5uo6u7wUv4QxYjoNkJxIK3DcX5m
hy46X6EhM2Xmknyd1J6R9cTGU3vrnVPHnChlTKl/Cnez/5xaP/aacJc/yl8oZ0Pl
2rkj+NK1Hw/FgXKYnKrViBYW0uoSnYuXmepVSvlJtskCJxOrmxc3jgbwG303DCvj
vzoFv2jdvtce55mQ6YE7Ty7odgGXIPgXA/X2/TZyAJ6ge7rfwfXVyBAp+9iyIWtn
4ReCsSnvxUwyLudmsM19HcmdCld2C767uebZ1DCCsl7AmS0GCLd9DxwV37VzaWtn
JtmdTIQmiTKwXoPU0d4r3QN7UQiMmbczN+6gpbT+MZAB86xNoU+4J9pVrrs5EwHv
QaDmk0EPZ88HOnyFDGEzynDcdLMSvy2PBXp+tlwb/dAxoKFznz9IxEqkyNhSbg80
htUIJpPol+lPOkROAGHso3EXtX4YmzxqsvCfNbrKmPFZfzJs3aTagJLZ4QovIVDx
6rpOfBqKGRU9ZzgXxhnqJT/FTbMp1tj67iGmzAz/I3HsTEUmSXcpvJF3h2RZznO3
do7pm95zD1eHkD+VOTOGmFsVY6LQ3H43cmqbDPx218giw+lut1Qs2cshaEr2Ylr2
Tfkk1ffTNom1x5dTfS7Cvt2QfwB7gRom5z/y4TkqykQbBA/PBnwCF11rQLfXGkXO
IW7XF6cpnNFD9nT824+t4ebSG+/OQ5XrmD9DAuyzHX9oDAFvpdgCzS5z9Pjk8fOF
9+WrHkzYWoegxR0fpDvRbW+UGg854/i0kBlFZXV3DRIfl1Mmhd3U7pslLXgmC/mc
lQyrJ86k7ctHjpJhX16JX74INRJvSSjuaHlq551ztPNtIKLLm2yzCKUPI1eyhcav
6lxUw2GoPJAsLXOWehTTjkaApe8XhrUlB4eVEMnS6/OEIw3/ZS01j03nBrvSJjna
BAOP8mGcK7d2eiGrQYT/88EebMC00JE9jxyg9IKhJyMABWiidAnLhmNexm9Ycz/0
K5Fbim1koI9aFUROk7xy7FJXV71TdPDAQbw26Pd675vd3PLMffT3poQ7sqLZo5PK
2Qku6Ndrusy835lhhMMZH5v6f6xUWhO+NtPm4gpE+6liu10D/ECte/fHleiF8oXA
Gu+4GUU7/GuR2W0lIat4UWS2jTAmqu58aFpQbFFRKuJCTCKisb4F+/UHW9sp4YAR
vB3lu3Z0wDxaxjN80l1E04FneOPxyQJiqlK+Jj65w4PUcBWfJ5CUE8fLyvzIE7xP
1XStWzWROvx/0WrJ0IoFAYvBxfHRVjSr6MHvG5h5179goxTLewxDlrk0fVrnBByJ
ZvGqvOjdFw9F1ucymQ2WTOJvFW0NiZwxcU8bzIfb6gasX3wJ+5yLgohN7cnqsfMI
6wCVXe0L0/rnvgynP0oDFGS+uFvuVEvXFomqCxIRbLDSL1glsikHB33wvHQw9l8R
7qKqsznHurQ585gQPirIHqMLIeulG39fib8ImZBwJt2TGIiYObCqJcBP2q4wjx6Z
utA9igZkKXpuCjgnbMpKrQ==
`protect END_PROTECTED

`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QeYZ2cS93/v8rG1ko+TT6fwh/wGMZrk8/I8RoAD21QWuRYiaIPcxdkXWJIsjJkSm
ty/4TiPJAqStpiVVASkLYh/tVD2A2DBmTau5FncOSo0fwPSawt4rwWjAnkyvByau
sDC0P1T/30NgNt2SmL/Tg3VodMYbjLq1mv0tky/EfaKa9tbPjzomsFZWj3uVfzoo
1C3uQDNVrWrB93Lnkv5Exxb8qPwNd6toZDovtnXq0Hx03eQ9hrFe5RzMF+BMD5Cf
d6C4TX+A/ycDZW9/FKZlMJ4n6n7UtguR0hEYot+SPF+UqAI28IiGvzmx1dbtEBUZ
egJDjB9HCks0CtgsTWLmKYnPs3Fsu4gtWalleLmZduwJb4db/dlkq0Dzpt8+1sQH
DuFK6dFVjopMXVdVtdueilF1gopJuBPZv8JhdapyZ+iJ7TqucG8t7bpBnMySzx1t
KX+zO7erBl9ncTdQW2xqsy0c7RcCa04wgR2Uhs8xXWq8Cq7M7odoarikuv0zoBBq
7CzA61yx+Pdb2AHQrEVEIsh3biLogX2uZA32fdknwJcUzk+jNmdtOP5FI8B1A1Do
TUW8ayn2JvziLzRFQDstW76/JVeAIvWOnW+CdYA7mkc=
`protect END_PROTECTED
